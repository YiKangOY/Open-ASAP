module sk128 (in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, in100, in101, in102, in103, in104, in105, in106, in107, in108, in109, in110, in111, in112, in113, in114, in115, in116, in117, in118, in119, in120, in121, in122, in123, in124, in125, in126, in127, in128, in129, in130, in131, in132, in133, in134, in135, in136, in137, in138, in139, in140, in141, in142, in143, in144, in145, in146, in147, in148, in149, in150, in151, in152, in153, in154, in155, in156, in157, in158, in159, in160, in161, in162, in163, in164, in165, in166, in167, in168, in169, in170, in171, in172, in173, in174, in175, in176, in177, in178, in179, in180, in181, in182, in183, in184, in185, in186, in187, in188, in189, in190, in191, in192, in193, in194, in195, in196, in197, in198, in199, in200, in201, in202, in203, in204, in205, in206, in207, in208, in209, in210, in211, in212, in213, in214, in215, in216, in217, in218, in219, in220, in221, in222, in223, in224, in225, in226, in227, in228, in229, in230, in231, in232, in233, in234, in235, in236, in237, in238, in239, in240, in241, in242, in243, in244, in245, in246, in247, in248, in249, in250, in251, in252, in253, in254, in255, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, out30, out31, out32, out33, out34, out35, out36, out37, out38, out39, out40, out41, out42, out43, out44, out45, out46, out47, out48, out49, out50, out51, out52, out53, out54, out55, out56, out57, out58, out59, out60, out61, out62, out63, out64, out65, out66, out67, out68, out69, out70, out71, out72, out73, out74, out75, out76, out77, out78, out79, out80, out81, out82, out83, out84, out85, out86, out87, out88, out89, out90, out91, out92, out93, out94, out95, out96, out97, out98, out99, out100, out101, out102, out103, out104, out105, out106, out107, out108, out109, out110, out111, out112, out113, out114, out115, out116, out117, out118, out119, out120, out121, out122, out123, out124, out125, out126, out127, out128, );
input in0;
input in1;
input in2;
input in3;
input in4;
input in5;
input in6;
input in7;
input in8;
input in9;
input in10;
input in11;
input in12;
input in13;
input in14;
input in15;
input in16;
input in17;
input in18;
input in19;
input in20;
input in21;
input in22;
input in23;
input in24;
input in25;
input in26;
input in27;
input in28;
input in29;
input in30;
input in31;
input in32;
input in33;
input in34;
input in35;
input in36;
input in37;
input in38;
input in39;
input in40;
input in41;
input in42;
input in43;
input in44;
input in45;
input in46;
input in47;
input in48;
input in49;
input in50;
input in51;
input in52;
input in53;
input in54;
input in55;
input in56;
input in57;
input in58;
input in59;
input in60;
input in61;
input in62;
input in63;
input in64;
input in65;
input in66;
input in67;
input in68;
input in69;
input in70;
input in71;
input in72;
input in73;
input in74;
input in75;
input in76;
input in77;
input in78;
input in79;
input in80;
input in81;
input in82;
input in83;
input in84;
input in85;
input in86;
input in87;
input in88;
input in89;
input in90;
input in91;
input in92;
input in93;
input in94;
input in95;
input in96;
input in97;
input in98;
input in99;
input in100;
input in101;
input in102;
input in103;
input in104;
input in105;
input in106;
input in107;
input in108;
input in109;
input in110;
input in111;
input in112;
input in113;
input in114;
input in115;
input in116;
input in117;
input in118;
input in119;
input in120;
input in121;
input in122;
input in123;
input in124;
input in125;
input in126;
input in127;
input in128;
input in129;
input in130;
input in131;
input in132;
input in133;
input in134;
input in135;
input in136;
input in137;
input in138;
input in139;
input in140;
input in141;
input in142;
input in143;
input in144;
input in145;
input in146;
input in147;
input in148;
input in149;
input in150;
input in151;
input in152;
input in153;
input in154;
input in155;
input in156;
input in157;
input in158;
input in159;
input in160;
input in161;
input in162;
input in163;
input in164;
input in165;
input in166;
input in167;
input in168;
input in169;
input in170;
input in171;
input in172;
input in173;
input in174;
input in175;
input in176;
input in177;
input in178;
input in179;
input in180;
input in181;
input in182;
input in183;
input in184;
input in185;
input in186;
input in187;
input in188;
input in189;
input in190;
input in191;
input in192;
input in193;
input in194;
input in195;
input in196;
input in197;
input in198;
input in199;
input in200;
input in201;
input in202;
input in203;
input in204;
input in205;
input in206;
input in207;
input in208;
input in209;
input in210;
input in211;
input in212;
input in213;
input in214;
input in215;
input in216;
input in217;
input in218;
input in219;
input in220;
input in221;
input in222;
input in223;
input in224;
input in225;
input in226;
input in227;
input in228;
input in229;
input in230;
input in231;
input in232;
input in233;
input in234;
input in235;
input in236;
input in237;
input in238;
input in239;
input in240;
input in241;
input in242;
input in243;
input in244;
input in245;
input in246;
input in247;
input in248;
input in249;
input in250;
input in251;
input in252;
input in253;
input in254;
input in255;
output out0;
output out1;
output out2;
output out3;
output out4;
output out5;
output out6;
output out7;
output out8;
output out9;
output out10;
output out11;
output out12;
output out13;
output out14;
output out15;
output out16;
output out17;
output out18;
output out19;
output out20;
output out21;
output out22;
output out23;
output out24;
output out25;
output out26;
output out27;
output out28;
output out29;
output out30;
output out31;
output out32;
output out33;
output out34;
output out35;
output out36;
output out37;
output out38;
output out39;
output out40;
output out41;
output out42;
output out43;
output out44;
output out45;
output out46;
output out47;
output out48;
output out49;
output out50;
output out51;
output out52;
output out53;
output out54;
output out55;
output out56;
output out57;
output out58;
output out59;
output out60;
output out61;
output out62;
output out63;
output out64;
output out65;
output out66;
output out67;
output out68;
output out69;
output out70;
output out71;
output out72;
output out73;
output out74;
output out75;
output out76;
output out77;
output out78;
output out79;
output out80;
output out81;
output out82;
output out83;
output out84;
output out85;
output out86;
output out87;
output out88;
output out89;
output out90;
output out91;
output out92;
output out93;
output out94;
output out95;
output out96;
output out97;
output out98;
output out99;
output out100;
output out101;
output out102;
output out103;
output out104;
output out105;
output out106;
output out107;
output out108;
output out109;
output out110;
output out111;
output out112;
output out113;
output out114;
output out115;
output out116;
output out117;
output out118;
output out119;
output out120;
output out121;
output out122;
output out123;
output out124;
output out125;
output out126;
output out127;
output out128;
wire var0;
wire var1;
wire var2;
wire var3;
wire var4;
wire var5;
wire var6;
wire var7;
wire var8;
wire var9;
wire var10;
wire var11;
wire var12;
wire var13;
wire var14;
wire var15;
wire var16;
wire var17;
wire var18;
wire var19;
wire var20;
wire var21;
wire var22;
wire var23;
wire var24;
wire var25;
wire var26;
wire var27;
wire var28;
wire var29;
wire var30;
wire var31;
wire var32;
wire var33;
wire var34;
wire var35;
wire var36;
wire var37;
wire var38;
wire var39;
wire var40;
wire var41;
wire var42;
wire var43;
wire var44;
wire var45;
wire var46;
wire var47;
wire var48;
wire var49;
wire var50;
wire var51;
wire var52;
wire var53;
wire var54;
wire var55;
wire var56;
wire var57;
wire var58;
wire var59;
wire var60;
wire var61;
wire var62;
wire var63;
wire var64;
wire var65;
wire var66;
wire var67;
wire var68;
wire var69;
wire var70;
wire var71;
wire var72;
wire var73;
wire var74;
wire var75;
wire var76;
wire var77;
wire var78;
wire var79;
wire var80;
wire var81;
wire var82;
wire var83;
wire var84;
wire var85;
wire var86;
wire var87;
wire var88;
wire var89;
wire var90;
wire var91;
wire var92;
wire var93;
wire var94;
wire var95;
wire var96;
wire var97;
wire var98;
wire var99;
wire var100;
wire var101;
wire var102;
wire var103;
wire var104;
wire var105;
wire var106;
wire var107;
wire var108;
wire var109;
wire var110;
wire var111;
wire var112;
wire var113;
wire var114;
wire var115;
wire var116;
wire var117;
wire var118;
wire var119;
wire var120;
wire var121;
wire var122;
wire var123;
wire var124;
wire var125;
wire var126;
wire var127;
wire var128;
wire var129;
wire var130;
wire var131;
wire var132;
wire var133;
wire var134;
wire var135;
wire var136;
wire var137;
wire var138;
wire var139;
wire var140;
wire var141;
wire var142;
wire var143;
wire var144;
wire var145;
wire var146;
wire var147;
wire var148;
wire var149;
wire var150;
wire var151;
wire var152;
wire var153;
wire var154;
wire var155;
wire var156;
wire var157;
wire var158;
wire var159;
wire var160;
wire var161;
wire var162;
wire var163;
wire var164;
wire var165;
wire var166;
wire var167;
wire var168;
wire var169;
wire var170;
wire var171;
wire var172;
wire var173;
wire var174;
wire var175;
wire var176;
wire var177;
wire var178;
wire var179;
wire var180;
wire var181;
wire var182;
wire var183;
wire var184;
wire var185;
wire var186;
wire var187;
wire var188;
wire var189;
wire var190;
wire var191;
wire var192;
wire var193;
wire var194;
wire var195;
wire var196;
wire var197;
wire var198;
wire var199;
wire var200;
wire var201;
wire var202;
wire var203;
wire var204;
wire var205;
wire var206;
wire var207;
wire var208;
wire var209;
wire var210;
wire var211;
wire var212;
wire var213;
wire var214;
wire var215;
wire var216;
wire var217;
wire var218;
wire var219;
wire var220;
wire var221;
wire var222;
wire var223;
wire var224;
wire var225;
wire var226;
wire var227;
wire var228;
wire var229;
wire var230;
wire var231;
wire var232;
wire var233;
wire var234;
wire var235;
wire var236;
wire var237;
wire var238;
wire var239;
wire var240;
wire var241;
wire var242;
wire var243;
wire var244;
wire var245;
wire var246;
wire var247;
wire var248;
wire var249;
wire var250;
wire var251;
wire var252;
wire var253;
wire var254;
wire var255;
wire var256;
wire var257;
wire var258;
wire var259;
wire var260;
wire var261;
wire var262;
wire var263;
wire var264;
wire var265;
wire var266;
wire var267;
wire var268;
wire var269;
wire var270;
wire var271;
wire var272;
wire var273;
wire var274;
wire var275;
wire var276;
wire var277;
wire var278;
wire var279;
wire var280;
wire var281;
wire var282;
wire var283;
wire var284;
wire var285;
wire var286;
wire var287;
wire var288;
wire var289;
wire var290;
wire var291;
wire var292;
wire var293;
wire var294;
wire var295;
wire var296;
wire var297;
wire var298;
wire var299;
wire var300;
wire var301;
wire var302;
wire var303;
wire var304;
wire var305;
wire var306;
wire var307;
wire var308;
wire var309;
wire var310;
wire var311;
wire var312;
wire var313;
wire var314;
wire var315;
wire var316;
wire var317;
wire var318;
wire var319;
wire var320;
wire var321;
wire var322;
wire var323;
wire var324;
wire var325;
wire var326;
wire var327;
wire var328;
wire var329;
wire var330;
wire var331;
wire var332;
wire var333;
wire var334;
wire var335;
wire var336;
wire var337;
wire var338;
wire var339;
wire var340;
wire var341;
wire var342;
wire var343;
wire var344;
wire var345;
wire var346;
wire var347;
wire var348;
wire var349;
wire var350;
wire var351;
wire var352;
wire var353;
wire var354;
wire var355;
wire var356;
wire var357;
wire var358;
wire var359;
wire var360;
wire var361;
wire var362;
wire var363;
wire var364;
wire var365;
wire var366;
wire var367;
wire var368;
wire var369;
wire var370;
wire var371;
wire var372;
wire var373;
wire var374;
wire var375;
wire var376;
wire var377;
wire var378;
wire var379;
wire var380;
wire var381;
wire var382;
wire var383;
wire var384;
wire var385;
wire var386;
wire var387;
wire var388;
wire var389;
wire var390;
wire var391;
wire var392;
wire var393;
wire var394;
wire var395;
wire var396;
wire var397;
wire var398;
wire var399;
wire var400;
wire var401;
wire var402;
wire var403;
wire var404;
wire var405;
wire var406;
wire var407;
wire var408;
wire var409;
wire var410;
wire var411;
wire var412;
wire var413;
wire var414;
wire var415;
wire var416;
wire var417;
wire var418;
wire var419;
wire var420;
wire var421;
wire var422;
wire var423;
wire var424;
wire var425;
wire var426;
wire var427;
wire var428;
wire var429;
wire var430;
wire var431;
wire var432;
wire var433;
wire var434;
wire var435;
wire var436;
wire var437;
wire var438;
wire var439;
wire var440;
wire var441;
wire var442;
wire var443;
wire var444;
wire var445;
wire var446;
wire var447;
wire var448;
wire var449;
wire var450;
wire var451;
wire var452;
wire var453;
wire var454;
wire var455;
wire var456;
wire var457;
wire var458;
wire var459;
wire var460;
wire var461;
wire var462;
wire var463;
wire var464;
wire var465;
wire var466;
wire var467;
wire var468;
wire var469;
wire var470;
wire var471;
wire var472;
wire var473;
wire var474;
wire var475;
wire var476;
wire var477;
wire var478;
wire var479;
wire var480;
wire var481;
wire var482;
wire var483;
wire var484;
wire var485;
wire var486;
wire var487;
wire var488;
wire var489;
wire var490;
wire var491;
wire var492;
wire var493;
wire var494;
wire var495;
wire var496;
wire var497;
wire var498;
wire var499;
wire var500;
wire var501;
wire var502;
wire var503;
wire var504;
wire var505;
wire var506;
wire var507;
wire var508;
wire var509;
wire var510;
wire var511;
wire var512;
wire var513;
wire var514;
wire var515;
wire var516;
wire var517;
wire var518;
wire var519;
wire var520;
wire var521;
wire var522;
wire var523;
wire var524;
wire var525;
wire var526;
wire var527;
wire var528;
wire var529;
wire var530;
wire var531;
wire var532;
wire var533;
wire var534;
wire var535;
wire var536;
wire var537;
wire var538;
wire var539;
wire var540;
wire var541;
wire var542;
wire var543;
wire var544;
wire var545;
wire var546;
wire var547;
wire var548;
wire var549;
wire var550;
wire var551;
wire var552;
wire var553;
wire var554;
wire var555;
wire var556;
wire var557;
wire var558;
wire var559;
wire var560;
wire var561;
wire var562;
wire var563;
wire var564;
wire var565;
wire var566;
wire var567;
wire var568;
wire var569;
wire var570;
wire var571;
wire var572;
wire var573;
wire var574;
wire var575;
wire var576;
wire var577;
wire var578;
wire var579;
wire var580;
wire var581;
wire var582;
wire var583;
wire var584;
wire var585;
wire var586;
wire var587;
wire var588;
wire var589;
wire var590;
wire var591;
wire var592;
wire var593;
wire var594;
wire var595;
wire var596;
wire var597;
wire var598;
wire var599;
wire var600;
wire var601;
wire var602;
wire var603;
wire var604;
wire var605;
wire var606;
wire var607;
wire var608;
wire var609;
wire var610;
wire var611;
wire var612;
wire var613;
wire var614;
wire var615;
wire var616;
wire var617;
wire var618;
wire var619;
wire var620;
wire var621;
wire var622;
wire var623;
wire var624;
wire var625;
wire var626;
wire var627;
wire var628;
wire var629;
wire var630;
wire var631;
wire var632;
wire var633;
wire var634;
wire var635;
wire var636;
wire var637;
wire var638;
wire var639;
wire var640;
wire var641;
wire var642;
wire var643;
wire var644;
wire var645;
wire var646;
wire var647;
wire var648;
wire var649;
wire var650;
wire var651;
wire var652;
wire var653;
wire var654;
wire var655;
wire var656;
wire var657;
wire var658;
wire var659;
wire var660;
wire var661;
wire var662;
wire var663;
wire var664;
wire var665;
wire var666;
wire var667;
wire var668;
wire var669;
wire var670;
wire var671;
wire var672;
wire var673;
wire var674;
wire var675;
wire var676;
wire var677;
wire var678;
wire var679;
wire var680;
wire var681;
wire var682;
wire var683;
wire var684;
wire var685;
wire var686;
wire var687;
wire var688;
wire var689;
wire var690;
wire var691;
wire var692;
wire var693;
wire var694;
wire var695;
wire var696;
wire var697;
wire var698;
wire var699;
wire var700;
wire var701;
wire var702;
wire var703;
wire var704;
wire var705;
wire var706;
wire var707;
wire var708;
wire var709;
wire var710;
wire var711;
wire var712;
wire var713;
wire var714;
wire var715;
wire var716;
wire var717;
wire var718;
wire var719;
wire var720;
wire var721;
wire var722;
wire var723;
wire var724;
wire var725;
wire var726;
wire var727;
wire var728;
wire var729;
wire var730;
wire var731;
wire var732;
wire var733;
wire var734;
wire var735;
wire var736;
wire var737;
wire var738;
wire var739;
wire var740;
wire var741;
wire var742;
wire var743;
wire var744;
wire var745;
wire var746;
wire var747;
wire var748;
wire var749;
wire var750;
wire var751;
wire var752;
wire var753;
wire var754;
wire var755;
wire var756;
wire var757;
wire var758;
wire var759;
wire var760;
wire var761;
wire var762;
wire var763;
wire var764;
wire var765;
wire var766;
wire var767;
wire var768;
wire var769;
wire var770;
wire var771;
wire var772;
wire var773;
wire var774;
wire var775;
wire var776;
wire var777;
wire var778;
wire var779;
wire var780;
wire var781;
wire var782;
wire var783;
wire var784;
wire var785;
wire var786;
wire var787;
wire var788;
wire var789;
wire var790;
wire var791;
wire var792;
wire var793;
wire var794;
wire var795;
wire var796;
wire var797;
wire var798;
wire var799;
wire var800;
wire var801;
wire var802;
wire var803;
wire var804;
wire var805;
wire var806;
wire var807;
wire var808;
wire var809;
wire var810;
wire var811;
wire var812;
wire var813;
wire var814;
wire var815;
wire var816;
wire var817;
wire var818;
wire var819;
wire var820;
wire var821;
wire var822;
wire var823;
wire var824;
wire var825;
wire var826;
wire var827;
wire var828;
wire var829;
wire var830;
wire var831;
wire var832;
wire var833;
wire var834;
wire var835;
wire var836;
wire var837;
wire var838;
wire var839;
wire var840;
wire var841;
wire var842;
wire var843;
wire var844;
wire var845;
wire var846;
wire var847;
wire var848;
wire var849;
wire var850;
wire var851;
wire var852;
wire var853;
wire var854;
wire var855;
wire var856;
wire var857;
wire var858;
wire var859;
wire var860;
wire var861;
wire var862;
wire var863;
wire var864;
wire var865;
wire var866;
wire var867;
wire var868;
wire var869;
wire var870;
wire var871;
wire var872;
wire var873;
wire var874;
wire var875;
wire var876;
wire var877;
wire var878;
wire var879;
wire var880;
wire var881;
wire var882;
wire var883;
wire var884;
wire var885;
wire var886;
wire var887;
wire var888;
wire var889;
wire var890;
wire var891;
wire var892;
wire var893;
wire var894;
wire var895;
wire var896;
wire var897;
wire var898;
wire var899;
wire var900;
wire var901;
wire var902;
wire var903;
wire var904;
wire var905;
wire var906;
wire var907;
wire var908;
wire var909;
wire var910;
wire var911;
wire var912;
wire var913;
wire var914;
wire var915;
wire var916;
wire var917;
wire var918;
wire var919;
wire var920;
wire var921;
wire var922;
wire var923;
wire var924;
wire var925;
wire var926;
wire var927;
wire var928;
wire var929;
wire var930;
wire var931;
wire var932;
wire var933;
wire var934;
wire var935;
wire var936;
wire var937;
wire var938;
wire var939;
wire var940;
wire var941;
wire var942;
wire var943;
wire var944;
wire var945;
wire var946;
wire var947;
wire var948;
wire var949;
wire var950;
wire var951;
wire var952;
wire var953;
wire var954;
wire var955;
wire var956;
wire var957;
wire var958;
wire var959;
wire var960;
wire var961;
wire var962;
wire var963;
wire var964;
wire var965;
wire var966;
wire var967;
wire var968;
wire var969;
wire var970;
wire var971;
wire var972;
wire var973;
wire var974;
wire var975;
wire var976;
wire var977;
wire var978;
wire var979;
wire var980;
wire var981;
wire var982;
wire var983;
wire var984;
wire var985;
wire var986;
wire var987;
wire var988;
wire var989;
wire var990;
wire var991;
wire var992;
wire var993;
wire var994;
wire var995;
wire var996;
wire var997;
wire var998;
wire var999;
wire var1000;
wire var1001;
wire var1002;
wire var1003;
wire var1004;
wire var1005;
wire var1006;
wire var1007;
wire var1008;
wire var1009;
wire var1010;
wire var1011;
wire var1012;
wire var1013;
wire var1014;
wire var1015;
wire var1016;
wire var1017;
wire var1018;
wire var1019;
wire var1020;
wire var1021;
wire var1022;
wire var1023;
wire var1024;
wire var1025;
wire var1026;
wire var1027;
wire var1028;
wire var1029;
wire var1030;
wire var1031;
wire var1032;
wire var1033;
wire var1034;
wire var1035;
wire var1036;
wire var1037;
wire var1038;
wire var1039;
wire var1040;
wire var1041;
wire var1042;
wire var1043;
wire var1044;
wire var1045;
wire var1046;
wire var1047;
wire var1048;
wire var1049;
wire var1050;
wire var1051;
wire var1052;
wire var1053;
wire var1054;
wire var1055;
wire var1056;
wire var1057;
wire var1058;
wire var1059;
wire var1060;
wire var1061;
wire var1062;
wire var1063;
wire var1064;
wire var1065;
wire var1066;
wire var1067;
wire var1068;
wire var1069;
wire var1070;
wire var1071;
wire var1072;
wire var1073;
wire var1074;
wire var1075;
wire var1076;
wire var1077;
wire var1078;
wire var1079;
wire var1080;
wire var1081;
wire var1082;
wire var1083;
wire var1084;
wire var1085;
wire var1086;
wire var1087;
wire var1088;
wire var1089;
wire var1090;
wire var1091;
wire var1092;
wire var1093;
wire var1094;
wire var1095;
wire var1096;
wire var1097;
wire var1098;
wire var1099;
wire var1100;
wire var1101;
wire var1102;
wire var1103;
wire var1104;
wire var1105;
wire var1106;
wire var1107;
wire var1108;
wire var1109;
wire var1110;
wire var1111;
wire var1112;
wire var1113;
wire var1114;
wire var1115;
wire var1116;
wire var1117;
wire var1118;
wire var1119;
wire var1120;
wire var1121;
wire var1122;
wire var1123;
wire var1124;
wire var1125;
wire var1126;
wire var1127;
wire var1128;
wire var1129;
wire var1130;
wire var1131;
wire var1132;
wire var1133;
wire var1134;
wire var1135;
wire var1136;
wire var1137;
wire var1138;
wire var1139;
wire var1140;
wire var1141;
wire var1142;
wire var1143;
wire var1144;
wire var1145;
wire var1146;
wire var1147;
wire var1148;
wire var1149;
wire var1150;
wire var1151;
wire var1152;
wire var1153;
wire var1154;
wire var1155;
wire var1156;
wire var1157;
wire var1158;
wire var1159;
wire var1160;
wire var1161;
wire var1162;
wire var1163;
wire var1164;
wire var1165;
wire var1166;
wire var1167;
wire var1168;
wire var1169;
wire var1170;
wire var1171;
wire var1172;
wire var1173;
wire var1174;
wire var1175;
wire var1176;
wire var1177;
wire var1178;
wire var1179;
wire var1180;
wire var1181;
wire var1182;
wire var1183;
wire var1184;
wire var1185;
wire var1186;
wire var1187;
wire var1188;
wire var1189;
wire var1190;
wire var1191;
wire var1192;
wire var1193;
wire var1194;
wire var1195;
wire var1196;
wire var1197;
wire var1198;
wire var1199;
wire var1200;
wire var1201;
wire var1202;
wire var1203;
wire var1204;
wire var1205;
wire var1206;
wire var1207;
wire var1208;
wire var1209;
wire var1210;
wire var1211;
wire var1212;
wire var1213;
wire var1214;
wire var1215;
wire var1216;
wire var1217;
wire var1218;
wire var1219;
wire var1220;
wire var1221;
wire var1222;
wire var1223;
wire var1224;
wire var1225;
wire var1226;
wire var1227;
wire var1228;
wire var1229;
wire var1230;
wire var1231;
wire var1232;
wire var1233;
wire var1234;
wire var1235;
wire var1236;
wire var1237;
wire var1238;
wire var1239;
wire var1240;
wire var1241;
wire var1242;
wire var1243;
wire var1244;
wire var1245;
wire var1246;
wire var1247;
wire var1248;
wire var1249;
wire var1250;
wire var1251;
wire var1252;
wire var1253;
wire var1254;
wire var1255;
wire var1256;
wire var1257;
wire var1258;
wire var1259;
wire var1260;
wire var1261;
wire var1262;
wire var1263;
wire var1264;
wire var1265;
wire var1266;
wire var1267;
wire var1268;
wire var1269;
wire var1270;
wire var1271;
wire var1272;
wire var1273;
wire var1274;
wire var1275;
wire var1276;
wire var1277;
wire var1278;
wire var1279;
wire var1280;
wire var1281;
wire var1282;
wire var1283;
wire var1284;
wire var1285;
wire var1286;
wire var1287;
wire var1288;
wire var1289;
wire var1290;
wire var1291;
wire var1292;
wire var1293;
wire var1294;
wire var1295;
wire var1296;
wire var1297;
wire var1298;
wire var1299;
wire var1300;
wire var1301;
wire var1302;
wire var1303;
wire var1304;
wire var1305;
wire var1306;
wire var1307;
wire var1308;
wire var1309;
wire var1310;
wire var1311;
wire var1312;
wire var1313;
wire var1314;
wire var1315;
wire var1316;
wire var1317;
wire var1318;
wire var1319;
wire var1320;
wire var1321;
wire var1322;
wire var1323;
wire var1324;
wire var1325;
wire var1326;
wire var1327;
wire var1328;
wire var1329;
wire var1330;
wire var1331;
wire var1332;
wire var1333;
wire var1334;
wire var1335;
wire var1336;
wire var1337;
wire var1338;
wire var1339;
wire var1340;
wire var1341;
wire var1342;
wire var1343;
wire var1344;
wire var1345;
wire var1346;
wire var1347;
wire var1348;
wire var1349;
wire var1350;
wire var1351;
wire var1352;
wire var1353;
wire var1354;
wire var1355;
wire var1356;
wire var1357;
wire var1358;
wire var1359;
wire var1360;
wire var1361;
wire var1362;
wire var1363;
wire var1364;
wire var1365;
wire var1366;
wire var1367;
wire var1368;
wire var1369;
wire var1370;
wire var1371;
wire var1372;
wire var1373;
wire var1374;
wire var1375;
wire var1376;
wire var1377;
wire var1378;
wire var1379;
wire var1380;
wire var1381;
wire var1382;
wire var1383;
wire var1384;
wire var1385;
wire var1386;
wire var1387;
wire var1388;
wire var1389;
wire var1390;
wire var1391;
wire var1392;
wire var1393;
wire var1394;
wire var1395;
wire var1396;
wire var1397;
wire var1398;
wire var1399;
wire var1400;
wire var1401;
wire var1402;
wire var1403;
wire var1404;
wire var1405;
wire var1406;
wire var1407;
wire var1408;
wire var1409;
wire var1410;
wire var1411;
wire var1412;
wire var1413;
wire var1414;
wire var1415;
wire var1416;
wire var1417;
wire var1418;
wire var1419;
wire var1420;
wire var1421;
wire var1422;
wire var1423;
wire var1424;
wire var1425;
wire var1426;
wire var1427;
wire var1428;
wire var1429;
wire var1430;
wire var1431;
wire var1432;
wire var1433;
wire var1434;
wire var1435;
wire var1436;
wire var1437;
wire var1438;
wire var1439;
wire var1440;
wire var1441;
wire var1442;
wire var1443;
wire var1444;
wire var1445;
wire var1446;
wire var1447;
wire var1448;
wire var1449;
wire var1450;
wire var1451;
wire var1452;
wire var1453;
wire var1454;
wire var1455;
wire var1456;
wire var1457;
wire var1458;
wire var1459;
wire var1460;
wire var1461;
wire var1462;
wire var1463;
wire var1464;
wire var1465;
wire var1466;
wire var1467;
wire var1468;
wire var1469;
wire var1470;
wire var1471;
wire var1472;
wire var1473;
wire var1474;
wire var1475;
wire var1476;
wire var1477;
wire var1478;
wire var1479;
wire var1480;
wire var1481;
wire var1482;
wire var1483;
wire var1484;
wire var1485;
wire var1486;
wire var1487;
wire var1488;
wire var1489;
wire var1490;
wire var1491;
wire var1492;
wire var1493;
wire var1494;
wire var1495;
wire var1496;
wire var1497;
wire var1498;
wire var1499;
wire var1500;
wire var1501;
wire var1502;
wire var1503;
wire var1504;
wire var1505;
wire var1506;
wire var1507;
wire var1508;
wire var1509;
wire var1510;
wire var1511;
wire var1512;
wire var1513;
wire var1514;
wire var1515;
wire var1516;
wire var1517;
wire var1518;
wire var1519;
wire var1520;
wire var1521;
wire var1522;
wire var1523;
wire var1524;
wire var1525;
wire var1526;
wire var1527;
wire var1528;
wire var1529;
wire var1530;
wire var1531;
wire var1532;
wire var1533;
wire var1534;
wire var1535;
wire var1536;
wire var1537;
wire var1538;
wire var1539;
wire var1540;
wire var1541;
wire var1542;
wire var1543;
wire var1544;
wire var1545;
wire var1546;
wire var1547;
wire var1548;
wire var1549;
wire var1550;
wire var1551;
wire var1552;
wire var1553;
wire var1554;
wire var1555;
wire var1556;
wire var1557;
wire var1558;
wire var1559;
wire var1560;
wire var1561;
wire var1562;
wire var1563;
wire var1564;
wire var1565;
wire var1566;
wire var1567;
wire var1568;
wire var1569;
wire var1570;
wire var1571;
wire var1572;
wire var1573;
wire var1574;
wire var1575;
wire var1576;
wire var1577;
wire var1578;
wire var1579;
wire var1580;
wire var1581;
wire var1582;
wire var1583;
wire var1584;
wire var1585;
wire var1586;
wire var1587;
wire var1588;
wire var1589;
wire var1590;
wire var1591;
wire var1592;
wire var1593;
wire var1594;
wire var1595;
wire var1596;
wire var1597;
wire var1598;
wire var1599;
assign var0 = in255 & in127;
assign var1 = in254 & in126;
assign var2 = in253 & in125;
assign var3 = in252 & in124;
assign var4 = in251 & in123;
assign var5 = in250 & in122;
assign var6 = in249 & in121;
assign var7 = in248 & in120;
assign var8 = in247 & in119;
assign var9 = in246 & in118;
assign var10 = in245 & in117;
assign var11 = in244 & in116;
assign var12 = in243 & in115;
assign var13 = in242 & in114;
assign var14 = in241 & in113;
assign var15 = in240 & in112;
assign var16 = in239 & in111;
assign var17 = in238 & in110;
assign var18 = in237 & in109;
assign var19 = in236 & in108;
assign var20 = in235 & in107;
assign var21 = in234 & in106;
assign var22 = in233 & in105;
assign var23 = in232 & in104;
assign var24 = in231 & in103;
assign var25 = in230 & in102;
assign var26 = in229 & in101;
assign var27 = in228 & in100;
assign var28 = in227 & in99;
assign var29 = in226 & in98;
assign var30 = in225 & in97;
assign var31 = in224 & in96;
assign var32 = in223 & in95;
assign var33 = in222 & in94;
assign var34 = in221 & in93;
assign var35 = in220 & in92;
assign var36 = in219 & in91;
assign var37 = in218 & in90;
assign var38 = in217 & in89;
assign var39 = in216 & in88;
assign var40 = in215 & in87;
assign var41 = in214 & in86;
assign var42 = in213 & in85;
assign var43 = in212 & in84;
assign var44 = in211 & in83;
assign var45 = in210 & in82;
assign var46 = in209 & in81;
assign var47 = in208 & in80;
assign var48 = in207 & in79;
assign var49 = in206 & in78;
assign var50 = in205 & in77;
assign var51 = in204 & in76;
assign var52 = in203 & in75;
assign var53 = in202 & in74;
assign var54 = in201 & in73;
assign var55 = in200 & in72;
assign var56 = in199 & in71;
assign var57 = in198 & in70;
assign var58 = in197 & in69;
assign var59 = in196 & in68;
assign var60 = in195 & in67;
assign var61 = in194 & in66;
assign var62 = in193 & in65;
assign var63 = in192 & in64;
assign var64 = in191 & in63;
assign var65 = in190 & in62;
assign var66 = in189 & in61;
assign var67 = in188 & in60;
assign var68 = in187 & in59;
assign var69 = in186 & in58;
assign var70 = in185 & in57;
assign var71 = in184 & in56;
assign var72 = in183 & in55;
assign var73 = in182 & in54;
assign var74 = in181 & in53;
assign var75 = in180 & in52;
assign var76 = in179 & in51;
assign var77 = in178 & in50;
assign var78 = in177 & in49;
assign var79 = in176 & in48;
assign var80 = in175 & in47;
assign var81 = in174 & in46;
assign var82 = in173 & in45;
assign var83 = in172 & in44;
assign var84 = in171 & in43;
assign var85 = in170 & in42;
assign var86 = in169 & in41;
assign var87 = in168 & in40;
assign var88 = in167 & in39;
assign var89 = in166 & in38;
assign var90 = in165 & in37;
assign var91 = in164 & in36;
assign var92 = in163 & in35;
assign var93 = in162 & in34;
assign var94 = in161 & in33;
assign var95 = in160 & in32;
assign var96 = in159 & in31;
assign var97 = in158 & in30;
assign var98 = in157 & in29;
assign var99 = in156 & in28;
assign var100 = in155 & in27;
assign var101 = in154 & in26;
assign var102 = in153 & in25;
assign var103 = in152 & in24;
assign var104 = in151 & in23;
assign var105 = in150 & in22;
assign var106 = in149 & in21;
assign var107 = in148 & in20;
assign var108 = in147 & in19;
assign var109 = in146 & in18;
assign var110 = in145 & in17;
assign var111 = in144 & in16;
assign var112 = in143 & in15;
assign var113 = in142 & in14;
assign var114 = in141 & in13;
assign var115 = in140 & in12;
assign var116 = in139 & in11;
assign var117 = in138 & in10;
assign var118 = in137 & in9;
assign var119 = in136 & in8;
assign var120 = in135 & in7;
assign var121 = in134 & in6;
assign var122 = in133 & in5;
assign var123 = in132 & in4;
assign var124 = in131 & in3;
assign var125 = in130 & in2;
assign var126 = in129 & in1;
assign var127 = in128 & in0;
assign var128 = in255 ^ in127;
assign var129 = in254 ^ in126;
assign var130 = in253 ^ in125;
assign var131 = in252 ^ in124;
assign var132 = in251 ^ in123;
assign var133 = in250 ^ in122;
assign var134 = in249 ^ in121;
assign var135 = in248 ^ in120;
assign var136 = in247 ^ in119;
assign var137 = in246 ^ in118;
assign var138 = in245 ^ in117;
assign var139 = in244 ^ in116;
assign var140 = in243 ^ in115;
assign var141 = in242 ^ in114;
assign var142 = in241 ^ in113;
assign var143 = in240 ^ in112;
assign var144 = in239 ^ in111;
assign var145 = in238 ^ in110;
assign var146 = in237 ^ in109;
assign var147 = in236 ^ in108;
assign var148 = in235 ^ in107;
assign var149 = in234 ^ in106;
assign var150 = in233 ^ in105;
assign var151 = in232 ^ in104;
assign var152 = in231 ^ in103;
assign var153 = in230 ^ in102;
assign var154 = in229 ^ in101;
assign var155 = in228 ^ in100;
assign var156 = in227 ^ in99;
assign var157 = in226 ^ in98;
assign var158 = in225 ^ in97;
assign var159 = in224 ^ in96;
assign var160 = in223 ^ in95;
assign var161 = in222 ^ in94;
assign var162 = in221 ^ in93;
assign var163 = in220 ^ in92;
assign var164 = in219 ^ in91;
assign var165 = in218 ^ in90;
assign var166 = in217 ^ in89;
assign var167 = in216 ^ in88;
assign var168 = in215 ^ in87;
assign var169 = in214 ^ in86;
assign var170 = in213 ^ in85;
assign var171 = in212 ^ in84;
assign var172 = in211 ^ in83;
assign var173 = in210 ^ in82;
assign var174 = in209 ^ in81;
assign var175 = in208 ^ in80;
assign var176 = in207 ^ in79;
assign var177 = in206 ^ in78;
assign var178 = in205 ^ in77;
assign var179 = in204 ^ in76;
assign var180 = in203 ^ in75;
assign var181 = in202 ^ in74;
assign var182 = in201 ^ in73;
assign var183 = in200 ^ in72;
assign var184 = in199 ^ in71;
assign var185 = in198 ^ in70;
assign var186 = in197 ^ in69;
assign var187 = in196 ^ in68;
assign var188 = in195 ^ in67;
assign var189 = in194 ^ in66;
assign var190 = in193 ^ in65;
assign var191 = in192 ^ in64;
assign var192 = in191 ^ in63;
assign var193 = in190 ^ in62;
assign var194 = in189 ^ in61;
assign var195 = in188 ^ in60;
assign var196 = in187 ^ in59;
assign var197 = in186 ^ in58;
assign var198 = in185 ^ in57;
assign var199 = in184 ^ in56;
assign var200 = in183 ^ in55;
assign var201 = in182 ^ in54;
assign var202 = in181 ^ in53;
assign var203 = in180 ^ in52;
assign var204 = in179 ^ in51;
assign var205 = in178 ^ in50;
assign var206 = in177 ^ in49;
assign var207 = in176 ^ in48;
assign var208 = in175 ^ in47;
assign var209 = in174 ^ in46;
assign var210 = in173 ^ in45;
assign var211 = in172 ^ in44;
assign var212 = in171 ^ in43;
assign var213 = in170 ^ in42;
assign var214 = in169 ^ in41;
assign var215 = in168 ^ in40;
assign var216 = in167 ^ in39;
assign var217 = in166 ^ in38;
assign var218 = in165 ^ in37;
assign var219 = in164 ^ in36;
assign var220 = in163 ^ in35;
assign var221 = in162 ^ in34;
assign var222 = in161 ^ in33;
assign var223 = in160 ^ in32;
assign var224 = in159 ^ in31;
assign var225 = in158 ^ in30;
assign var226 = in157 ^ in29;
assign var227 = in156 ^ in28;
assign var228 = in155 ^ in27;
assign var229 = in154 ^ in26;
assign var230 = in153 ^ in25;
assign var231 = in152 ^ in24;
assign var232 = in151 ^ in23;
assign var233 = in150 ^ in22;
assign var234 = in149 ^ in21;
assign var235 = in148 ^ in20;
assign var236 = in147 ^ in19;
assign var237 = in146 ^ in18;
assign var238 = in145 ^ in17;
assign var239 = in144 ^ in16;
assign var240 = in143 ^ in15;
assign var241 = in142 ^ in14;
assign var242 = in141 ^ in13;
assign var243 = in140 ^ in12;
assign var244 = in139 ^ in11;
assign var245 = in138 ^ in10;
assign var246 = in137 ^ in9;
assign var247 = in136 ^ in8;
assign var248 = in135 ^ in7;
assign var249 = in134 ^ in6;
assign var250 = in133 ^ in5;
assign var251 = in132 ^ in4;
assign var252 = in131 ^ in3;
assign var253 = in130 ^ in2;
assign var254 = in129 ^ in1;
assign var255 = in128 ^ in0;
assign var256 = var255 & var126;
assign var257 = var127 | var256;
assign var258 = var255 & var254;
assign var259 = var253 & var124;
assign var260 = var125 | var259;
assign var261 = var253 & var252;
assign var262 = var251 & var122;
assign var263 = var123 | var262;
assign var264 = var251 & var250;
assign var265 = var249 & var120;
assign var266 = var121 | var265;
assign var267 = var249 & var248;
assign var268 = var247 & var118;
assign var269 = var119 | var268;
assign var270 = var247 & var246;
assign var271 = var245 & var116;
assign var272 = var117 | var271;
assign var273 = var245 & var244;
assign var274 = var243 & var114;
assign var275 = var115 | var274;
assign var276 = var243 & var242;
assign var277 = var241 & var112;
assign var278 = var113 | var277;
assign var279 = var241 & var240;
assign var280 = var239 & var110;
assign var281 = var111 | var280;
assign var282 = var239 & var238;
assign var283 = var237 & var108;
assign var284 = var109 | var283;
assign var285 = var237 & var236;
assign var286 = var235 & var106;
assign var287 = var107 | var286;
assign var288 = var235 & var234;
assign var289 = var233 & var104;
assign var290 = var105 | var289;
assign var291 = var233 & var232;
assign var292 = var231 & var102;
assign var293 = var103 | var292;
assign var294 = var231 & var230;
assign var295 = var229 & var100;
assign var296 = var101 | var295;
assign var297 = var229 & var228;
assign var298 = var227 & var98;
assign var299 = var99 | var298;
assign var300 = var227 & var226;
assign var301 = var225 & var96;
assign var302 = var97 | var301;
assign var303 = var225 & var224;
assign var304 = var223 & var94;
assign var305 = var95 | var304;
assign var306 = var223 & var222;
assign var307 = var221 & var92;
assign var308 = var93 | var307;
assign var309 = var221 & var220;
assign var310 = var219 & var90;
assign var311 = var91 | var310;
assign var312 = var219 & var218;
assign var313 = var217 & var88;
assign var314 = var89 | var313;
assign var315 = var217 & var216;
assign var316 = var215 & var86;
assign var317 = var87 | var316;
assign var318 = var215 & var214;
assign var319 = var213 & var84;
assign var320 = var85 | var319;
assign var321 = var213 & var212;
assign var322 = var211 & var82;
assign var323 = var83 | var322;
assign var324 = var211 & var210;
assign var325 = var209 & var80;
assign var326 = var81 | var325;
assign var327 = var209 & var208;
assign var328 = var207 & var78;
assign var329 = var79 | var328;
assign var330 = var207 & var206;
assign var331 = var205 & var76;
assign var332 = var77 | var331;
assign var333 = var205 & var204;
assign var334 = var203 & var74;
assign var335 = var75 | var334;
assign var336 = var203 & var202;
assign var337 = var201 & var72;
assign var338 = var73 | var337;
assign var339 = var201 & var200;
assign var340 = var199 & var70;
assign var341 = var71 | var340;
assign var342 = var199 & var198;
assign var343 = var197 & var68;
assign var344 = var69 | var343;
assign var345 = var197 & var196;
assign var346 = var195 & var66;
assign var347 = var67 | var346;
assign var348 = var195 & var194;
assign var349 = var193 & var64;
assign var350 = var65 | var349;
assign var351 = var193 & var192;
assign var352 = var191 & var62;
assign var353 = var63 | var352;
assign var354 = var191 & var190;
assign var355 = var189 & var60;
assign var356 = var61 | var355;
assign var357 = var189 & var188;
assign var358 = var187 & var58;
assign var359 = var59 | var358;
assign var360 = var187 & var186;
assign var361 = var185 & var56;
assign var362 = var57 | var361;
assign var363 = var185 & var184;
assign var364 = var183 & var54;
assign var365 = var55 | var364;
assign var366 = var183 & var182;
assign var367 = var181 & var52;
assign var368 = var53 | var367;
assign var369 = var181 & var180;
assign var370 = var179 & var50;
assign var371 = var51 | var370;
assign var372 = var179 & var178;
assign var373 = var177 & var48;
assign var374 = var49 | var373;
assign var375 = var177 & var176;
assign var376 = var175 & var46;
assign var377 = var47 | var376;
assign var378 = var175 & var174;
assign var379 = var173 & var44;
assign var380 = var45 | var379;
assign var381 = var173 & var172;
assign var382 = var171 & var42;
assign var383 = var43 | var382;
assign var384 = var171 & var170;
assign var385 = var169 & var40;
assign var386 = var41 | var385;
assign var387 = var169 & var168;
assign var388 = var167 & var38;
assign var389 = var39 | var388;
assign var390 = var167 & var166;
assign var391 = var165 & var36;
assign var392 = var37 | var391;
assign var393 = var165 & var164;
assign var394 = var163 & var34;
assign var395 = var35 | var394;
assign var396 = var163 & var162;
assign var397 = var161 & var32;
assign var398 = var33 | var397;
assign var399 = var161 & var160;
assign var400 = var159 & var30;
assign var401 = var31 | var400;
assign var402 = var159 & var158;
assign var403 = var157 & var28;
assign var404 = var29 | var403;
assign var405 = var157 & var156;
assign var406 = var155 & var26;
assign var407 = var27 | var406;
assign var408 = var155 & var154;
assign var409 = var153 & var24;
assign var410 = var25 | var409;
assign var411 = var153 & var152;
assign var412 = var151 & var22;
assign var413 = var23 | var412;
assign var414 = var151 & var150;
assign var415 = var149 & var20;
assign var416 = var21 | var415;
assign var417 = var149 & var148;
assign var418 = var147 & var18;
assign var419 = var19 | var418;
assign var420 = var147 & var146;
assign var421 = var145 & var16;
assign var422 = var17 | var421;
assign var423 = var145 & var144;
assign var424 = var143 & var14;
assign var425 = var15 | var424;
assign var426 = var143 & var142;
assign var427 = var141 & var12;
assign var428 = var13 | var427;
assign var429 = var141 & var140;
assign var430 = var139 & var10;
assign var431 = var11 | var430;
assign var432 = var139 & var138;
assign var433 = var137 & var8;
assign var434 = var9 | var433;
assign var435 = var137 & var136;
assign var436 = var135 & var6;
assign var437 = var7 | var436;
assign var438 = var135 & var134;
assign var439 = var133 & var4;
assign var440 = var5 | var439;
assign var441 = var133 & var132;
assign var442 = var131 & var2;
assign var443 = var3 | var442;
assign var444 = var131 & var130;
assign var445 = var129 & var0;
assign var446 = var1 | var445;
assign var447 = var258 & var260;
assign var448 = var257 | var447;
assign var449 = var258 & var261;
assign var450 = var254 & var260;
assign var451 = var126 | var450;
assign var452 = var254 & var261;
assign var453 = var264 & var266;
assign var454 = var263 | var453;
assign var455 = var264 & var267;
assign var456 = var250 & var266;
assign var457 = var122 | var456;
assign var458 = var250 & var267;
assign var459 = var270 & var272;
assign var460 = var269 | var459;
assign var461 = var270 & var273;
assign var462 = var246 & var272;
assign var463 = var118 | var462;
assign var464 = var246 & var273;
assign var465 = var276 & var278;
assign var466 = var275 | var465;
assign var467 = var276 & var279;
assign var468 = var242 & var278;
assign var469 = var114 | var468;
assign var470 = var242 & var279;
assign var471 = var282 & var284;
assign var472 = var281 | var471;
assign var473 = var282 & var285;
assign var474 = var238 & var284;
assign var475 = var110 | var474;
assign var476 = var238 & var285;
assign var477 = var288 & var290;
assign var478 = var287 | var477;
assign var479 = var288 & var291;
assign var480 = var234 & var290;
assign var481 = var106 | var480;
assign var482 = var234 & var291;
assign var483 = var294 & var296;
assign var484 = var293 | var483;
assign var485 = var294 & var297;
assign var486 = var230 & var296;
assign var487 = var102 | var486;
assign var488 = var230 & var297;
assign var489 = var300 & var302;
assign var490 = var299 | var489;
assign var491 = var300 & var303;
assign var492 = var226 & var302;
assign var493 = var98 | var492;
assign var494 = var226 & var303;
assign var495 = var306 & var308;
assign var496 = var305 | var495;
assign var497 = var306 & var309;
assign var498 = var222 & var308;
assign var499 = var94 | var498;
assign var500 = var222 & var309;
assign var501 = var312 & var314;
assign var502 = var311 | var501;
assign var503 = var312 & var315;
assign var504 = var218 & var314;
assign var505 = var90 | var504;
assign var506 = var218 & var315;
assign var507 = var318 & var320;
assign var508 = var317 | var507;
assign var509 = var318 & var321;
assign var510 = var214 & var320;
assign var511 = var86 | var510;
assign var512 = var214 & var321;
assign var513 = var324 & var326;
assign var514 = var323 | var513;
assign var515 = var324 & var327;
assign var516 = var210 & var326;
assign var517 = var82 | var516;
assign var518 = var210 & var327;
assign var519 = var330 & var332;
assign var520 = var329 | var519;
assign var521 = var330 & var333;
assign var522 = var206 & var332;
assign var523 = var78 | var522;
assign var524 = var206 & var333;
assign var525 = var336 & var338;
assign var526 = var335 | var525;
assign var527 = var336 & var339;
assign var528 = var202 & var338;
assign var529 = var74 | var528;
assign var530 = var202 & var339;
assign var531 = var342 & var344;
assign var532 = var341 | var531;
assign var533 = var342 & var345;
assign var534 = var198 & var344;
assign var535 = var70 | var534;
assign var536 = var198 & var345;
assign var537 = var348 & var350;
assign var538 = var347 | var537;
assign var539 = var348 & var351;
assign var540 = var194 & var350;
assign var541 = var66 | var540;
assign var542 = var194 & var351;
assign var543 = var354 & var356;
assign var544 = var353 | var543;
assign var545 = var354 & var357;
assign var546 = var190 & var356;
assign var547 = var62 | var546;
assign var548 = var190 & var357;
assign var549 = var360 & var362;
assign var550 = var359 | var549;
assign var551 = var360 & var363;
assign var552 = var186 & var362;
assign var553 = var58 | var552;
assign var554 = var186 & var363;
assign var555 = var366 & var368;
assign var556 = var365 | var555;
assign var557 = var366 & var369;
assign var558 = var182 & var368;
assign var559 = var54 | var558;
assign var560 = var182 & var369;
assign var561 = var372 & var374;
assign var562 = var371 | var561;
assign var563 = var372 & var375;
assign var564 = var178 & var374;
assign var565 = var50 | var564;
assign var566 = var178 & var375;
assign var567 = var378 & var380;
assign var568 = var377 | var567;
assign var569 = var378 & var381;
assign var570 = var174 & var380;
assign var571 = var46 | var570;
assign var572 = var174 & var381;
assign var573 = var384 & var386;
assign var574 = var383 | var573;
assign var575 = var384 & var387;
assign var576 = var170 & var386;
assign var577 = var42 | var576;
assign var578 = var170 & var387;
assign var579 = var390 & var392;
assign var580 = var389 | var579;
assign var581 = var390 & var393;
assign var582 = var166 & var392;
assign var583 = var38 | var582;
assign var584 = var166 & var393;
assign var585 = var396 & var398;
assign var586 = var395 | var585;
assign var587 = var396 & var399;
assign var588 = var162 & var398;
assign var589 = var34 | var588;
assign var590 = var162 & var399;
assign var591 = var402 & var404;
assign var592 = var401 | var591;
assign var593 = var402 & var405;
assign var594 = var158 & var404;
assign var595 = var30 | var594;
assign var596 = var158 & var405;
assign var597 = var408 & var410;
assign var598 = var407 | var597;
assign var599 = var408 & var411;
assign var600 = var154 & var410;
assign var601 = var26 | var600;
assign var602 = var154 & var411;
assign var603 = var414 & var416;
assign var604 = var413 | var603;
assign var605 = var414 & var417;
assign var606 = var150 & var416;
assign var607 = var22 | var606;
assign var608 = var150 & var417;
assign var609 = var420 & var422;
assign var610 = var419 | var609;
assign var611 = var420 & var423;
assign var612 = var146 & var422;
assign var613 = var18 | var612;
assign var614 = var146 & var423;
assign var615 = var426 & var428;
assign var616 = var425 | var615;
assign var617 = var426 & var429;
assign var618 = var142 & var428;
assign var619 = var14 | var618;
assign var620 = var142 & var429;
assign var621 = var432 & var434;
assign var622 = var431 | var621;
assign var623 = var432 & var435;
assign var624 = var138 & var434;
assign var625 = var10 | var624;
assign var626 = var138 & var435;
assign var627 = var438 & var440;
assign var628 = var437 | var627;
assign var629 = var438 & var441;
assign var630 = var134 & var440;
assign var631 = var6 | var630;
assign var632 = var134 & var441;
assign var633 = var444 & var446;
assign var634 = var443 | var633;
assign var635 = var130 & var446;
assign var636 = var2 | var635;
assign var637 = var449 & var454;
assign var638 = var448 | var637;
assign var639 = var449 & var455;
assign var640 = var452 & var454;
assign var641 = var451 | var640;
assign var642 = var452 & var455;
assign var643 = var261 & var454;
assign var644 = var260 | var643;
assign var645 = var261 & var455;
assign var646 = var252 & var454;
assign var647 = var124 | var646;
assign var648 = var252 & var455;
assign var649 = var461 & var466;
assign var650 = var460 | var649;
assign var651 = var461 & var467;
assign var652 = var464 & var466;
assign var653 = var463 | var652;
assign var654 = var464 & var467;
assign var655 = var273 & var466;
assign var656 = var272 | var655;
assign var657 = var273 & var467;
assign var658 = var244 & var466;
assign var659 = var116 | var658;
assign var660 = var244 & var467;
assign var661 = var473 & var478;
assign var662 = var472 | var661;
assign var663 = var473 & var479;
assign var664 = var476 & var478;
assign var665 = var475 | var664;
assign var666 = var476 & var479;
assign var667 = var285 & var478;
assign var668 = var284 | var667;
assign var669 = var285 & var479;
assign var670 = var236 & var478;
assign var671 = var108 | var670;
assign var672 = var236 & var479;
assign var673 = var485 & var490;
assign var674 = var484 | var673;
assign var675 = var485 & var491;
assign var676 = var488 & var490;
assign var677 = var487 | var676;
assign var678 = var488 & var491;
assign var679 = var297 & var490;
assign var680 = var296 | var679;
assign var681 = var297 & var491;
assign var682 = var228 & var490;
assign var683 = var100 | var682;
assign var684 = var228 & var491;
assign var685 = var497 & var502;
assign var686 = var496 | var685;
assign var687 = var497 & var503;
assign var688 = var500 & var502;
assign var689 = var499 | var688;
assign var690 = var500 & var503;
assign var691 = var309 & var502;
assign var692 = var308 | var691;
assign var693 = var309 & var503;
assign var694 = var220 & var502;
assign var695 = var92 | var694;
assign var696 = var220 & var503;
assign var697 = var509 & var514;
assign var698 = var508 | var697;
assign var699 = var509 & var515;
assign var700 = var512 & var514;
assign var701 = var511 | var700;
assign var702 = var512 & var515;
assign var703 = var321 & var514;
assign var704 = var320 | var703;
assign var705 = var321 & var515;
assign var706 = var212 & var514;
assign var707 = var84 | var706;
assign var708 = var212 & var515;
assign var709 = var521 & var526;
assign var710 = var520 | var709;
assign var711 = var521 & var527;
assign var712 = var524 & var526;
assign var713 = var523 | var712;
assign var714 = var524 & var527;
assign var715 = var333 & var526;
assign var716 = var332 | var715;
assign var717 = var333 & var527;
assign var718 = var204 & var526;
assign var719 = var76 | var718;
assign var720 = var204 & var527;
assign var721 = var533 & var538;
assign var722 = var532 | var721;
assign var723 = var533 & var539;
assign var724 = var536 & var538;
assign var725 = var535 | var724;
assign var726 = var536 & var539;
assign var727 = var345 & var538;
assign var728 = var344 | var727;
assign var729 = var345 & var539;
assign var730 = var196 & var538;
assign var731 = var68 | var730;
assign var732 = var196 & var539;
assign var733 = var545 & var550;
assign var734 = var544 | var733;
assign var735 = var545 & var551;
assign var736 = var548 & var550;
assign var737 = var547 | var736;
assign var738 = var548 & var551;
assign var739 = var357 & var550;
assign var740 = var356 | var739;
assign var741 = var357 & var551;
assign var742 = var188 & var550;
assign var743 = var60 | var742;
assign var744 = var188 & var551;
assign var745 = var557 & var562;
assign var746 = var556 | var745;
assign var747 = var557 & var563;
assign var748 = var560 & var562;
assign var749 = var559 | var748;
assign var750 = var560 & var563;
assign var751 = var369 & var562;
assign var752 = var368 | var751;
assign var753 = var369 & var563;
assign var754 = var180 & var562;
assign var755 = var52 | var754;
assign var756 = var180 & var563;
assign var757 = var569 & var574;
assign var758 = var568 | var757;
assign var759 = var569 & var575;
assign var760 = var572 & var574;
assign var761 = var571 | var760;
assign var762 = var572 & var575;
assign var763 = var381 & var574;
assign var764 = var380 | var763;
assign var765 = var381 & var575;
assign var766 = var172 & var574;
assign var767 = var44 | var766;
assign var768 = var172 & var575;
assign var769 = var581 & var586;
assign var770 = var580 | var769;
assign var771 = var581 & var587;
assign var772 = var584 & var586;
assign var773 = var583 | var772;
assign var774 = var584 & var587;
assign var775 = var393 & var586;
assign var776 = var392 | var775;
assign var777 = var393 & var587;
assign var778 = var164 & var586;
assign var779 = var36 | var778;
assign var780 = var164 & var587;
assign var781 = var593 & var598;
assign var782 = var592 | var781;
assign var783 = var593 & var599;
assign var784 = var596 & var598;
assign var785 = var595 | var784;
assign var786 = var596 & var599;
assign var787 = var405 & var598;
assign var788 = var404 | var787;
assign var789 = var405 & var599;
assign var790 = var156 & var598;
assign var791 = var28 | var790;
assign var792 = var156 & var599;
assign var793 = var605 & var610;
assign var794 = var604 | var793;
assign var795 = var605 & var611;
assign var796 = var608 & var610;
assign var797 = var607 | var796;
assign var798 = var608 & var611;
assign var799 = var417 & var610;
assign var800 = var416 | var799;
assign var801 = var417 & var611;
assign var802 = var148 & var610;
assign var803 = var20 | var802;
assign var804 = var148 & var611;
assign var805 = var617 & var622;
assign var806 = var616 | var805;
assign var807 = var617 & var623;
assign var808 = var620 & var622;
assign var809 = var619 | var808;
assign var810 = var620 & var623;
assign var811 = var429 & var622;
assign var812 = var428 | var811;
assign var813 = var429 & var623;
assign var814 = var140 & var622;
assign var815 = var12 | var814;
assign var816 = var140 & var623;
assign var817 = var629 & var634;
assign var818 = var628 | var817;
assign var819 = var632 & var634;
assign var820 = var631 | var819;
assign var821 = var441 & var634;
assign var822 = var440 | var821;
assign var823 = var132 & var634;
assign var824 = var4 | var823;
assign var825 = var639 & var650;
assign var826 = var638 | var825;
assign var827 = var639 & var651;
assign var828 = var642 & var650;
assign var829 = var641 | var828;
assign var830 = var642 & var651;
assign var831 = var645 & var650;
assign var832 = var644 | var831;
assign var833 = var645 & var651;
assign var834 = var648 & var650;
assign var835 = var647 | var834;
assign var836 = var648 & var651;
assign var837 = var455 & var650;
assign var838 = var454 | var837;
assign var839 = var455 & var651;
assign var840 = var458 & var650;
assign var841 = var457 | var840;
assign var842 = var458 & var651;
assign var843 = var267 & var650;
assign var844 = var266 | var843;
assign var845 = var267 & var651;
assign var846 = var248 & var650;
assign var847 = var120 | var846;
assign var848 = var248 & var651;
assign var849 = var663 & var674;
assign var850 = var662 | var849;
assign var851 = var663 & var675;
assign var852 = var666 & var674;
assign var853 = var665 | var852;
assign var854 = var666 & var675;
assign var855 = var669 & var674;
assign var856 = var668 | var855;
assign var857 = var669 & var675;
assign var858 = var672 & var674;
assign var859 = var671 | var858;
assign var860 = var672 & var675;
assign var861 = var479 & var674;
assign var862 = var478 | var861;
assign var863 = var479 & var675;
assign var864 = var482 & var674;
assign var865 = var481 | var864;
assign var866 = var482 & var675;
assign var867 = var291 & var674;
assign var868 = var290 | var867;
assign var869 = var291 & var675;
assign var870 = var232 & var674;
assign var871 = var104 | var870;
assign var872 = var232 & var675;
assign var873 = var687 & var698;
assign var874 = var686 | var873;
assign var875 = var687 & var699;
assign var876 = var690 & var698;
assign var877 = var689 | var876;
assign var878 = var690 & var699;
assign var879 = var693 & var698;
assign var880 = var692 | var879;
assign var881 = var693 & var699;
assign var882 = var696 & var698;
assign var883 = var695 | var882;
assign var884 = var696 & var699;
assign var885 = var503 & var698;
assign var886 = var502 | var885;
assign var887 = var503 & var699;
assign var888 = var506 & var698;
assign var889 = var505 | var888;
assign var890 = var506 & var699;
assign var891 = var315 & var698;
assign var892 = var314 | var891;
assign var893 = var315 & var699;
assign var894 = var216 & var698;
assign var895 = var88 | var894;
assign var896 = var216 & var699;
assign var897 = var711 & var722;
assign var898 = var710 | var897;
assign var899 = var711 & var723;
assign var900 = var714 & var722;
assign var901 = var713 | var900;
assign var902 = var714 & var723;
assign var903 = var717 & var722;
assign var904 = var716 | var903;
assign var905 = var717 & var723;
assign var906 = var720 & var722;
assign var907 = var719 | var906;
assign var908 = var720 & var723;
assign var909 = var527 & var722;
assign var910 = var526 | var909;
assign var911 = var527 & var723;
assign var912 = var530 & var722;
assign var913 = var529 | var912;
assign var914 = var530 & var723;
assign var915 = var339 & var722;
assign var916 = var338 | var915;
assign var917 = var339 & var723;
assign var918 = var200 & var722;
assign var919 = var72 | var918;
assign var920 = var200 & var723;
assign var921 = var735 & var746;
assign var922 = var734 | var921;
assign var923 = var735 & var747;
assign var924 = var738 & var746;
assign var925 = var737 | var924;
assign var926 = var738 & var747;
assign var927 = var741 & var746;
assign var928 = var740 | var927;
assign var929 = var741 & var747;
assign var930 = var744 & var746;
assign var931 = var743 | var930;
assign var932 = var744 & var747;
assign var933 = var551 & var746;
assign var934 = var550 | var933;
assign var935 = var551 & var747;
assign var936 = var554 & var746;
assign var937 = var553 | var936;
assign var938 = var554 & var747;
assign var939 = var363 & var746;
assign var940 = var362 | var939;
assign var941 = var363 & var747;
assign var942 = var184 & var746;
assign var943 = var56 | var942;
assign var944 = var184 & var747;
assign var945 = var759 & var770;
assign var946 = var758 | var945;
assign var947 = var759 & var771;
assign var948 = var762 & var770;
assign var949 = var761 | var948;
assign var950 = var762 & var771;
assign var951 = var765 & var770;
assign var952 = var764 | var951;
assign var953 = var765 & var771;
assign var954 = var768 & var770;
assign var955 = var767 | var954;
assign var956 = var768 & var771;
assign var957 = var575 & var770;
assign var958 = var574 | var957;
assign var959 = var575 & var771;
assign var960 = var578 & var770;
assign var961 = var577 | var960;
assign var962 = var578 & var771;
assign var963 = var387 & var770;
assign var964 = var386 | var963;
assign var965 = var387 & var771;
assign var966 = var168 & var770;
assign var967 = var40 | var966;
assign var968 = var168 & var771;
assign var969 = var783 & var794;
assign var970 = var782 | var969;
assign var971 = var783 & var795;
assign var972 = var786 & var794;
assign var973 = var785 | var972;
assign var974 = var786 & var795;
assign var975 = var789 & var794;
assign var976 = var788 | var975;
assign var977 = var789 & var795;
assign var978 = var792 & var794;
assign var979 = var791 | var978;
assign var980 = var792 & var795;
assign var981 = var599 & var794;
assign var982 = var598 | var981;
assign var983 = var599 & var795;
assign var984 = var602 & var794;
assign var985 = var601 | var984;
assign var986 = var602 & var795;
assign var987 = var411 & var794;
assign var988 = var410 | var987;
assign var989 = var411 & var795;
assign var990 = var152 & var794;
assign var991 = var24 | var990;
assign var992 = var152 & var795;
assign var993 = var807 & var818;
assign var994 = var806 | var993;
assign var995 = var810 & var818;
assign var996 = var809 | var995;
assign var997 = var813 & var818;
assign var998 = var812 | var997;
assign var999 = var816 & var818;
assign var1000 = var815 | var999;
assign var1001 = var623 & var818;
assign var1002 = var622 | var1001;
assign var1003 = var626 & var818;
assign var1004 = var625 | var1003;
assign var1005 = var435 & var818;
assign var1006 = var434 | var1005;
assign var1007 = var136 & var818;
assign var1008 = var8 | var1007;
assign var1009 = var827 & var850;
assign var1010 = var826 | var1009;
assign var1011 = var827 & var851;
assign var1012 = var830 & var850;
assign var1013 = var829 | var1012;
assign var1014 = var830 & var851;
assign var1015 = var833 & var850;
assign var1016 = var832 | var1015;
assign var1017 = var833 & var851;
assign var1018 = var836 & var850;
assign var1019 = var835 | var1018;
assign var1020 = var836 & var851;
assign var1021 = var839 & var850;
assign var1022 = var838 | var1021;
assign var1023 = var839 & var851;
assign var1024 = var842 & var850;
assign var1025 = var841 | var1024;
assign var1026 = var842 & var851;
assign var1027 = var845 & var850;
assign var1028 = var844 | var1027;
assign var1029 = var845 & var851;
assign var1030 = var848 & var850;
assign var1031 = var847 | var1030;
assign var1032 = var848 & var851;
assign var1033 = var651 & var850;
assign var1034 = var650 | var1033;
assign var1035 = var651 & var851;
assign var1036 = var654 & var850;
assign var1037 = var653 | var1036;
assign var1038 = var654 & var851;
assign var1039 = var657 & var850;
assign var1040 = var656 | var1039;
assign var1041 = var657 & var851;
assign var1042 = var660 & var850;
assign var1043 = var659 | var1042;
assign var1044 = var660 & var851;
assign var1045 = var467 & var850;
assign var1046 = var466 | var1045;
assign var1047 = var467 & var851;
assign var1048 = var470 & var850;
assign var1049 = var469 | var1048;
assign var1050 = var470 & var851;
assign var1051 = var279 & var850;
assign var1052 = var278 | var1051;
assign var1053 = var279 & var851;
assign var1054 = var240 & var850;
assign var1055 = var112 | var1054;
assign var1056 = var240 & var851;
assign var1057 = var875 & var898;
assign var1058 = var874 | var1057;
assign var1059 = var875 & var899;
assign var1060 = var878 & var898;
assign var1061 = var877 | var1060;
assign var1062 = var878 & var899;
assign var1063 = var881 & var898;
assign var1064 = var880 | var1063;
assign var1065 = var881 & var899;
assign var1066 = var884 & var898;
assign var1067 = var883 | var1066;
assign var1068 = var884 & var899;
assign var1069 = var887 & var898;
assign var1070 = var886 | var1069;
assign var1071 = var887 & var899;
assign var1072 = var890 & var898;
assign var1073 = var889 | var1072;
assign var1074 = var890 & var899;
assign var1075 = var893 & var898;
assign var1076 = var892 | var1075;
assign var1077 = var893 & var899;
assign var1078 = var896 & var898;
assign var1079 = var895 | var1078;
assign var1080 = var896 & var899;
assign var1081 = var699 & var898;
assign var1082 = var698 | var1081;
assign var1083 = var699 & var899;
assign var1084 = var702 & var898;
assign var1085 = var701 | var1084;
assign var1086 = var702 & var899;
assign var1087 = var705 & var898;
assign var1088 = var704 | var1087;
assign var1089 = var705 & var899;
assign var1090 = var708 & var898;
assign var1091 = var707 | var1090;
assign var1092 = var708 & var899;
assign var1093 = var515 & var898;
assign var1094 = var514 | var1093;
assign var1095 = var515 & var899;
assign var1096 = var518 & var898;
assign var1097 = var517 | var1096;
assign var1098 = var518 & var899;
assign var1099 = var327 & var898;
assign var1100 = var326 | var1099;
assign var1101 = var327 & var899;
assign var1102 = var208 & var898;
assign var1103 = var80 | var1102;
assign var1104 = var208 & var899;
assign var1105 = var923 & var946;
assign var1106 = var922 | var1105;
assign var1107 = var923 & var947;
assign var1108 = var926 & var946;
assign var1109 = var925 | var1108;
assign var1110 = var926 & var947;
assign var1111 = var929 & var946;
assign var1112 = var928 | var1111;
assign var1113 = var929 & var947;
assign var1114 = var932 & var946;
assign var1115 = var931 | var1114;
assign var1116 = var932 & var947;
assign var1117 = var935 & var946;
assign var1118 = var934 | var1117;
assign var1119 = var935 & var947;
assign var1120 = var938 & var946;
assign var1121 = var937 | var1120;
assign var1122 = var938 & var947;
assign var1123 = var941 & var946;
assign var1124 = var940 | var1123;
assign var1125 = var941 & var947;
assign var1126 = var944 & var946;
assign var1127 = var943 | var1126;
assign var1128 = var944 & var947;
assign var1129 = var747 & var946;
assign var1130 = var746 | var1129;
assign var1131 = var747 & var947;
assign var1132 = var750 & var946;
assign var1133 = var749 | var1132;
assign var1134 = var750 & var947;
assign var1135 = var753 & var946;
assign var1136 = var752 | var1135;
assign var1137 = var753 & var947;
assign var1138 = var756 & var946;
assign var1139 = var755 | var1138;
assign var1140 = var756 & var947;
assign var1141 = var563 & var946;
assign var1142 = var562 | var1141;
assign var1143 = var563 & var947;
assign var1144 = var566 & var946;
assign var1145 = var565 | var1144;
assign var1146 = var566 & var947;
assign var1147 = var375 & var946;
assign var1148 = var374 | var1147;
assign var1149 = var375 & var947;
assign var1150 = var176 & var946;
assign var1151 = var48 | var1150;
assign var1152 = var176 & var947;
assign var1153 = var971 & var994;
assign var1154 = var970 | var1153;
assign var1155 = var974 & var994;
assign var1156 = var973 | var1155;
assign var1157 = var977 & var994;
assign var1158 = var976 | var1157;
assign var1159 = var980 & var994;
assign var1160 = var979 | var1159;
assign var1161 = var983 & var994;
assign var1162 = var982 | var1161;
assign var1163 = var986 & var994;
assign var1164 = var985 | var1163;
assign var1165 = var989 & var994;
assign var1166 = var988 | var1165;
assign var1167 = var992 & var994;
assign var1168 = var991 | var1167;
assign var1169 = var795 & var994;
assign var1170 = var794 | var1169;
assign var1171 = var798 & var994;
assign var1172 = var797 | var1171;
assign var1173 = var801 & var994;
assign var1174 = var800 | var1173;
assign var1175 = var804 & var994;
assign var1176 = var803 | var1175;
assign var1177 = var611 & var994;
assign var1178 = var610 | var1177;
assign var1179 = var614 & var994;
assign var1180 = var613 | var1179;
assign var1181 = var423 & var994;
assign var1182 = var422 | var1181;
assign var1183 = var144 & var994;
assign var1184 = var16 | var1183;
assign var1185 = var1011 & var1058;
assign var1186 = var1010 | var1185;
assign var1187 = var1011 & var1059;
assign var1188 = var1014 & var1058;
assign var1189 = var1013 | var1188;
assign var1190 = var1014 & var1059;
assign var1191 = var1017 & var1058;
assign var1192 = var1016 | var1191;
assign var1193 = var1017 & var1059;
assign var1194 = var1020 & var1058;
assign var1195 = var1019 | var1194;
assign var1196 = var1020 & var1059;
assign var1197 = var1023 & var1058;
assign var1198 = var1022 | var1197;
assign var1199 = var1023 & var1059;
assign var1200 = var1026 & var1058;
assign var1201 = var1025 | var1200;
assign var1202 = var1026 & var1059;
assign var1203 = var1029 & var1058;
assign var1204 = var1028 | var1203;
assign var1205 = var1029 & var1059;
assign var1206 = var1032 & var1058;
assign var1207 = var1031 | var1206;
assign var1208 = var1032 & var1059;
assign var1209 = var1035 & var1058;
assign var1210 = var1034 | var1209;
assign var1211 = var1035 & var1059;
assign var1212 = var1038 & var1058;
assign var1213 = var1037 | var1212;
assign var1214 = var1038 & var1059;
assign var1215 = var1041 & var1058;
assign var1216 = var1040 | var1215;
assign var1217 = var1041 & var1059;
assign var1218 = var1044 & var1058;
assign var1219 = var1043 | var1218;
assign var1220 = var1044 & var1059;
assign var1221 = var1047 & var1058;
assign var1222 = var1046 | var1221;
assign var1223 = var1047 & var1059;
assign var1224 = var1050 & var1058;
assign var1225 = var1049 | var1224;
assign var1226 = var1050 & var1059;
assign var1227 = var1053 & var1058;
assign var1228 = var1052 | var1227;
assign var1229 = var1053 & var1059;
assign var1230 = var1056 & var1058;
assign var1231 = var1055 | var1230;
assign var1232 = var1056 & var1059;
assign var1233 = var851 & var1058;
assign var1234 = var850 | var1233;
assign var1235 = var851 & var1059;
assign var1236 = var854 & var1058;
assign var1237 = var853 | var1236;
assign var1238 = var854 & var1059;
assign var1239 = var857 & var1058;
assign var1240 = var856 | var1239;
assign var1241 = var857 & var1059;
assign var1242 = var860 & var1058;
assign var1243 = var859 | var1242;
assign var1244 = var860 & var1059;
assign var1245 = var863 & var1058;
assign var1246 = var862 | var1245;
assign var1247 = var863 & var1059;
assign var1248 = var866 & var1058;
assign var1249 = var865 | var1248;
assign var1250 = var866 & var1059;
assign var1251 = var869 & var1058;
assign var1252 = var868 | var1251;
assign var1253 = var869 & var1059;
assign var1254 = var872 & var1058;
assign var1255 = var871 | var1254;
assign var1256 = var872 & var1059;
assign var1257 = var675 & var1058;
assign var1258 = var674 | var1257;
assign var1259 = var675 & var1059;
assign var1260 = var678 & var1058;
assign var1261 = var677 | var1260;
assign var1262 = var678 & var1059;
assign var1263 = var681 & var1058;
assign var1264 = var680 | var1263;
assign var1265 = var681 & var1059;
assign var1266 = var684 & var1058;
assign var1267 = var683 | var1266;
assign var1268 = var684 & var1059;
assign var1269 = var491 & var1058;
assign var1270 = var490 | var1269;
assign var1271 = var491 & var1059;
assign var1272 = var494 & var1058;
assign var1273 = var493 | var1272;
assign var1274 = var494 & var1059;
assign var1275 = var303 & var1058;
assign var1276 = var302 | var1275;
assign var1277 = var303 & var1059;
assign var1278 = var224 & var1058;
assign var1279 = var96 | var1278;
assign var1280 = var224 & var1059;
assign var1281 = var1107 & var1154;
assign var1282 = var1106 | var1281;
assign var1283 = var1110 & var1154;
assign var1284 = var1109 | var1283;
assign var1285 = var1113 & var1154;
assign var1286 = var1112 | var1285;
assign var1287 = var1116 & var1154;
assign var1288 = var1115 | var1287;
assign var1289 = var1119 & var1154;
assign var1290 = var1118 | var1289;
assign var1291 = var1122 & var1154;
assign var1292 = var1121 | var1291;
assign var1293 = var1125 & var1154;
assign var1294 = var1124 | var1293;
assign var1295 = var1128 & var1154;
assign var1296 = var1127 | var1295;
assign var1297 = var1131 & var1154;
assign var1298 = var1130 | var1297;
assign var1299 = var1134 & var1154;
assign var1300 = var1133 | var1299;
assign var1301 = var1137 & var1154;
assign var1302 = var1136 | var1301;
assign var1303 = var1140 & var1154;
assign var1304 = var1139 | var1303;
assign var1305 = var1143 & var1154;
assign var1306 = var1142 | var1305;
assign var1307 = var1146 & var1154;
assign var1308 = var1145 | var1307;
assign var1309 = var1149 & var1154;
assign var1310 = var1148 | var1309;
assign var1311 = var1152 & var1154;
assign var1312 = var1151 | var1311;
assign var1313 = var947 & var1154;
assign var1314 = var946 | var1313;
assign var1315 = var950 & var1154;
assign var1316 = var949 | var1315;
assign var1317 = var953 & var1154;
assign var1318 = var952 | var1317;
assign var1319 = var956 & var1154;
assign var1320 = var955 | var1319;
assign var1321 = var959 & var1154;
assign var1322 = var958 | var1321;
assign var1323 = var962 & var1154;
assign var1324 = var961 | var1323;
assign var1325 = var965 & var1154;
assign var1326 = var964 | var1325;
assign var1327 = var968 & var1154;
assign var1328 = var967 | var1327;
assign var1329 = var771 & var1154;
assign var1330 = var770 | var1329;
assign var1331 = var774 & var1154;
assign var1332 = var773 | var1331;
assign var1333 = var777 & var1154;
assign var1334 = var776 | var1333;
assign var1335 = var780 & var1154;
assign var1336 = var779 | var1335;
assign var1337 = var587 & var1154;
assign var1338 = var586 | var1337;
assign var1339 = var590 & var1154;
assign var1340 = var589 | var1339;
assign var1341 = var399 & var1154;
assign var1342 = var398 | var1341;
assign var1343 = var160 & var1154;
assign var1344 = var32 | var1343;
assign var1345 = var1187 & var1282;
assign var1346 = var1186 | var1345;
assign var1347 = var1190 & var1282;
assign var1348 = var1189 | var1347;
assign var1349 = var1193 & var1282;
assign var1350 = var1192 | var1349;
assign var1351 = var1196 & var1282;
assign var1352 = var1195 | var1351;
assign var1353 = var1199 & var1282;
assign var1354 = var1198 | var1353;
assign var1355 = var1202 & var1282;
assign var1356 = var1201 | var1355;
assign var1357 = var1205 & var1282;
assign var1358 = var1204 | var1357;
assign var1359 = var1208 & var1282;
assign var1360 = var1207 | var1359;
assign var1361 = var1211 & var1282;
assign var1362 = var1210 | var1361;
assign var1363 = var1214 & var1282;
assign var1364 = var1213 | var1363;
assign var1365 = var1217 & var1282;
assign var1366 = var1216 | var1365;
assign var1367 = var1220 & var1282;
assign var1368 = var1219 | var1367;
assign var1369 = var1223 & var1282;
assign var1370 = var1222 | var1369;
assign var1371 = var1226 & var1282;
assign var1372 = var1225 | var1371;
assign var1373 = var1229 & var1282;
assign var1374 = var1228 | var1373;
assign var1375 = var1232 & var1282;
assign var1376 = var1231 | var1375;
assign var1377 = var1235 & var1282;
assign var1378 = var1234 | var1377;
assign var1379 = var1238 & var1282;
assign var1380 = var1237 | var1379;
assign var1381 = var1241 & var1282;
assign var1382 = var1240 | var1381;
assign var1383 = var1244 & var1282;
assign var1384 = var1243 | var1383;
assign var1385 = var1247 & var1282;
assign var1386 = var1246 | var1385;
assign var1387 = var1250 & var1282;
assign var1388 = var1249 | var1387;
assign var1389 = var1253 & var1282;
assign var1390 = var1252 | var1389;
assign var1391 = var1256 & var1282;
assign var1392 = var1255 | var1391;
assign var1393 = var1259 & var1282;
assign var1394 = var1258 | var1393;
assign var1395 = var1262 & var1282;
assign var1396 = var1261 | var1395;
assign var1397 = var1265 & var1282;
assign var1398 = var1264 | var1397;
assign var1399 = var1268 & var1282;
assign var1400 = var1267 | var1399;
assign var1401 = var1271 & var1282;
assign var1402 = var1270 | var1401;
assign var1403 = var1274 & var1282;
assign var1404 = var1273 | var1403;
assign var1405 = var1277 & var1282;
assign var1406 = var1276 | var1405;
assign var1407 = var1280 & var1282;
assign var1408 = var1279 | var1407;
assign var1409 = var1059 & var1282;
assign var1410 = var1058 | var1409;
assign var1411 = var1062 & var1282;
assign var1412 = var1061 | var1411;
assign var1413 = var1065 & var1282;
assign var1414 = var1064 | var1413;
assign var1415 = var1068 & var1282;
assign var1416 = var1067 | var1415;
assign var1417 = var1071 & var1282;
assign var1418 = var1070 | var1417;
assign var1419 = var1074 & var1282;
assign var1420 = var1073 | var1419;
assign var1421 = var1077 & var1282;
assign var1422 = var1076 | var1421;
assign var1423 = var1080 & var1282;
assign var1424 = var1079 | var1423;
assign var1425 = var1083 & var1282;
assign var1426 = var1082 | var1425;
assign var1427 = var1086 & var1282;
assign var1428 = var1085 | var1427;
assign var1429 = var1089 & var1282;
assign var1430 = var1088 | var1429;
assign var1431 = var1092 & var1282;
assign var1432 = var1091 | var1431;
assign var1433 = var1095 & var1282;
assign var1434 = var1094 | var1433;
assign var1435 = var1098 & var1282;
assign var1436 = var1097 | var1435;
assign var1437 = var1101 & var1282;
assign var1438 = var1100 | var1437;
assign var1439 = var1104 & var1282;
assign var1440 = var1103 | var1439;
assign var1441 = var899 & var1282;
assign var1442 = var898 | var1441;
assign var1443 = var902 & var1282;
assign var1444 = var901 | var1443;
assign var1445 = var905 & var1282;
assign var1446 = var904 | var1445;
assign var1447 = var908 & var1282;
assign var1448 = var907 | var1447;
assign var1449 = var911 & var1282;
assign var1450 = var910 | var1449;
assign var1451 = var914 & var1282;
assign var1452 = var913 | var1451;
assign var1453 = var917 & var1282;
assign var1454 = var916 | var1453;
assign var1455 = var920 & var1282;
assign var1456 = var919 | var1455;
assign var1457 = var723 & var1282;
assign var1458 = var722 | var1457;
assign var1459 = var726 & var1282;
assign var1460 = var725 | var1459;
assign var1461 = var729 & var1282;
assign var1462 = var728 | var1461;
assign var1463 = var732 & var1282;
assign var1464 = var731 | var1463;
assign var1465 = var539 & var1282;
assign var1466 = var538 | var1465;
assign var1467 = var542 & var1282;
assign var1468 = var541 | var1467;
assign var1469 = var351 & var1282;
assign var1470 = var350 | var1469;
assign var1471 = var192 & var1282;
assign var1472 = var64 | var1471;
assign var1473 = var129 ^ var0;
assign var1474 = var130 ^ var446;
assign var1475 = var131 ^ var636;
assign var1476 = var132 ^ var634;
assign var1477 = var133 ^ var824;
assign var1478 = var134 ^ var822;
assign var1479 = var135 ^ var820;
assign var1480 = var136 ^ var818;
assign var1481 = var137 ^ var1008;
assign var1482 = var138 ^ var1006;
assign var1483 = var139 ^ var1004;
assign var1484 = var140 ^ var1002;
assign var1485 = var141 ^ var1000;
assign var1486 = var142 ^ var998;
assign var1487 = var143 ^ var996;
assign var1488 = var144 ^ var994;
assign var1489 = var145 ^ var1184;
assign var1490 = var146 ^ var1182;
assign var1491 = var147 ^ var1180;
assign var1492 = var148 ^ var1178;
assign var1493 = var149 ^ var1176;
assign var1494 = var150 ^ var1174;
assign var1495 = var151 ^ var1172;
assign var1496 = var152 ^ var1170;
assign var1497 = var153 ^ var1168;
assign var1498 = var154 ^ var1166;
assign var1499 = var155 ^ var1164;
assign var1500 = var156 ^ var1162;
assign var1501 = var157 ^ var1160;
assign var1502 = var158 ^ var1158;
assign var1503 = var159 ^ var1156;
assign var1504 = var160 ^ var1154;
assign var1505 = var161 ^ var1344;
assign var1506 = var162 ^ var1342;
assign var1507 = var163 ^ var1340;
assign var1508 = var164 ^ var1338;
assign var1509 = var165 ^ var1336;
assign var1510 = var166 ^ var1334;
assign var1511 = var167 ^ var1332;
assign var1512 = var168 ^ var1330;
assign var1513 = var169 ^ var1328;
assign var1514 = var170 ^ var1326;
assign var1515 = var171 ^ var1324;
assign var1516 = var172 ^ var1322;
assign var1517 = var173 ^ var1320;
assign var1518 = var174 ^ var1318;
assign var1519 = var175 ^ var1316;
assign var1520 = var176 ^ var1314;
assign var1521 = var177 ^ var1312;
assign var1522 = var178 ^ var1310;
assign var1523 = var179 ^ var1308;
assign var1524 = var180 ^ var1306;
assign var1525 = var181 ^ var1304;
assign var1526 = var182 ^ var1302;
assign var1527 = var183 ^ var1300;
assign var1528 = var184 ^ var1298;
assign var1529 = var185 ^ var1296;
assign var1530 = var186 ^ var1294;
assign var1531 = var187 ^ var1292;
assign var1532 = var188 ^ var1290;
assign var1533 = var189 ^ var1288;
assign var1534 = var190 ^ var1286;
assign var1535 = var191 ^ var1284;
assign var1536 = var192 ^ var1282;
assign var1537 = var193 ^ var1472;
assign var1538 = var194 ^ var1470;
assign var1539 = var195 ^ var1468;
assign var1540 = var196 ^ var1466;
assign var1541 = var197 ^ var1464;
assign var1542 = var198 ^ var1462;
assign var1543 = var199 ^ var1460;
assign var1544 = var200 ^ var1458;
assign var1545 = var201 ^ var1456;
assign var1546 = var202 ^ var1454;
assign var1547 = var203 ^ var1452;
assign var1548 = var204 ^ var1450;
assign var1549 = var205 ^ var1448;
assign var1550 = var206 ^ var1446;
assign var1551 = var207 ^ var1444;
assign var1552 = var208 ^ var1442;
assign var1553 = var209 ^ var1440;
assign var1554 = var210 ^ var1438;
assign var1555 = var211 ^ var1436;
assign var1556 = var212 ^ var1434;
assign var1557 = var213 ^ var1432;
assign var1558 = var214 ^ var1430;
assign var1559 = var215 ^ var1428;
assign var1560 = var216 ^ var1426;
assign var1561 = var217 ^ var1424;
assign var1562 = var218 ^ var1422;
assign var1563 = var219 ^ var1420;
assign var1564 = var220 ^ var1418;
assign var1565 = var221 ^ var1416;
assign var1566 = var222 ^ var1414;
assign var1567 = var223 ^ var1412;
assign var1568 = var224 ^ var1410;
assign var1569 = var225 ^ var1408;
assign var1570 = var226 ^ var1406;
assign var1571 = var227 ^ var1404;
assign var1572 = var228 ^ var1402;
assign var1573 = var229 ^ var1400;
assign var1574 = var230 ^ var1398;
assign var1575 = var231 ^ var1396;
assign var1576 = var232 ^ var1394;
assign var1577 = var233 ^ var1392;
assign var1578 = var234 ^ var1390;
assign var1579 = var235 ^ var1388;
assign var1580 = var236 ^ var1386;
assign var1581 = var237 ^ var1384;
assign var1582 = var238 ^ var1382;
assign var1583 = var239 ^ var1380;
assign var1584 = var240 ^ var1378;
assign var1585 = var241 ^ var1376;
assign var1586 = var242 ^ var1374;
assign var1587 = var243 ^ var1372;
assign var1588 = var244 ^ var1370;
assign var1589 = var245 ^ var1368;
assign var1590 = var246 ^ var1366;
assign var1591 = var247 ^ var1364;
assign var1592 = var248 ^ var1362;
assign var1593 = var249 ^ var1360;
assign var1594 = var250 ^ var1358;
assign var1595 = var251 ^ var1356;
assign var1596 = var252 ^ var1354;
assign var1597 = var253 ^ var1352;
assign var1598 = var254 ^ var1350;
assign var1599 = var255 ^ var1348;
assign out0 = var1346;
assign out1 = var1599;
assign out2 = var1598;
assign out3 = var1597;
assign out4 = var1596;
assign out5 = var1595;
assign out6 = var1594;
assign out7 = var1593;
assign out8 = var1592;
assign out9 = var1591;
assign out10 = var1590;
assign out11 = var1589;
assign out12 = var1588;
assign out13 = var1587;
assign out14 = var1586;
assign out15 = var1585;
assign out16 = var1584;
assign out17 = var1583;
assign out18 = var1582;
assign out19 = var1581;
assign out20 = var1580;
assign out21 = var1579;
assign out22 = var1578;
assign out23 = var1577;
assign out24 = var1576;
assign out25 = var1575;
assign out26 = var1574;
assign out27 = var1573;
assign out28 = var1572;
assign out29 = var1571;
assign out30 = var1570;
assign out31 = var1569;
assign out32 = var1568;
assign out33 = var1567;
assign out34 = var1566;
assign out35 = var1565;
assign out36 = var1564;
assign out37 = var1563;
assign out38 = var1562;
assign out39 = var1561;
assign out40 = var1560;
assign out41 = var1559;
assign out42 = var1558;
assign out43 = var1557;
assign out44 = var1556;
assign out45 = var1555;
assign out46 = var1554;
assign out47 = var1553;
assign out48 = var1552;
assign out49 = var1551;
assign out50 = var1550;
assign out51 = var1549;
assign out52 = var1548;
assign out53 = var1547;
assign out54 = var1546;
assign out55 = var1545;
assign out56 = var1544;
assign out57 = var1543;
assign out58 = var1542;
assign out59 = var1541;
assign out60 = var1540;
assign out61 = var1539;
assign out62 = var1538;
assign out63 = var1537;
assign out64 = var1536;
assign out65 = var1535;
assign out66 = var1534;
assign out67 = var1533;
assign out68 = var1532;
assign out69 = var1531;
assign out70 = var1530;
assign out71 = var1529;
assign out72 = var1528;
assign out73 = var1527;
assign out74 = var1526;
assign out75 = var1525;
assign out76 = var1524;
assign out77 = var1523;
assign out78 = var1522;
assign out79 = var1521;
assign out80 = var1520;
assign out81 = var1519;
assign out82 = var1518;
assign out83 = var1517;
assign out84 = var1516;
assign out85 = var1515;
assign out86 = var1514;
assign out87 = var1513;
assign out88 = var1512;
assign out89 = var1511;
assign out90 = var1510;
assign out91 = var1509;
assign out92 = var1508;
assign out93 = var1507;
assign out94 = var1506;
assign out95 = var1505;
assign out96 = var1504;
assign out97 = var1503;
assign out98 = var1502;
assign out99 = var1501;
assign out100 = var1500;
assign out101 = var1499;
assign out102 = var1498;
assign out103 = var1497;
assign out104 = var1496;
assign out105 = var1495;
assign out106 = var1494;
assign out107 = var1493;
assign out108 = var1492;
assign out109 = var1491;
assign out110 = var1490;
assign out111 = var1489;
assign out112 = var1488;
assign out113 = var1487;
assign out114 = var1486;
assign out115 = var1485;
assign out116 = var1484;
assign out117 = var1483;
assign out118 = var1482;
assign out119 = var1481;
assign out120 = var1480;
assign out121 = var1479;
assign out122 = var1478;
assign out123 = var1477;
assign out124 = var1476;
assign out125 = var1475;
assign out126 = var1474;
assign out127 = var1473;
assign out128 = var128;
endmodule 
