module bk4 (in0, in1, in2, in3, in4, in5, in6, in7, out0, out1, out2, out3, out4, );
input in0;
input in1;
input in2;
input in3;
input in4;
input in5;
input in6;
input in7;
output out0;
output out1;
output out2;
output out3;
output out4;
wire var0;
wire var1;
wire var2;
wire var3;
wire var4;
wire var5;
wire var6;
wire var7;
wire var8;
wire var9;
wire var10;
wire var11;
wire var12;
wire var13;
wire var14;
wire var15;
wire var16;
wire var17;
wire var18;
wire var19;
wire var20;
assign var0 = in7 & in3;
assign var1 = in6 & in2;
assign var2 = in5 & in1;
assign var3 = in4 & in0;
assign var4 = in7 ^ in3;
assign var5 = in6 ^ in2;
assign var6 = in5 ^ in1;
assign var7 = in4 ^ in0;
assign var8 = var7 & var2;
assign var9 = var3 | var8;
assign var10 = var7 & var6;
assign var11 = var5 & var0;
assign var12 = var1 | var11;
assign var13 = var10 & var12;
assign var14 = var9 | var13;
assign var15 = var6 & var12;
assign var16 = var2 | var15;
assign var17 = var6 & var5;
assign var18 = var5 ^ var0;
assign var19 = var6 ^ var12;
assign var20 = var7 ^ var16;
assign out0 = var14;
assign out1 = var20;
assign out2 = var19;
assign out3 = var18;
assign out4 = var4;
endmodule 
