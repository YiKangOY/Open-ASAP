// Verilog
// c5315
// Ninputs 178
// Noutputs 123
// NtotalGates 2307
// BUFF1 313
// AND2 319
// NOT1 581
// NAND2 454
// AND4 27
// OR2 95
// AND3 359
// OR3 50
// OR4 61
// NOR2 19
// AND5 11
// OR5 8
// NOR3 6
// NOR4 2
// AND9 2

module c5315 (N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, 
              N27, N31, N34, N37, N40, N43, N46, N49, N52, N53, 
              N54, N61, N64, N67, N70, N73, N76, N79, N80, N81, 
              N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, 
              N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, 
              N120, N121, N122, N123, N126, N127, N128, N129, N130, N131, 
              N132, N135, N136, N137, N140, N141, N145, N146, N149, N152, 
              N155, N158, N161, N164, N167, N170, N173, N176, N179, N182, 
              N185, N188, N191, N194, N197, N200, N203, N206, N209, N210, 
              N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, 
              N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, 
              N289, N292, N293, N299, N302, N307, N308, N315, N316, N323, 
              N324, N331, N332, N335, N338, N341, N348, N351, N358, N361, 
              N366, N369, N372, N373, N374, N386, N389, N400, N411, N422, 
              N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, 
              N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, 
              N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, 
              N603, N607, N610, N613, N616, N619, N625, N631, N709, N816, 
              N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, 
              N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060, N2061, N2139, 
              N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357, N3358, N3359, 
              N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737, N4738, N4739, 
              N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716, N6877, N6924, 
              N6925, N6926, N6927, N7015, N7363, N7365, N7432, N7449, N7465, N7466, 
              N7467, N7469, N7470, N7471, N7472, N7473, N7474, N7476, N7503, N7504, 
              N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520, N7521, N7522, 
              N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, N7626, N7698, 
              N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706, N7707, N7735, 
              N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754, N7755, N7756, 
              N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123, N8124, N8127, 
              N8128);

input N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, 
      N27, N31, N34, N37, N40, N43, N46, N49, N52, N53, 
      N54, N61, N64, N67, N70, N73, N76, N79, N80, N81, 
      N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, 
      N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, 
      N120, N121, N122, N123, N126, N127, N128, N129, N130, N131, 
      N132, N135, N136, N137, N140, N141, N145, N146, N149, N152, 
      N155, N158, N161, N164, N167, N170, N173, N176, N179, N182, 
      N185, N188, N191, N194, N197, N200, N203, N206, N209, N210, 
      N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, 
      N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, 
      N289, N292, N293, N299, N302, N307, N308, N315, N316, N323, 
      N324, N331, N332, N335, N338, N341, N348, N351, N358, N361, 
      N366, N369, N372, N373, N374, N386, N389, N400, N411, N422, 
      N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, 
      N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, 
      N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, 
      N603, N607, N610, N613, N616, N619, N625, N631;

output N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143, 
       N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060, 
       N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357, 
       N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737, 
       N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716, 
       N6877, N6924, N6925, N6926, N6927, N7015, N7363, N7365, N7432, N7449, 
       N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474, N7476, 
       N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520, 
       N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, 
       N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706, 
       N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754, 
       N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123, 
       N8124, N8127, N8128;

wire N1042, N1043, N1067, N1080, N1092, N1104, N1146, N1148, N1149, N1150, 
     N1151, N1156, N1157, N1161, N1173, N1185, N1197, N1209, N1213, N1216, 
     N1219, N1223, N1235, N1247, N1259, N1271, N1280, N1292, N1303, N1315, 
     N1327, N1339, N1351, N1363, N1375, N1378, N1381, N1384, N1387, N1390, 
     N1393, N1396, N1415, N1418, N1421, N1424, N1427, N1430, N1433, N1436, 
     N1455, N1462, N1469, N1475, N1479, N1482, N1492, N1495, N1498, N1501, 
     N1504, N1507, N1510, N1513, N1516, N1519, N1522, N1525, N1542, N1545, 
     N1548, N1551, N1554, N1557, N1560, N1563, N1566, N1573, N1580, N1583, 
     N1588, N1594, N1597, N1600, N1603, N1606, N1609, N1612, N1615, N1618, 
     N1621, N1624, N1627, N1630, N1633, N1636, N1639, N1642, N1645, N1648, 
     N1651, N1654, N1657, N1660, N1663, N1675, N1685, N1697, N1709, N1721, 
     N1727, N1731, N1743, N1755, N1758, N1761, N1769, N1777, N1785, N1793, 
     N1800, N1807, N1814, N1821, N1824, N1827, N1830, N1833, N1836, N1839, 
     N1842, N1845, N1848, N1851, N1854, N1857, N1860, N1863, N1866, N1869, 
     N1872, N1875, N1878, N1881, N1884, N1887, N1890, N1893, N1896, N1899, 
     N1902, N1905, N1908, N1911, N1914, N1917, N1920, N1923, N1926, N1929, 
     N1932, N1935, N1938, N1941, N1944, N1947, N1950, N1953, N1956, N1959, 
     N1962, N1965, N1968, N2349, N2350, N2585, N2586, N2587, N2588, N2589, 
     N2591, N2592, N2593, N2594, N2595, N2596, N2597, N2598, N2599, N2600, 
     N2601, N2602, N2603, N2604, N2605, N2606, N2607, N2608, N2609, N2610, 
     N2611, N2612, N2613, N2614, N2615, N2616, N2617, N2618, N2619, N2620, 
     N2621, N2622, N2624, N2625, N2626, N2627, N2628, N2629, N2630, N2631, 
     N2632, N2633, N2634, N2635, N2636, N2637, N2638, N2639, N2640, N2641, 
     N2642, N2643, N2644, N2645, N2646, N2647, N2653, N2664, N2675, N2681, 
     N2692, N2703, N2704, N2709, N2710, N2711, N2712, N2713, N2714, N2715, 
     N2716, N2717, N2718, N2719, N2720, N2721, N2722, N2728, N2739, N2750, 
     N2756, N2767, N2778, N2779, N2790, N2801, N2812, N2823, N2824, N2825, 
     N2826, N2827, N2828, N2829, N2830, N2831, N2832, N2833, N2834, N2835, 
     N2836, N2837, N2838, N2839, N2840, N2841, N2842, N2843, N2844, N2845, 
     N2846, N2847, N2848, N2849, N2850, N2851, N2852, N2853, N2854, N2855, 
     N2861, N2867, N2868, N2869, N2870, N2871, N2872, N2873, N2874, N2875, 
     N2876, N2877, N2882, N2891, N2901, N2902, N2903, N2904, N2905, N2906, 
     N2907, N2908, N2909, N2910, N2911, N2912, N2913, N2914, N2915, N2916, 
     N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925, N2926, 
     N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, N2936, 
     N2937, N2938, N2939, N2940, N2941, N2942, N2948, N2954, N2955, N2956, 
     N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964, N2969, N2970, 
     N2971, N2972, N2973, N2974, N2975, N2976, N2977, N2978, N2979, N2980, 
     N2981, N2982, N2983, N2984, N2985, N2986, N2987, N2988, N2989, N2990, 
     N2991, N2992, N2993, N2994, N2995, N2996, N2997, N2998, N2999, N3000, 
     N3003, N3006, N3007, N3010, N3013, N3014, N3015, N3016, N3017, N3018, 
     N3019, N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028, 
     N3029, N3030, N3031, N3032, N3033, N3034, N3035, N3038, N3041, N3052, 
     N3063, N3068, N3071, N3072, N3073, N3074, N3075, N3086, N3097, N3108, 
     N3119, N3130, N3141, N3142, N3143, N3144, N3145, N3146, N3147, N3158, 
     N3169, N3180, N3191, N3194, N3195, N3196, N3197, N3198, N3199, N3200, 
     N3203, N3401, N3402, N3403, N3404, N3405, N3406, N3407, N3408, N3409, 
     N3410, N3411, N3412, N3413, N3414, N3415, N3416, N3444, N3445, N3446, 
     N3447, N3448, N3449, N3450, N3451, N3452, N3453, N3454, N3455, N3456, 
     N3459, N3460, N3461, N3462, N3463, N3464, N3465, N3466, N3481, N3482, 
     N3483, N3484, N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492, 
     N3493, N3502, N3503, N3504, N3505, N3506, N3507, N3508, N3509, N3510, 
     N3511, N3512, N3513, N3514, N3515, N3558, N3559, N3560, N3561, N3562, 
     N3563, N3605, N3606, N3607, N3608, N3609, N3610, N3614, N3615, N3616, 
     N3617, N3618, N3619, N3620, N3621, N3622, N3623, N3624, N3625, N3626, 
     N3627, N3628, N3629, N3630, N3631, N3632, N3633, N3634, N3635, N3636, 
     N3637, N3638, N3639, N3640, N3641, N3642, N3643, N3644, N3645, N3646, 
     N3647, N3648, N3649, N3650, N3651, N3652, N3653, N3654, N3655, N3656, 
     N3657, N3658, N3659, N3660, N3661, N3662, N3663, N3664, N3665, N3666, 
     N3667, N3668, N3669, N3670, N3671, N3672, N3673, N3674, N3675, N3676, 
     N3677, N3678, N3679, N3680, N3681, N3682, N3683, N3684, N3685, N3686, 
     N3687, N3688, N3689, N3691, N3700, N3701, N3702, N3703, N3704, N3705, 
     N3708, N3709, N3710, N3711, N3712, N3713, N3715, N3716, N3717, N3718, 
     N3719, N3720, N3721, N3722, N3723, N3724, N3725, N3726, N3727, N3728, 
     N3729, N3730, N3731, N3732, N3738, N3739, N3740, N3741, N3742, N3743, 
     N3744, N3745, N3746, N3747, N3748, N3749, N3750, N3751, N3752, N3753, 
     N3754, N3755, N3756, N3757, N3758, N3759, N3760, N3761, N3762, N3763, 
     N3764, N3765, N3766, N3767, N3768, N3769, N3770, N3771, N3775, N3779, 
     N3780, N3781, N3782, N3783, N3784, N3785, N3786, N3787, N3788, N3789, 
     N3793, N3797, N3800, N3801, N3802, N3803, N3804, N3805, N3806, N3807, 
     N3808, N3809, N3810, N3813, N3816, N3819, N3822, N3823, N3824, N3827, 
     N3828, N3829, N3830, N3831, N3834, N3835, N3836, N3837, N3838, N3839, 
     N3840, N3841, N3842, N3849, N3855, N3861, N3867, N3873, N3881, N3887, 
     N3893, N3908, N3909, N3911, N3914, N3915, N3916, N3917, N3918, N3919, 
     N3920, N3921, N3927, N3933, N3942, N3948, N3956, N3962, N3968, N3975, 
     N3976, N3977, N3978, N3979, N3980, N3981, N3982, N3983, N3984, N3987, 
     N3988, N3989, N3990, N3991, N3998, N4008, N4011, N4021, N4024, N4027, 
     N4031, N4032, N4033, N4034, N4035, N4036, N4037, N4038, N4039, N4040, 
     N4041, N4042, N4067, N4080, N4088, N4091, N4094, N4097, N4100, N4103, 
     N4106, N4109, N4144, N4147, N4150, N4153, N4156, N4159, N4183, N4184, 
     N4185, N4186, N4188, N4191, N4196, N4197, N4198, N4199, N4200, N4203, 
     N4206, N4209, N4212, N4215, N4219, N4223, N4224, N4225, N4228, N4231, 
     N4234, N4237, N4240, N4243, N4246, N4249, N4252, N4255, N4258, N4263, 
     N4264, N4267, N4268, N4269, N4270, N4271, N4273, N4274, N4276, N4277, 
     N4280, N4284, N4290, N4297, N4298, N4301, N4305, N4310, N4316, N4320, 
     N4325, N4331, N4332, N4336, N4342, N4349, N4357, N4364, N4375, N4379, 
     N4385, N4392, N4396, N4400, N4405, N4412, N4418, N4425, N4436, N4440, 
     N4445, N4451, N4456, N4462, N4469, N4477, N4512, N4515, N4516, N4521, 
     N4523, N4524, N4532, N4547, N4548, N4551, N4554, N4557, N4560, N4563, 
     N4566, N4569, N4572, N4575, N4578, N4581, N4584, N4587, N4590, N4593, 
     N4596, N4599, N4602, N4605, N4608, N4611, N4614, N4617, N4621, N4624, 
     N4627, N4630, N4633, N4637, N4640, N4643, N4646, N4649, N4652, N4655, 
     N4658, N4662, N4665, N4668, N4671, N4674, N4677, N4680, N4683, N4686, 
     N4689, N4692, N4695, N4698, N4701, N4702, N4720, N4721, N4724, N4725, 
     N4726, N4727, N4728, N4729, N4730, N4731, N4732, N4733, N4734, N4735, 
     N4736, N4741, N4855, N4856, N4908, N4909, N4939, N4942, N4947, N4953, 
     N4954, N4955, N4956, N4957, N4958, N4959, N4960, N4961, N4965, N4966, 
     N4967, N4968, N4972, N4973, N4974, N4975, N4976, N4977, N4978, N4979, 
     N4980, N4981, N4982, N4983, N4984, N4985, N4986, N4987, N5049, N5052, 
     N5053, N5054, N5055, N5056, N5057, N5058, N5059, N5060, N5061, N5062, 
     N5063, N5065, N5066, N5067, N5068, N5069, N5070, N5071, N5072, N5073, 
     N5074, N5075, N5076, N5077, N5078, N5079, N5080, N5081, N5082, N5083, 
     N5084, N5085, N5086, N5087, N5088, N5089, N5090, N5091, N5092, N5093, 
     N5094, N5095, N5096, N5097, N5098, N5099, N5100, N5101, N5102, N5103, 
     N5104, N5105, N5106, N5107, N5108, N5109, N5110, N5111, N5112, N5113, 
     N5114, N5115, N5116, N5117, N5118, N5119, N5120, N5121, N5122, N5123, 
     N5124, N5125, N5126, N5127, N5128, N5129, N5130, N5131, N5132, N5133, 
     N5135, N5136, N5137, N5138, N5139, N5140, N5141, N5142, N5143, N5144, 
     N5145, N5146, N5147, N5148, N5150, N5153, N5154, N5155, N5156, N5157, 
     N5160, N5161, N5162, N5163, N5164, N5165, N5166, N5169, N5172, N5173, 
     N5176, N5177, N5180, N5183, N5186, N5189, N5192, N5195, N5198, N5199, 
     N5202, N5205, N5208, N5211, N5214, N5217, N5220, N5223, N5224, N5225, 
     N5226, N5227, N5228, N5229, N5230, N5232, N5233, N5234, N5235, N5236, 
     N5239, N5241, N5242, N5243, N5244, N5245, N5246, N5247, N5248, N5249, 
     N5250, N5252, N5253, N5254, N5255, N5256, N5257, N5258, N5259, N5260, 
     N5261, N5262, N5263, N5264, N5274, N5275, N5282, N5283, N5284, N5298, 
     N5299, N5300, N5303, N5304, N5305, N5306, N5307, N5308, N5309, N5310, 
     N5311, N5312, N5315, N5319, N5324, N5328, N5331, N5332, N5346, N5363, 
     N5364, N5365, N5366, N5367, N5368, N5369, N5370, N5371, N5374, N5377, 
     N5382, N5385, N5389, N5396, N5407, N5418, N5424, N5431, N5441, N5452, 
     N5462, N5469, N5470, N5477, N5488, N5498, N5506, N5520, N5536, N5549, 
     N5555, N5562, N5573, N5579, N5595, N5606, N5616, N5617, N5618, N5619, 
     N5620, N5621, N5622, N5624, N5634, N5655, N5671, N5684, N5690, N5691, 
     N5692, N5696, N5700, N5703, N5707, N5711, N5726, N5727, N5728, N5730, 
     N5731, N5732, N5733, N5734, N5735, N5736, N5739, N5742, N5745, N5755, 
     N5756, N5954, N5955, N5956, N6005, N6006, N6023, N6024, N6025, N6028, 
     N6031, N6034, N6037, N6040, N6044, N6045, N6048, N6051, N6054, N6065, 
     N6066, N6067, N6068, N6069, N6071, N6072, N6073, N6074, N6075, N6076, 
     N6077, N6078, N6079, N6080, N6083, N6084, N6085, N6086, N6087, N6088, 
     N6089, N6090, N6091, N6094, N6095, N6096, N6097, N6098, N6099, N6100, 
     N6101, N6102, N6103, N6104, N6105, N6106, N6107, N6108, N6111, N6112, 
     N6113, N6114, N6115, N6116, N6117, N6120, N6121, N6122, N6123, N6124, 
     N6125, N6126, N6127, N6128, N6129, N6130, N6131, N6132, N6133, N6134, 
     N6135, N6136, N6137, N6138, N6139, N6140, N6143, N6144, N6145, N6146, 
     N6147, N6148, N6149, N6152, N6153, N6154, N6155, N6156, N6157, N6158, 
     N6159, N6160, N6161, N6162, N6163, N6164, N6168, N6171, N6172, N6173, 
     N6174, N6175, N6178, N6179, N6180, N6181, N6182, N6183, N6184, N6185, 
     N6186, N6187, N6188, N6189, N6190, N6191, N6192, N6193, N6194, N6197, 
     N6200, N6203, N6206, N6209, N6212, N6215, N6218, N6221, N6234, N6235, 
     N6238, N6241, N6244, N6247, N6250, N6253, N6256, N6259, N6262, N6265, 
     N6268, N6271, N6274, N6277, N6280, N6283, N6286, N6289, N6292, N6295, 
     N6298, N6301, N6304, N6307, N6310, N6313, N6316, N6319, N6322, N6325, 
     N6328, N6331, N6335, N6338, N6341, N6344, N6347, N6350, N6353, N6356, 
     N6359, N6364, N6367, N6370, N6373, N6374, N6375, N6376, N6377, N6378, 
     N6382, N6386, N6388, N6392, N6397, N6411, N6415, N6419, N6427, N6434, 
     N6437, N6441, N6445, N6448, N6449, N6466, N6469, N6470, N6471, N6472, 
     N6473, N6474, N6475, N6476, N6477, N6478, N6482, N6486, N6490, N6494, 
     N6500, N6504, N6508, N6512, N6516, N6526, N6536, N6539, N6553, N6556, 
     N6566, N6569, N6572, N6575, N6580, N6584, N6587, N6592, N6599, N6606, 
     N6609, N6619, N6622, N6630, N6631, N6632, N6633, N6634, N6637, N6640, 
     N6650, N6651, N6653, N6655, N6657, N6659, N6660, N6661, N6662, N6663, 
     N6664, N6666, N6668, N6670, N6672, N6675, N6680, N6681, N6682, N6683, 
     N6689, N6690, N6691, N6692, N6693, N6695, N6698, N6699, N6700, N6703, 
     N6708, N6709, N6710, N6711, N6712, N6713, N6714, N6715, N6718, N6719, 
     N6720, N6721, N6722, N6724, N6739, N6740, N6741, N6744, N6745, N6746, 
     N6751, N6752, N6753, N6754, N6755, N6760, N6761, N6762, N6772, N6773, 
     N6776, N6777, N6782, N6783, N6784, N6785, N6790, N6791, N6792, N6795, 
     N6801, N6802, N6803, N6804, N6805, N6806, N6807, N6808, N6809, N6810, 
     N6811, N6812, N6813, N6814, N6815, N6816, N6817, N6823, N6824, N6825, 
     N6826, N6827, N6828, N6829, N6830, N6831, N6834, N6835, N6836, N6837, 
     N6838, N6839, N6840, N6841, N6842, N6843, N6844, N6850, N6851, N6852, 
     N6853, N6854, N6855, N6856, N6857, N6860, N6861, N6862, N6863, N6866, 
     N6872, N6873, N6874, N6875, N6876, N6879, N6880, N6881, N6884, N6885, 
     N6888, N6889, N6890, N6891, N6894, N6895, N6896, N6897, N6900, N6901, 
     N6904, N6905, N6908, N6909, N6912, N6913, N6914, N6915, N6916, N6919, 
     N6922, N6923, N6930, N6932, N6935, N6936, N6937, N6938, N6939, N6940, 
     N6946, N6947, N6948, N6949, N6953, N6954, N6955, N6956, N6957, N6958, 
     N6964, N6965, N6966, N6967, N6973, N6974, N6975, N6976, N6977, N6978, 
     N6979, N6987, N6990, N6999, N7002, N7003, N7006, N7011, N7012, N7013, 
     N7016, N7018, N7019, N7020, N7021, N7022, N7023, N7028, N7031, N7034, 
     N7037, N7040, N7041, N7044, N7045, N7046, N7047, N7048, N7049, N7054, 
     N7057, N7060, N7064, N7065, N7072, N7073, N7074, N7075, N7076, N7079, 
     N7080, N7083, N7084, N7085, N7086, N7087, N7088, N7089, N7090, N7093, 
     N7094, N7097, N7101, N7105, N7110, N7114, N7115, N7116, N7125, N7126, 
     N7127, N7130, N7131, N7139, N7140, N7141, N7146, N7147, N7149, N7150, 
     N7151, N7152, N7153, N7158, N7159, N7160, N7166, N7167, N7168, N7169, 
     N7170, N7171, N7172, N7173, N7174, N7175, N7176, N7177, N7178, N7179, 
     N7180, N7181, N7182, N7183, N7184, N7185, N7186, N7187, N7188, N7189, 
     N7190, N7196, N7197, N7198, N7204, N7205, N7206, N7207, N7208, N7209, 
     N7212, N7215, N7216, N7217, N7218, N7219, N7222, N7225, N7228, N7229, 
     N7236, N7239, N7242, N7245, N7250, N7257, N7260, N7263, N7268, N7269, 
     N7270, N7276, N7282, N7288, N7294, N7300, N7301, N7304, N7310, N7320, 
     N7321, N7328, N7338, N7339, N7340, N7341, N7342, N7349, N7357, N7364, 
     N7394, N7397, N7402, N7405, N7406, N7407, N7408, N7409, N7412, N7415, 
     N7416, N7417, N7418, N7419, N7420, N7421, N7424, N7425, N7426, N7427, 
     N7428, N7429, N7430, N7431, N7433, N7434, N7435, N7436, N7437, N7438, 
     N7439, N7440, N7441, N7442, N7443, N7444, N7445, N7446, N7447, N7448, 
     N7450, N7451, N7452, N7453, N7454, N7455, N7456, N7457, N7458, N7459, 
     N7460, N7461, N7462, N7463, N7464, N7468, N7479, N7481, N7482, N7483, 
     N7484, N7485, N7486, N7487, N7488, N7489, N7492, N7493, N7498, N7499, 
     N7500, N7505, N7507, N7508, N7509, N7510, N7512, N7513, N7514, N7525, 
     N7526, N7527, N7528, N7529, N7530, N7531, N7537, N7543, N7549, N7555, 
     N7561, N7567, N7573, N7579, N7582, N7585, N7586, N7587, N7588, N7589, 
     N7592, N7595, N7598, N7599, N7624, N7625, N7631, N7636, N7657, N7658, 
     N7665, N7666, N7667, N7668, N7669, N7670, N7671, N7672, N7673, N7674, 
     N7675, N7676, N7677, N7678, N7679, N7680, N7681, N7682, N7683, N7684, 
     N7685, N7686, N7687, N7688, N7689, N7690, N7691, N7692, N7693, N7694, 
     N7695, N7696, N7697, N7708, N7709, N7710, N7711, N7712, N7715, N7718, 
     N7719, N7720, N7721, N7722, N7723, N7724, N7727, N7728, N7729, N7730, 
     N7731, N7732, N7733, N7734, N7743, N7744, N7749, N7750, N7751, N7762, 
     N7765, N7768, N7769, N7770, N7771, N7772, N7775, N7778, N7781, N7782, 
     N7787, N7788, N7795, N7796, N7797, N7798, N7799, N7800, N7803, N7806, 
     N7807, N7808, N7809, N7810, N7811, N7812, N7815, N7816, N7821, N7822, 
     N7823, N7826, N7829, N7832, N7833, N7834, N7835, N7836, N7839, N7842, 
     N7845, N7846, N7851, N7852, N7859, N7860, N7861, N7862, N7863, N7864, 
     N7867, N7870, N7871, N7872, N7873, N7874, N7875, N7876, N7879, N7880, 
     N7885, N7886, N7887, N7890, N7893, N7896, N7897, N7898, N7899, N7900, 
     N7903, N7906, N7909, N7910, N7917, N7918, N7923, N7924, N7925, N7926, 
     N7927, N7928, N7929, N7930, N7931, N7932, N7935, N7938, N7939, N7940, 
     N7943, N7944, N7945, N7946, N7951, N7954, N7957, N7960, N7963, N7966, 
     N7967, N7968, N7969, N7970, N7973, N7974, N7984, N7985, N7987, N7988, 
     N7989, N7990, N7991, N7992, N7993, N7994, N7995, N7996, N7997, N7998, 
     N8001, N8004, N8009, N8013, N8017, N8020, N8021, N8022, N8023, N8025, 
     N8026, N8027, N8031, N8032, N8033, N8034, N8035, N8036, N8037, N8038, 
     N8039, N8040, N8041, N8042, N8043, N8044, N8045, N8048, N8055, N8056, 
     N8057, N8058, N8059, N8060, N8061, N8064, N8071, N8072, N8073, N8074, 
     N8077, N8078, N8079, N8082, N8089, N8090, N8091, N8092, N8093, N8096, 
     N8099, N8102, N8113, N8114, N8115, N8116, N8117, N8118, N8119, N8120, 
     N8121, N8122, N8125, N8126;

buf BUFF1_1 (N709,  N141);
buf BUFF1_2 (N816,  N293);
and AND2_3 (N1042,  N135,  N631);
not NOT1_4 (N1043,  N591);
buf BUFF1_5 (N1066,  N592);
not NOT1_6 (N1067,  N595);
not NOT1_7 (N1080,  N596);
not NOT1_8 (N1092,  N597);
not NOT1_9 (N1104,  N598);
not NOT1_10 (N1137,  N545);
not NOT1_11 (N1138,  N348);
not NOT1_12 (N1139,  N366);
and AND2_13 (N1140,  N552,  N562);
not NOT1_14 (N1141,  N549);
not NOT1_15 (N1142,  N545);
not NOT1_16 (N1143,  N545);
not NOT1_17 (N1144,  N338);
not NOT1_18 (N1145,  N358);
nand NAND2_19 (N1146,  N373,  N1);
and AND2_20 (N1147,  N141,  N145);
not NOT1_21 (N1148,  N592);
not NOT1_22 (N1149,  N1042);
and AND2_23 (N1150,  N1043,  N27);
and AND2_24 (N1151,  N386,  N556);
not NOT1_25 (N1152,  N245);
not NOT1_26 (N1153,  N552);
not NOT1_27 (N1154,  N562);
not NOT1_28 (N1155,  N559);
and AND4_29 (N1156,  N386,  N559,  N556,  N552);
not NOT1_30 (N1157,  N566);
buf BUFF1_31 (N1161,  N571);
buf BUFF1_32 (N1173,  N574);
buf BUFF1_33 (N1185,  N571);
buf BUFF1_34 (N1197,  N574);
buf BUFF1_35 (N1209,  N137);
buf BUFF1_36 (N1213,  N137);
buf BUFF1_37 (N1216,  N141);
not NOT1_38 (N1219,  N583);
buf BUFF1_39 (N1223,  N577);
buf BUFF1_40 (N1235,  N580);
buf BUFF1_41 (N1247,  N577);
buf BUFF1_42 (N1259,  N580);
buf BUFF1_43 (N1271,  N254);
buf BUFF1_44 (N1280,  N251);
buf BUFF1_45 (N1292,  N251);
buf BUFF1_46 (N1303,  N248);
buf BUFF1_47 (N1315,  N248);
buf BUFF1_48 (N1327,  N610);
buf BUFF1_49 (N1339,  N607);
buf BUFF1_50 (N1351,  N613);
buf BUFF1_51 (N1363,  N616);
buf BUFF1_52 (N1375,  N210);
buf BUFF1_53 (N1378,  N210);
buf BUFF1_54 (N1381,  N218);
buf BUFF1_55 (N1384,  N218);
buf BUFF1_56 (N1387,  N226);
buf BUFF1_57 (N1390,  N226);
buf BUFF1_58 (N1393,  N234);
buf BUFF1_59 (N1396,  N234);
buf BUFF1_60 (N1415,  N257);
buf BUFF1_61 (N1418,  N257);
buf BUFF1_62 (N1421,  N265);
buf BUFF1_63 (N1424,  N265);
buf BUFF1_64 (N1427,  N273);
buf BUFF1_65 (N1430,  N273);
buf BUFF1_66 (N1433,  N281);
buf BUFF1_67 (N1436,  N281);
buf BUFF1_68 (N1455,  N335);
buf BUFF1_69 (N1462,  N335);
buf BUFF1_70 (N1469,  N206);
and AND2_71 (N1475,  N27,  N31);
buf BUFF1_72 (N1479,  N1);
buf BUFF1_73 (N1482,  N588);
buf BUFF1_74 (N1492,  N293);
buf BUFF1_75 (N1495,  N302);
buf BUFF1_76 (N1498,  N308);
buf BUFF1_77 (N1501,  N308);
buf BUFF1_78 (N1504,  N316);
buf BUFF1_79 (N1507,  N316);
buf BUFF1_80 (N1510,  N324);
buf BUFF1_81 (N1513,  N324);
buf BUFF1_82 (N1516,  N341);
buf BUFF1_83 (N1519,  N341);
buf BUFF1_84 (N1522,  N351);
buf BUFF1_85 (N1525,  N351);
buf BUFF1_86 (N1542,  N257);
buf BUFF1_87 (N1545,  N257);
buf BUFF1_88 (N1548,  N265);
buf BUFF1_89 (N1551,  N265);
buf BUFF1_90 (N1554,  N273);
buf BUFF1_91 (N1557,  N273);
buf BUFF1_92 (N1560,  N281);
buf BUFF1_93 (N1563,  N281);
buf BUFF1_94 (N1566,  N332);
buf BUFF1_95 (N1573,  N332);
buf BUFF1_96 (N1580,  N549);
and AND2_97 (N1583,  N31,  N27);
not NOT1_98 (N1588,  N588);
buf BUFF1_99 (N1594,  N324);
buf BUFF1_100 (N1597,  N324);
buf BUFF1_101 (N1600,  N341);
buf BUFF1_102 (N1603,  N341);
buf BUFF1_103 (N1606,  N351);
buf BUFF1_104 (N1609,  N351);
buf BUFF1_105 (N1612,  N293);
buf BUFF1_106 (N1615,  N302);
buf BUFF1_107 (N1618,  N308);
buf BUFF1_108 (N1621,  N308);
buf BUFF1_109 (N1624,  N316);
buf BUFF1_110 (N1627,  N316);
buf BUFF1_111 (N1630,  N361);
buf BUFF1_112 (N1633,  N361);
buf BUFF1_113 (N1636,  N210);
buf BUFF1_114 (N1639,  N210);
buf BUFF1_115 (N1642,  N218);
buf BUFF1_116 (N1645,  N218);
buf BUFF1_117 (N1648,  N226);
buf BUFF1_118 (N1651,  N226);
buf BUFF1_119 (N1654,  N234);
buf BUFF1_120 (N1657,  N234);
not NOT1_121 (N1660,  N324);
buf BUFF1_122 (N1663,  N242);
buf BUFF1_123 (N1675,  N242);
buf BUFF1_124 (N1685,  N254);
buf BUFF1_125 (N1697,  N610);
buf BUFF1_126 (N1709,  N607);
buf BUFF1_127 (N1721,  N625);
buf BUFF1_128 (N1727,  N619);
buf BUFF1_129 (N1731,  N613);
buf BUFF1_130 (N1743,  N616);
not NOT1_131 (N1755,  N599);
not NOT1_132 (N1758,  N603);
buf BUFF1_133 (N1761,  N619);
buf BUFF1_134 (N1769,  N625);
buf BUFF1_135 (N1777,  N619);
buf BUFF1_136 (N1785,  N625);
buf BUFF1_137 (N1793,  N619);
buf BUFF1_138 (N1800,  N625);
buf BUFF1_139 (N1807,  N619);
buf BUFF1_140 (N1814,  N625);
buf BUFF1_141 (N1821,  N299);
buf BUFF1_142 (N1824,  N446);
buf BUFF1_143 (N1827,  N457);
buf BUFF1_144 (N1830,  N468);
buf BUFF1_145 (N1833,  N422);
buf BUFF1_146 (N1836,  N435);
buf BUFF1_147 (N1839,  N389);
buf BUFF1_148 (N1842,  N400);
buf BUFF1_149 (N1845,  N411);
buf BUFF1_150 (N1848,  N374);
buf BUFF1_151 (N1851,  N4);
buf BUFF1_152 (N1854,  N446);
buf BUFF1_153 (N1857,  N457);
buf BUFF1_154 (N1860,  N468);
buf BUFF1_155 (N1863,  N435);
buf BUFF1_156 (N1866,  N389);
buf BUFF1_157 (N1869,  N400);
buf BUFF1_158 (N1872,  N411);
buf BUFF1_159 (N1875,  N422);
buf BUFF1_160 (N1878,  N374);
buf BUFF1_161 (N1881,  N479);
buf BUFF1_162 (N1884,  N490);
buf BUFF1_163 (N1887,  N503);
buf BUFF1_164 (N1890,  N514);
buf BUFF1_165 (N1893,  N523);
buf BUFF1_166 (N1896,  N534);
buf BUFF1_167 (N1899,  N54);
buf BUFF1_168 (N1902,  N479);
buf BUFF1_169 (N1905,  N503);
buf BUFF1_170 (N1908,  N514);
buf BUFF1_171 (N1911,  N523);
buf BUFF1_172 (N1914,  N534);
buf BUFF1_173 (N1917,  N490);
buf BUFF1_174 (N1920,  N361);
buf BUFF1_175 (N1923,  N369);
buf BUFF1_176 (N1926,  N341);
buf BUFF1_177 (N1929,  N351);
buf BUFF1_178 (N1932,  N308);
buf BUFF1_179 (N1935,  N316);
buf BUFF1_180 (N1938,  N293);
buf BUFF1_181 (N1941,  N302);
buf BUFF1_182 (N1944,  N281);
buf BUFF1_183 (N1947,  N289);
buf BUFF1_184 (N1950,  N265);
buf BUFF1_185 (N1953,  N273);
buf BUFF1_186 (N1956,  N234);
buf BUFF1_187 (N1959,  N257);
buf BUFF1_188 (N1962,  N218);
buf BUFF1_189 (N1965,  N226);
buf BUFF1_190 (N1968,  N210);
not NOT1_191 (N1972,  N1146);
and AND2_192 (N2054,  N136,  N1148);
not NOT1_193 (N2060,  N1150);
not NOT1_194 (N2061,  N1151);
buf BUFF1_195 (N2139,  N1209);
buf BUFF1_196 (N2142,  N1216);
buf BUFF1_197 (N2309,  N1479);
and AND2_198 (N2349,  N1104,  N514);
or OR2_199 (N2350,  N1067,  N514);
buf BUFF1_200 (N2387,  N1580);
buf BUFF1_201 (N2527,  N1821);
not NOT1_202 (N2584,  N1580);
and AND3_203 (N2585,  N170,  N1161,  N1173);
and AND3_204 (N2586,  N173,  N1161,  N1173);
and AND3_205 (N2587,  N167,  N1161,  N1173);
and AND3_206 (N2588,  N164,  N1161,  N1173);
and AND3_207 (N2589,  N161,  N1161,  N1173);
nand NAND2_208 (N2590,  N1475,  N140);
and AND3_209 (N2591,  N185,  N1185,  N1197);
and AND3_210 (N2592,  N158,  N1185,  N1197);
and AND3_211 (N2593,  N152,  N1185,  N1197);
and AND3_212 (N2594,  N146,  N1185,  N1197);
and AND3_213 (N2595,  N170,  N1223,  N1235);
and AND3_214 (N2596,  N173,  N1223,  N1235);
and AND3_215 (N2597,  N167,  N1223,  N1235);
and AND3_216 (N2598,  N164,  N1223,  N1235);
and AND3_217 (N2599,  N161,  N1223,  N1235);
and AND3_218 (N2600,  N185,  N1247,  N1259);
and AND3_219 (N2601,  N158,  N1247,  N1259);
and AND3_220 (N2602,  N152,  N1247,  N1259);
and AND3_221 (N2603,  N146,  N1247,  N1259);
and AND3_222 (N2604,  N106,  N1731,  N1743);
and AND3_223 (N2605,  N61,  N1327,  N1339);
and AND3_224 (N2606,  N106,  N1697,  N1709);
and AND3_225 (N2607,  N49,  N1697,  N1709);
and AND3_226 (N2608,  N103,  N1697,  N1709);
and AND3_227 (N2609,  N40,  N1697,  N1709);
and AND3_228 (N2610,  N37,  N1697,  N1709);
and AND3_229 (N2611,  N20,  N1327,  N1339);
and AND3_230 (N2612,  N17,  N1327,  N1339);
and AND3_231 (N2613,  N70,  N1327,  N1339);
and AND3_232 (N2614,  N64,  N1327,  N1339);
and AND3_233 (N2615,  N49,  N1731,  N1743);
and AND3_234 (N2616,  N103,  N1731,  N1743);
and AND3_235 (N2617,  N40,  N1731,  N1743);
and AND3_236 (N2618,  N37,  N1731,  N1743);
and AND3_237 (N2619,  N20,  N1351,  N1363);
and AND3_238 (N2620,  N17,  N1351,  N1363);
and AND3_239 (N2621,  N70,  N1351,  N1363);
and AND3_240 (N2622,  N64,  N1351,  N1363);
not NOT1_241 (N2623,  N1475);
and AND3_242 (N2624,  N123,  N1758,  N599);
and AND2_243 (N2625,  N1777,  N1785);
and AND3_244 (N2626,  N61,  N1351,  N1363);
and AND2_245 (N2627,  N1761,  N1769);
not NOT1_246 (N2628,  N1824);
not NOT1_247 (N2629,  N1827);
not NOT1_248 (N2630,  N1830);
not NOT1_249 (N2631,  N1833);
not NOT1_250 (N2632,  N1836);
not NOT1_251 (N2633,  N1839);
not NOT1_252 (N2634,  N1842);
not NOT1_253 (N2635,  N1845);
not NOT1_254 (N2636,  N1848);
not NOT1_255 (N2637,  N1851);
not NOT1_256 (N2638,  N1854);
not NOT1_257 (N2639,  N1857);
not NOT1_258 (N2640,  N1860);
not NOT1_259 (N2641,  N1863);
not NOT1_260 (N2642,  N1866);
not NOT1_261 (N2643,  N1869);
not NOT1_262 (N2644,  N1872);
not NOT1_263 (N2645,  N1875);
not NOT1_264 (N2646,  N1878);
buf BUFF1_265 (N2647,  N1209);
not NOT1_266 (N2653,  N1161);
not NOT1_267 (N2664,  N1173);
buf BUFF1_268 (N2675,  N1209);
not NOT1_269 (N2681,  N1185);
not NOT1_270 (N2692,  N1197);
and AND3_271 (N2703,  N179,  N1185,  N1197);
buf BUFF1_272 (N2704,  N1479);
not NOT1_273 (N2709,  N1881);
not NOT1_274 (N2710,  N1884);
not NOT1_275 (N2711,  N1887);
not NOT1_276 (N2712,  N1890);
not NOT1_277 (N2713,  N1893);
not NOT1_278 (N2714,  N1896);
not NOT1_279 (N2715,  N1899);
not NOT1_280 (N2716,  N1902);
not NOT1_281 (N2717,  N1905);
not NOT1_282 (N2718,  N1908);
not NOT1_283 (N2719,  N1911);
not NOT1_284 (N2720,  N1914);
not NOT1_285 (N2721,  N1917);
buf BUFF1_286 (N2722,  N1213);
not NOT1_287 (N2728,  N1223);
not NOT1_288 (N2739,  N1235);
buf BUFF1_289 (N2750,  N1213);
not NOT1_290 (N2756,  N1247);
not NOT1_291 (N2767,  N1259);
and AND3_292 (N2778,  N179,  N1247,  N1259);
not NOT1_293 (N2779,  N1327);
not NOT1_294 (N2790,  N1339);
not NOT1_295 (N2801,  N1351);
not NOT1_296 (N2812,  N1363);
not NOT1_297 (N2823,  N1375);
not NOT1_298 (N2824,  N1378);
not NOT1_299 (N2825,  N1381);
not NOT1_300 (N2826,  N1384);
not NOT1_301 (N2827,  N1387);
not NOT1_302 (N2828,  N1390);
not NOT1_303 (N2829,  N1393);
not NOT1_304 (N2830,  N1396);
and AND3_305 (N2831,  N1104,  N457,  N1378);
and AND3_306 (N2832,  N1104,  N468,  N1384);
and AND3_307 (N2833,  N1104,  N422,  N1390);
and AND3_308 (N2834,  N1104,  N435,  N1396);
and AND2_309 (N2835,  N1067,  N1375);
and AND2_310 (N2836,  N1067,  N1381);
and AND2_311 (N2837,  N1067,  N1387);
and AND2_312 (N2838,  N1067,  N1393);
not NOT1_313 (N2839,  N1415);
not NOT1_314 (N2840,  N1418);
not NOT1_315 (N2841,  N1421);
not NOT1_316 (N2842,  N1424);
not NOT1_317 (N2843,  N1427);
not NOT1_318 (N2844,  N1430);
not NOT1_319 (N2845,  N1433);
not NOT1_320 (N2846,  N1436);
and AND3_321 (N2847,  N1104,  N389,  N1418);
and AND3_322 (N2848,  N1104,  N400,  N1424);
and AND3_323 (N2849,  N1104,  N411,  N1430);
and AND3_324 (N2850,  N1104,  N374,  N1436);
and AND2_325 (N2851,  N1067,  N1415);
and AND2_326 (N2852,  N1067,  N1421);
and AND2_327 (N2853,  N1067,  N1427);
and AND2_328 (N2854,  N1067,  N1433);
not NOT1_329 (N2855,  N1455);
not NOT1_330 (N2861,  N1462);
and AND2_331 (N2867,  N292,  N1455);
and AND2_332 (N2868,  N288,  N1455);
and AND2_333 (N2869,  N280,  N1455);
and AND2_334 (N2870,  N272,  N1455);
and AND2_335 (N2871,  N264,  N1455);
and AND2_336 (N2872,  N241,  N1462);
and AND2_337 (N2873,  N233,  N1462);
and AND2_338 (N2874,  N225,  N1462);
and AND2_339 (N2875,  N217,  N1462);
and AND2_340 (N2876,  N209,  N1462);
buf BUFF1_341 (N2877,  N1216);
not NOT1_342 (N2882,  N1482);
not NOT1_343 (N2891,  N1475);
not NOT1_344 (N2901,  N1492);
not NOT1_345 (N2902,  N1495);
not NOT1_346 (N2903,  N1498);
not NOT1_347 (N2904,  N1501);
not NOT1_348 (N2905,  N1504);
not NOT1_349 (N2906,  N1507);
and AND2_350 (N2907,  N1303,  N1495);
and AND3_351 (N2908,  N1303,  N479,  N1501);
and AND3_352 (N2909,  N1303,  N490,  N1507);
and AND2_353 (N2910,  N1663,  N1492);
and AND2_354 (N2911,  N1663,  N1498);
and AND2_355 (N2912,  N1663,  N1504);
not NOT1_356 (N2913,  N1510);
not NOT1_357 (N2914,  N1513);
not NOT1_358 (N2915,  N1516);
not NOT1_359 (N2916,  N1519);
not NOT1_360 (N2917,  N1522);
not NOT1_361 (N2918,  N1525);
and AND3_362 (N2919,  N1104,  N503,  N1513);
not NOT1_363 (N2920,  N2349);
and AND3_364 (N2921,  N1104,  N523,  N1519);
and AND3_365 (N2922,  N1104,  N534,  N1525);
and AND2_366 (N2923,  N1067,  N1510);
and AND2_367 (N2924,  N1067,  N1516);
and AND2_368 (N2925,  N1067,  N1522);
not NOT1_369 (N2926,  N1542);
not NOT1_370 (N2927,  N1545);
not NOT1_371 (N2928,  N1548);
not NOT1_372 (N2929,  N1551);
not NOT1_373 (N2930,  N1554);
not NOT1_374 (N2931,  N1557);
not NOT1_375 (N2932,  N1560);
not NOT1_376 (N2933,  N1563);
and AND3_377 (N2934,  N1303,  N389,  N1545);
and AND3_378 (N2935,  N1303,  N400,  N1551);
and AND3_379 (N2936,  N1303,  N411,  N1557);
and AND3_380 (N2937,  N1303,  N374,  N1563);
and AND2_381 (N2938,  N1663,  N1542);
and AND2_382 (N2939,  N1663,  N1548);
and AND2_383 (N2940,  N1663,  N1554);
and AND2_384 (N2941,  N1663,  N1560);
not NOT1_385 (N2942,  N1566);
not NOT1_386 (N2948,  N1573);
and AND2_387 (N2954,  N372,  N1566);
and AND2_388 (N2955,  N366,  N1566);
and AND2_389 (N2956,  N358,  N1566);
and AND2_390 (N2957,  N348,  N1566);
and AND2_391 (N2958,  N338,  N1566);
and AND2_392 (N2959,  N331,  N1573);
and AND2_393 (N2960,  N323,  N1573);
and AND2_394 (N2961,  N315,  N1573);
and AND2_395 (N2962,  N307,  N1573);
and AND2_396 (N2963,  N299,  N1573);
not NOT1_397 (N2964,  N1588);
and AND2_398 (N2969,  N83,  N1588);
and AND2_399 (N2970,  N86,  N1588);
and AND2_400 (N2971,  N88,  N1588);
and AND2_401 (N2972,  N88,  N1588);
not NOT1_402 (N2973,  N1594);
not NOT1_403 (N2974,  N1597);
not NOT1_404 (N2975,  N1600);
not NOT1_405 (N2976,  N1603);
not NOT1_406 (N2977,  N1606);
not NOT1_407 (N2978,  N1609);
and AND3_408 (N2979,  N1315,  N503,  N1597);
and AND2_409 (N2980,  N1315,  N514);
and AND3_410 (N2981,  N1315,  N523,  N1603);
and AND3_411 (N2982,  N1315,  N534,  N1609);
and AND2_412 (N2983,  N1675,  N1594);
or OR2_413 (N2984,  N1675,  N514);
and AND2_414 (N2985,  N1675,  N1600);
and AND2_415 (N2986,  N1675,  N1606);
not NOT1_416 (N2987,  N1612);
not NOT1_417 (N2988,  N1615);
not NOT1_418 (N2989,  N1618);
not NOT1_419 (N2990,  N1621);
not NOT1_420 (N2991,  N1624);
not NOT1_421 (N2992,  N1627);
and AND2_422 (N2993,  N1315,  N1615);
and AND3_423 (N2994,  N1315,  N479,  N1621);
and AND3_424 (N2995,  N1315,  N490,  N1627);
and AND2_425 (N2996,  N1675,  N1612);
and AND2_426 (N2997,  N1675,  N1618);
and AND2_427 (N2998,  N1675,  N1624);
not NOT1_428 (N2999,  N1630);
buf BUFF1_429 (N3000,  N1469);
buf BUFF1_430 (N3003,  N1469);
not NOT1_431 (N3006,  N1633);
buf BUFF1_432 (N3007,  N1469);
buf BUFF1_433 (N3010,  N1469);
and AND2_434 (N3013,  N1315,  N1630);
and AND2_435 (N3014,  N1315,  N1633);
not NOT1_436 (N3015,  N1636);
not NOT1_437 (N3016,  N1639);
not NOT1_438 (N3017,  N1642);
not NOT1_439 (N3018,  N1645);
not NOT1_440 (N3019,  N1648);
not NOT1_441 (N3020,  N1651);
not NOT1_442 (N3021,  N1654);
not NOT1_443 (N3022,  N1657);
and AND3_444 (N3023,  N1303,  N457,  N1639);
and AND3_445 (N3024,  N1303,  N468,  N1645);
and AND3_446 (N3025,  N1303,  N422,  N1651);
and AND3_447 (N3026,  N1303,  N435,  N1657);
and AND2_448 (N3027,  N1663,  N1636);
and AND2_449 (N3028,  N1663,  N1642);
and AND2_450 (N3029,  N1663,  N1648);
and AND2_451 (N3030,  N1663,  N1654);
not NOT1_452 (N3031,  N1920);
not NOT1_453 (N3032,  N1923);
not NOT1_454 (N3033,  N1926);
not NOT1_455 (N3034,  N1929);
buf BUFF1_456 (N3035,  N1660);
buf BUFF1_457 (N3038,  N1660);
not NOT1_458 (N3041,  N1697);
not NOT1_459 (N3052,  N1709);
not NOT1_460 (N3063,  N1721);
not NOT1_461 (N3068,  N1727);
and AND2_462 (N3071,  N97,  N1721);
and AND2_463 (N3072,  N94,  N1721);
and AND2_464 (N3073,  N97,  N1721);
and AND2_465 (N3074,  N94,  N1721);
not NOT1_466 (N3075,  N1731);
not NOT1_467 (N3086,  N1743);
not NOT1_468 (N3097,  N1761);
not NOT1_469 (N3108,  N1769);
not NOT1_470 (N3119,  N1777);
not NOT1_471 (N3130,  N1785);
not NOT1_472 (N3141,  N1944);
not NOT1_473 (N3142,  N1947);
not NOT1_474 (N3143,  N1950);
not NOT1_475 (N3144,  N1953);
not NOT1_476 (N3145,  N1956);
not NOT1_477 (N3146,  N1959);
not NOT1_478 (N3147,  N1793);
not NOT1_479 (N3158,  N1800);
not NOT1_480 (N3169,  N1807);
not NOT1_481 (N3180,  N1814);
buf BUFF1_482 (N3191,  N1821);
not NOT1_483 (N3194,  N1932);
not NOT1_484 (N3195,  N1935);
not NOT1_485 (N3196,  N1938);
not NOT1_486 (N3197,  N1941);
not NOT1_487 (N3198,  N1962);
not NOT1_488 (N3199,  N1965);
buf BUFF1_489 (N3200,  N1469);
not NOT1_490 (N3203,  N1968);
buf BUFF1_491 (N3357,  N2704);
buf BUFF1_492 (N3358,  N2704);
buf BUFF1_493 (N3359,  N2704);
buf BUFF1_494 (N3360,  N2704);
and AND3_495 (N3401,  N457,  N1092,  N2824);
and AND3_496 (N3402,  N468,  N1092,  N2826);
and AND3_497 (N3403,  N422,  N1092,  N2828);
and AND3_498 (N3404,  N435,  N1092,  N2830);
and AND2_499 (N3405,  N1080,  N2823);
and AND2_500 (N3406,  N1080,  N2825);
and AND2_501 (N3407,  N1080,  N2827);
and AND2_502 (N3408,  N1080,  N2829);
and AND3_503 (N3409,  N389,  N1092,  N2840);
and AND3_504 (N3410,  N400,  N1092,  N2842);
and AND3_505 (N3411,  N411,  N1092,  N2844);
and AND3_506 (N3412,  N374,  N1092,  N2846);
and AND2_507 (N3413,  N1080,  N2839);
and AND2_508 (N3414,  N1080,  N2841);
and AND2_509 (N3415,  N1080,  N2843);
and AND2_510 (N3416,  N1080,  N2845);
and AND2_511 (N3444,  N1280,  N2902);
and AND3_512 (N3445,  N479,  N1280,  N2904);
and AND3_513 (N3446,  N490,  N1280,  N2906);
and AND2_514 (N3447,  N1685,  N2901);
and AND2_515 (N3448,  N1685,  N2903);
and AND2_516 (N3449,  N1685,  N2905);
and AND3_517 (N3450,  N503,  N1092,  N2914);
and AND3_518 (N3451,  N523,  N1092,  N2916);
and AND3_519 (N3452,  N534,  N1092,  N2918);
and AND2_520 (N3453,  N1080,  N2913);
and AND2_521 (N3454,  N1080,  N2915);
and AND2_522 (N3455,  N1080,  N2917);
and AND2_523 (N3456,  N2920,  N2350);
and AND3_524 (N3459,  N389,  N1280,  N2927);
and AND3_525 (N3460,  N400,  N1280,  N2929);
and AND3_526 (N3461,  N411,  N1280,  N2931);
and AND3_527 (N3462,  N374,  N1280,  N2933);
and AND2_528 (N3463,  N1685,  N2926);
and AND2_529 (N3464,  N1685,  N2928);
and AND2_530 (N3465,  N1685,  N2930);
and AND2_531 (N3466,  N1685,  N2932);
and AND3_532 (N3481,  N503,  N1292,  N2974);
not NOT1_533 (N3482,  N2980);
and AND3_534 (N3483,  N523,  N1292,  N2976);
and AND3_535 (N3484,  N534,  N1292,  N2978);
and AND2_536 (N3485,  N1271,  N2973);
and AND2_537 (N3486,  N1271,  N2975);
and AND2_538 (N3487,  N1271,  N2977);
and AND2_539 (N3488,  N1292,  N2988);
and AND3_540 (N3489,  N479,  N1292,  N2990);
and AND3_541 (N3490,  N490,  N1292,  N2992);
and AND2_542 (N3491,  N1271,  N2987);
and AND2_543 (N3492,  N1271,  N2989);
and AND2_544 (N3493,  N1271,  N2991);
and AND2_545 (N3502,  N1292,  N2999);
and AND2_546 (N3503,  N1292,  N3006);
and AND3_547 (N3504,  N457,  N1280,  N3016);
and AND3_548 (N3505,  N468,  N1280,  N3018);
and AND3_549 (N3506,  N422,  N1280,  N3020);
and AND3_550 (N3507,  N435,  N1280,  N3022);
and AND2_551 (N3508,  N1685,  N3015);
and AND2_552 (N3509,  N1685,  N3017);
and AND2_553 (N3510,  N1685,  N3019);
and AND2_554 (N3511,  N1685,  N3021);
nand NAND2_555 (N3512,  N1923,  N3031);
nand NAND2_556 (N3513,  N1920,  N3032);
nand NAND2_557 (N3514,  N1929,  N3033);
nand NAND2_558 (N3515,  N1926,  N3034);
nand NAND2_559 (N3558,  N1947,  N3141);
nand NAND2_560 (N3559,  N1944,  N3142);
nand NAND2_561 (N3560,  N1953,  N3143);
nand NAND2_562 (N3561,  N1950,  N3144);
nand NAND2_563 (N3562,  N1959,  N3145);
nand NAND2_564 (N3563,  N1956,  N3146);
buf BUFF1_565 (N3604,  N3191);
nand NAND2_566 (N3605,  N1935,  N3194);
nand NAND2_567 (N3606,  N1932,  N3195);
nand NAND2_568 (N3607,  N1941,  N3196);
nand NAND2_569 (N3608,  N1938,  N3197);
nand NAND2_570 (N3609,  N1965,  N3198);
nand NAND2_571 (N3610,  N1962,  N3199);
not NOT1_572 (N3613,  N3191);
and AND2_573 (N3614,  N2882,  N2891);
and AND2_574 (N3615,  N1482,  N2891);
and AND3_575 (N3616,  N200,  N2653,  N1173);
and AND3_576 (N3617,  N203,  N2653,  N1173);
and AND3_577 (N3618,  N197,  N2653,  N1173);
and AND3_578 (N3619,  N194,  N2653,  N1173);
and AND3_579 (N3620,  N191,  N2653,  N1173);
and AND3_580 (N3621,  N182,  N2681,  N1197);
and AND3_581 (N3622,  N188,  N2681,  N1197);
and AND3_582 (N3623,  N155,  N2681,  N1197);
and AND3_583 (N3624,  N149,  N2681,  N1197);
and AND2_584 (N3625,  N2882,  N2891);
and AND2_585 (N3626,  N1482,  N2891);
and AND3_586 (N3627,  N200,  N2728,  N1235);
and AND3_587 (N3628,  N203,  N2728,  N1235);
and AND3_588 (N3629,  N197,  N2728,  N1235);
and AND3_589 (N3630,  N194,  N2728,  N1235);
and AND3_590 (N3631,  N191,  N2728,  N1235);
and AND3_591 (N3632,  N182,  N2756,  N1259);
and AND3_592 (N3633,  N188,  N2756,  N1259);
and AND3_593 (N3634,  N155,  N2756,  N1259);
and AND3_594 (N3635,  N149,  N2756,  N1259);
and AND2_595 (N3636,  N2882,  N2891);
and AND2_596 (N3637,  N1482,  N2891);
and AND3_597 (N3638,  N109,  N3075,  N1743);
and AND2_598 (N3639,  N2882,  N2891);
and AND2_599 (N3640,  N1482,  N2891);
and AND3_600 (N3641,  N11,  N2779,  N1339);
and AND3_601 (N3642,  N109,  N3041,  N1709);
and AND3_602 (N3643,  N46,  N3041,  N1709);
and AND3_603 (N3644,  N100,  N3041,  N1709);
and AND3_604 (N3645,  N91,  N3041,  N1709);
and AND3_605 (N3646,  N43,  N3041,  N1709);
and AND3_606 (N3647,  N76,  N2779,  N1339);
and AND3_607 (N3648,  N73,  N2779,  N1339);
and AND3_608 (N3649,  N67,  N2779,  N1339);
and AND3_609 (N3650,  N14,  N2779,  N1339);
and AND3_610 (N3651,  N46,  N3075,  N1743);
and AND3_611 (N3652,  N100,  N3075,  N1743);
and AND3_612 (N3653,  N91,  N3075,  N1743);
and AND3_613 (N3654,  N43,  N3075,  N1743);
and AND3_614 (N3655,  N76,  N2801,  N1363);
and AND3_615 (N3656,  N73,  N2801,  N1363);
and AND3_616 (N3657,  N67,  N2801,  N1363);
and AND3_617 (N3658,  N14,  N2801,  N1363);
and AND3_618 (N3659,  N120,  N3119,  N1785);
and AND3_619 (N3660,  N11,  N2801,  N1363);
and AND3_620 (N3661,  N118,  N3097,  N1769);
and AND3_621 (N3662,  N176,  N2681,  N1197);
and AND3_622 (N3663,  N176,  N2756,  N1259);
or OR2_623 (N3664,  N2831,  N3401);
or OR2_624 (N3665,  N2832,  N3402);
or OR2_625 (N3666,  N2833,  N3403);
or OR2_626 (N3667,  N2834,  N3404);
or OR3_627 (N3668,  N2835,  N3405,  N457);
or OR3_628 (N3669,  N2836,  N3406,  N468);
or OR3_629 (N3670,  N2837,  N3407,  N422);
or OR3_630 (N3671,  N2838,  N3408,  N435);
or OR2_631 (N3672,  N2847,  N3409);
or OR2_632 (N3673,  N2848,  N3410);
or OR2_633 (N3674,  N2849,  N3411);
or OR2_634 (N3675,  N2850,  N3412);
or OR3_635 (N3676,  N2851,  N3413,  N389);
or OR3_636 (N3677,  N2852,  N3414,  N400);
or OR3_637 (N3678,  N2853,  N3415,  N411);
or OR3_638 (N3679,  N2854,  N3416,  N374);
and AND2_639 (N3680,  N289,  N2855);
and AND2_640 (N3681,  N281,  N2855);
and AND2_641 (N3682,  N273,  N2855);
and AND2_642 (N3683,  N265,  N2855);
and AND2_643 (N3684,  N257,  N2855);
and AND2_644 (N3685,  N234,  N2861);
and AND2_645 (N3686,  N226,  N2861);
and AND2_646 (N3687,  N218,  N2861);
and AND2_647 (N3688,  N210,  N2861);
and AND2_648 (N3689,  N206,  N2861);
not NOT1_649 (N3691,  N2891);
or OR2_650 (N3700,  N2907,  N3444);
or OR2_651 (N3701,  N2908,  N3445);
or OR2_652 (N3702,  N2909,  N3446);
or OR3_653 (N3703,  N2911,  N3448,  N479);
or OR3_654 (N3704,  N2912,  N3449,  N490);
or OR2_655 (N3705,  N2910,  N3447);
or OR2_656 (N3708,  N2919,  N3450);
or OR2_657 (N3709,  N2921,  N3451);
or OR2_658 (N3710,  N2922,  N3452);
or OR3_659 (N3711,  N2923,  N3453,  N503);
or OR3_660 (N3712,  N2924,  N3454,  N523);
or OR3_661 (N3713,  N2925,  N3455,  N534);
or OR2_662 (N3715,  N2934,  N3459);
or OR2_663 (N3716,  N2935,  N3460);
or OR2_664 (N3717,  N2936,  N3461);
or OR2_665 (N3718,  N2937,  N3462);
or OR3_666 (N3719,  N2938,  N3463,  N389);
or OR3_667 (N3720,  N2939,  N3464,  N400);
or OR3_668 (N3721,  N2940,  N3465,  N411);
or OR3_669 (N3722,  N2941,  N3466,  N374);
and AND2_670 (N3723,  N369,  N2942);
and AND2_671 (N3724,  N361,  N2942);
and AND2_672 (N3725,  N351,  N2942);
and AND2_673 (N3726,  N341,  N2942);
and AND2_674 (N3727,  N324,  N2948);
and AND2_675 (N3728,  N316,  N2948);
and AND2_676 (N3729,  N308,  N2948);
and AND2_677 (N3730,  N302,  N2948);
and AND2_678 (N3731,  N293,  N2948);
or OR2_679 (N3732,  N2942,  N2958);
and AND2_680 (N3738,  N83,  N2964);
and AND2_681 (N3739,  N87,  N2964);
and AND2_682 (N3740,  N34,  N2964);
and AND2_683 (N3741,  N34,  N2964);
or OR2_684 (N3742,  N2979,  N3481);
or OR2_685 (N3743,  N2981,  N3483);
or OR2_686 (N3744,  N2982,  N3484);
or OR3_687 (N3745,  N2983,  N3485,  N503);
or OR3_688 (N3746,  N2985,  N3486,  N523);
or OR3_689 (N3747,  N2986,  N3487,  N534);
or OR2_690 (N3748,  N2993,  N3488);
or OR2_691 (N3749,  N2994,  N3489);
or OR2_692 (N3750,  N2995,  N3490);
or OR3_693 (N3751,  N2997,  N3492,  N479);
or OR3_694 (N3752,  N2998,  N3493,  N490);
not NOT1_695 (N3753,  N3000);
not NOT1_696 (N3754,  N3003);
not NOT1_697 (N3755,  N3007);
not NOT1_698 (N3756,  N3010);
or OR2_699 (N3757,  N3013,  N3502);
and AND3_700 (N3758,  N1315,  N446,  N3003);
or OR2_701 (N3759,  N3014,  N3503);
and AND3_702 (N3760,  N1315,  N446,  N3010);
and AND2_703 (N3761,  N1675,  N3000);
and AND2_704 (N3762,  N1675,  N3007);
or OR2_705 (N3763,  N3023,  N3504);
or OR2_706 (N3764,  N3024,  N3505);
or OR2_707 (N3765,  N3025,  N3506);
or OR2_708 (N3766,  N3026,  N3507);
or OR3_709 (N3767,  N3027,  N3508,  N457);
or OR3_710 (N3768,  N3028,  N3509,  N468);
or OR3_711 (N3769,  N3029,  N3510,  N422);
or OR3_712 (N3770,  N3030,  N3511,  N435);
nand NAND2_713 (N3771,  N3512,  N3513);
nand NAND2_714 (N3775,  N3514,  N3515);
not NOT1_715 (N3779,  N3035);
not NOT1_716 (N3780,  N3038);
and AND3_717 (N3781,  N117,  N3097,  N1769);
and AND3_718 (N3782,  N126,  N3097,  N1769);
and AND3_719 (N3783,  N127,  N3097,  N1769);
and AND3_720 (N3784,  N128,  N3097,  N1769);
and AND3_721 (N3785,  N131,  N3119,  N1785);
and AND3_722 (N3786,  N129,  N3119,  N1785);
and AND3_723 (N3787,  N119,  N3119,  N1785);
and AND3_724 (N3788,  N130,  N3119,  N1785);
nand NAND2_725 (N3789,  N3558,  N3559);
nand NAND2_726 (N3793,  N3560,  N3561);
nand NAND2_727 (N3797,  N3562,  N3563);
and AND3_728 (N3800,  N122,  N3147,  N1800);
and AND3_729 (N3801,  N113,  N3147,  N1800);
and AND3_730 (N3802,  N53,  N3147,  N1800);
and AND3_731 (N3803,  N114,  N3147,  N1800);
and AND3_732 (N3804,  N115,  N3147,  N1800);
and AND3_733 (N3805,  N52,  N3169,  N1814);
and AND3_734 (N3806,  N112,  N3169,  N1814);
and AND3_735 (N3807,  N116,  N3169,  N1814);
and AND3_736 (N3808,  N121,  N3169,  N1814);
and AND3_737 (N3809,  N123,  N3169,  N1814);
nand NAND2_738 (N3810,  N3607,  N3608);
nand NAND2_739 (N3813,  N3605,  N3606);
and AND2_740 (N3816,  N3482,  N2984);
or OR2_741 (N3819,  N2996,  N3491);
not NOT1_742 (N3822,  N3200);
nand NAND2_743 (N3823,  N3200,  N3203);
nand NAND2_744 (N3824,  N3609,  N3610);
not NOT1_745 (N3827,  N3456);
or OR2_746 (N3828,  N3739,  N2970);
or OR2_747 (N3829,  N3740,  N2971);
or OR2_748 (N3830,  N3741,  N2972);
or OR2_749 (N3831,  N3738,  N2969);
not NOT1_750 (N3834,  N3664);
not NOT1_751 (N3835,  N3665);
not NOT1_752 (N3836,  N3666);
not NOT1_753 (N3837,  N3667);
not NOT1_754 (N3838,  N3672);
not NOT1_755 (N3839,  N3673);
not NOT1_756 (N3840,  N3674);
not NOT1_757 (N3841,  N3675);
or OR2_758 (N3842,  N3681,  N2868);
or OR2_759 (N3849,  N3682,  N2869);
or OR2_760 (N3855,  N3683,  N2870);
or OR2_761 (N3861,  N3684,  N2871);
or OR2_762 (N3867,  N3685,  N2872);
or OR2_763 (N3873,  N3686,  N2873);
or OR2_764 (N3881,  N3687,  N2874);
or OR2_765 (N3887,  N3688,  N2875);
or OR2_766 (N3893,  N3689,  N2876);
not NOT1_767 (N3908,  N3701);
not NOT1_768 (N3909,  N3702);
not NOT1_769 (N3911,  N3700);
not NOT1_770 (N3914,  N3708);
not NOT1_771 (N3915,  N3709);
not NOT1_772 (N3916,  N3710);
not NOT1_773 (N3917,  N3715);
not NOT1_774 (N3918,  N3716);
not NOT1_775 (N3919,  N3717);
not NOT1_776 (N3920,  N3718);
or OR2_777 (N3921,  N3724,  N2955);
or OR2_778 (N3927,  N3725,  N2956);
or OR2_779 (N3933,  N3726,  N2957);
or OR2_780 (N3942,  N3727,  N2959);
or OR2_781 (N3948,  N3728,  N2960);
or OR2_782 (N3956,  N3729,  N2961);
or OR2_783 (N3962,  N3730,  N2962);
or OR2_784 (N3968,  N3731,  N2963);
not NOT1_785 (N3975,  N3742);
not NOT1_786 (N3976,  N3743);
not NOT1_787 (N3977,  N3744);
not NOT1_788 (N3978,  N3749);
not NOT1_789 (N3979,  N3750);
and AND3_790 (N3980,  N446,  N1292,  N3754);
and AND3_791 (N3981,  N446,  N1292,  N3756);
and AND2_792 (N3982,  N1271,  N3753);
and AND2_793 (N3983,  N1271,  N3755);
not NOT1_794 (N3984,  N3757);
not NOT1_795 (N3987,  N3759);
not NOT1_796 (N3988,  N3763);
not NOT1_797 (N3989,  N3764);
not NOT1_798 (N3990,  N3765);
not NOT1_799 (N3991,  N3766);
and AND3_800 (N3998,  N3456,  N3119,  N3130);
or OR2_801 (N4008,  N3723,  N2954);
or OR2_802 (N4011,  N3680,  N2867);
not NOT1_803 (N4021,  N3748);
nand NAND2_804 (N4024,  N1968,  N3822);
not NOT1_805 (N4027,  N3705);
and AND2_806 (N4031,  N3828,  N1583);
and AND3_807 (N4032,  N24,  N2882,  N3691);
and AND3_808 (N4033,  N25,  N1482,  N3691);
and AND3_809 (N4034,  N26,  N2882,  N3691);
and AND3_810 (N4035,  N81,  N1482,  N3691);
and AND2_811 (N4036,  N3829,  N1583);
and AND3_812 (N4037,  N79,  N2882,  N3691);
and AND3_813 (N4038,  N23,  N1482,  N3691);
and AND3_814 (N4039,  N82,  N2882,  N3691);
and AND3_815 (N4040,  N80,  N1482,  N3691);
and AND2_816 (N4041,  N3830,  N1583);
and AND2_817 (N4042,  N3831,  N1583);
and AND2_818 (N4067,  N3732,  N514);
and AND2_819 (N4080,  N514,  N3732);
and AND2_820 (N4088,  N3834,  N3668);
and AND2_821 (N4091,  N3835,  N3669);
and AND2_822 (N4094,  N3836,  N3670);
and AND2_823 (N4097,  N3837,  N3671);
and AND2_824 (N4100,  N3838,  N3676);
and AND2_825 (N4103,  N3839,  N3677);
and AND2_826 (N4106,  N3840,  N3678);
and AND2_827 (N4109,  N3841,  N3679);
and AND2_828 (N4144,  N3908,  N3703);
and AND2_829 (N4147,  N3909,  N3704);
buf BUFF1_830 (N4150,  N3705);
and AND2_831 (N4153,  N3914,  N3711);
and AND2_832 (N4156,  N3915,  N3712);
and AND2_833 (N4159,  N3916,  N3713);
or OR2_834 (N4183,  N3758,  N3980);
or OR2_835 (N4184,  N3760,  N3981);
or OR3_836 (N4185,  N3761,  N3982,  N446);
or OR3_837 (N4186,  N3762,  N3983,  N446);
not NOT1_838 (N4188,  N3771);
not NOT1_839 (N4191,  N3775);
and AND3_840 (N4196,  N3775,  N3771,  N3035);
and AND3_841 (N4197,  N3987,  N3119,  N3130);
and AND2_842 (N4198,  N3920,  N3722);
not NOT1_843 (N4199,  N3816);
not NOT1_844 (N4200,  N3789);
not NOT1_845 (N4203,  N3793);
buf BUFF1_846 (N4206,  N3797);
buf BUFF1_847 (N4209,  N3797);
buf BUFF1_848 (N4212,  N3732);
buf BUFF1_849 (N4215,  N3732);
buf BUFF1_850 (N4219,  N3732);
not NOT1_851 (N4223,  N3810);
not NOT1_852 (N4224,  N3813);
and AND2_853 (N4225,  N3918,  N3720);
and AND2_854 (N4228,  N3919,  N3721);
and AND2_855 (N4231,  N3991,  N3770);
and AND2_856 (N4234,  N3917,  N3719);
and AND2_857 (N4237,  N3989,  N3768);
and AND2_858 (N4240,  N3990,  N3769);
and AND2_859 (N4243,  N3988,  N3767);
and AND2_860 (N4246,  N3976,  N3746);
and AND2_861 (N4249,  N3977,  N3747);
and AND2_862 (N4252,  N3975,  N3745);
and AND2_863 (N4255,  N3978,  N3751);
and AND2_864 (N4258,  N3979,  N3752);
not NOT1_865 (N4263,  N3819);
nand NAND2_866 (N4264,  N4024,  N3823);
not NOT1_867 (N4267,  N3824);
and AND2_868 (N4268,  N446,  N3893);
not NOT1_869 (N4269,  N3911);
not NOT1_870 (N4270,  N3984);
and AND2_871 (N4271,  N3893,  N446);
not NOT1_872 (N4272,  N4031);
or OR4_873 (N4273,  N4032,  N4033,  N3614,  N3615);
or OR4_874 (N4274,  N4034,  N4035,  N3625,  N3626);
not NOT1_875 (N4275,  N4036);
or OR4_876 (N4276,  N4037,  N4038,  N3636,  N3637);
or OR4_877 (N4277,  N4039,  N4040,  N3639,  N3640);
not NOT1_878 (N4278,  N4041);
not NOT1_879 (N4279,  N4042);
and AND2_880 (N4280,  N3887,  N457);
and AND2_881 (N4284,  N3881,  N468);
and AND2_882 (N4290,  N422,  N3873);
and AND2_883 (N4297,  N3867,  N435);
and AND2_884 (N4298,  N3861,  N389);
and AND2_885 (N4301,  N3855,  N400);
and AND2_886 (N4305,  N3849,  N411);
and AND2_887 (N4310,  N3842,  N374);
and AND2_888 (N4316,  N457,  N3887);
and AND2_889 (N4320,  N468,  N3881);
and AND2_890 (N4325,  N422,  N3873);
and AND2_891 (N4331,  N435,  N3867);
and AND2_892 (N4332,  N389,  N3861);
and AND2_893 (N4336,  N400,  N3855);
and AND2_894 (N4342,  N411,  N3849);
and AND2_895 (N4349,  N374,  N3842);
not NOT1_896 (N4357,  N3968);
not NOT1_897 (N4364,  N3962);
buf BUFF1_898 (N4375,  N3962);
and AND2_899 (N4379,  N3956,  N479);
and AND2_900 (N4385,  N490,  N3948);
and AND2_901 (N4392,  N3942,  N503);
and AND2_902 (N4396,  N3933,  N523);
and AND2_903 (N4400,  N3927,  N534);
not NOT1_904 (N4405,  N3921);
buf BUFF1_905 (N4412,  N3921);
not NOT1_906 (N4418,  N3968);
not NOT1_907 (N4425,  N3962);
buf BUFF1_908 (N4436,  N3962);
and AND2_909 (N4440,  N479,  N3956);
and AND2_910 (N4445,  N490,  N3948);
and AND2_911 (N4451,  N503,  N3942);
and AND2_912 (N4456,  N523,  N3933);
and AND2_913 (N4462,  N534,  N3927);
buf BUFF1_914 (N4469,  N3921);
not NOT1_915 (N4477,  N3921);
buf BUFF1_916 (N4512,  N3968);
not NOT1_917 (N4515,  N4183);
not NOT1_918 (N4516,  N4184);
not NOT1_919 (N4521,  N4008);
not NOT1_920 (N4523,  N4011);
not NOT1_921 (N4524,  N4198);
not NOT1_922 (N4532,  N3984);
and AND3_923 (N4547,  N3911,  N3169,  N3180);
buf BUFF1_924 (N4548,  N3893);
buf BUFF1_925 (N4551,  N3887);
buf BUFF1_926 (N4554,  N3881);
buf BUFF1_927 (N4557,  N3873);
buf BUFF1_928 (N4560,  N3867);
buf BUFF1_929 (N4563,  N3861);
buf BUFF1_930 (N4566,  N3855);
buf BUFF1_931 (N4569,  N3849);
buf BUFF1_932 (N4572,  N3842);
nor NOR2_933 (N4575,  N422,  N3873);
buf BUFF1_934 (N4578,  N3893);
buf BUFF1_935 (N4581,  N3887);
buf BUFF1_936 (N4584,  N3881);
buf BUFF1_937 (N4587,  N3867);
buf BUFF1_938 (N4590,  N3861);
buf BUFF1_939 (N4593,  N3855);
buf BUFF1_940 (N4596,  N3849);
buf BUFF1_941 (N4599,  N3873);
buf BUFF1_942 (N4602,  N3842);
nor NOR2_943 (N4605,  N422,  N3873);
nor NOR2_944 (N4608,  N374,  N3842);
buf BUFF1_945 (N4611,  N3956);
buf BUFF1_946 (N4614,  N3948);
buf BUFF1_947 (N4617,  N3942);
buf BUFF1_948 (N4621,  N3933);
buf BUFF1_949 (N4624,  N3927);
nor NOR2_950 (N4627,  N490,  N3948);
buf BUFF1_951 (N4630,  N3956);
buf BUFF1_952 (N4633,  N3942);
buf BUFF1_953 (N4637,  N3933);
buf BUFF1_954 (N4640,  N3927);
buf BUFF1_955 (N4643,  N3948);
nor NOR2_956 (N4646,  N490,  N3948);
buf BUFF1_957 (N4649,  N3927);
buf BUFF1_958 (N4652,  N3933);
buf BUFF1_959 (N4655,  N3921);
buf BUFF1_960 (N4658,  N3942);
buf BUFF1_961 (N4662,  N3956);
buf BUFF1_962 (N4665,  N3948);
buf BUFF1_963 (N4668,  N3968);
buf BUFF1_964 (N4671,  N3962);
buf BUFF1_965 (N4674,  N3873);
buf BUFF1_966 (N4677,  N3867);
buf BUFF1_967 (N4680,  N3887);
buf BUFF1_968 (N4683,  N3881);
buf BUFF1_969 (N4686,  N3893);
buf BUFF1_970 (N4689,  N3849);
buf BUFF1_971 (N4692,  N3842);
buf BUFF1_972 (N4695,  N3861);
buf BUFF1_973 (N4698,  N3855);
nand NAND2_974 (N4701,  N3813,  N4223);
nand NAND2_975 (N4702,  N3810,  N4224);
not NOT1_976 (N4720,  N4021);
nand NAND2_977 (N4721,  N4021,  N4263);
not NOT1_978 (N4724,  N4147);
not NOT1_979 (N4725,  N4144);
not NOT1_980 (N4726,  N4159);
not NOT1_981 (N4727,  N4156);
not NOT1_982 (N4728,  N4153);
not NOT1_983 (N4729,  N4097);
not NOT1_984 (N4730,  N4094);
not NOT1_985 (N4731,  N4091);
not NOT1_986 (N4732,  N4088);
not NOT1_987 (N4733,  N4109);
not NOT1_988 (N4734,  N4106);
not NOT1_989 (N4735,  N4103);
not NOT1_990 (N4736,  N4100);
and AND2_991 (N4737,  N4273,  N2877);
and AND2_992 (N4738,  N4274,  N2877);
and AND2_993 (N4739,  N4276,  N2877);
and AND2_994 (N4740,  N4277,  N2877);
and AND3_995 (N4741,  N4150,  N1758,  N1755);
not NOT1_996 (N4855,  N4212);
nand NAND2_997 (N4856,  N4212,  N2712);
nand NAND2_998 (N4908,  N4215,  N2718);
not NOT1_999 (N4909,  N4215);
and AND2_1000 (N4939,  N4515,  N4185);
and AND2_1001 (N4942,  N4516,  N4186);
not NOT1_1002 (N4947,  N4219);
and AND3_1003 (N4953,  N4188,  N3775,  N3779);
and AND3_1004 (N4954,  N3771,  N4191,  N3780);
and AND3_1005 (N4955,  N4191,  N4188,  N3038);
and AND3_1006 (N4956,  N4109,  N3097,  N3108);
and AND3_1007 (N4957,  N4106,  N3097,  N3108);
and AND3_1008 (N4958,  N4103,  N3097,  N3108);
and AND3_1009 (N4959,  N4100,  N3097,  N3108);
and AND3_1010 (N4960,  N4159,  N3119,  N3130);
and AND3_1011 (N4961,  N4156,  N3119,  N3130);
not NOT1_1012 (N4965,  N4225);
not NOT1_1013 (N4966,  N4228);
not NOT1_1014 (N4967,  N4231);
not NOT1_1015 (N4968,  N4234);
not NOT1_1016 (N4972,  N4246);
not NOT1_1017 (N4973,  N4249);
not NOT1_1018 (N4974,  N4252);
nand NAND2_1019 (N4975,  N4252,  N4199);
not NOT1_1020 (N4976,  N4206);
not NOT1_1021 (N4977,  N4209);
and AND3_1022 (N4978,  N3793,  N3789,  N4206);
and AND3_1023 (N4979,  N4203,  N4200,  N4209);
and AND3_1024 (N4980,  N4097,  N3147,  N3158);
and AND3_1025 (N4981,  N4094,  N3147,  N3158);
and AND3_1026 (N4982,  N4091,  N3147,  N3158);
and AND3_1027 (N4983,  N4088,  N3147,  N3158);
and AND3_1028 (N4984,  N4153,  N3169,  N3180);
and AND3_1029 (N4985,  N4147,  N3169,  N3180);
and AND3_1030 (N4986,  N4144,  N3169,  N3180);
and AND3_1031 (N4987,  N4150,  N3169,  N3180);
nand NAND2_1032 (N5049,  N4701,  N4702);
not NOT1_1033 (N5052,  N4237);
not NOT1_1034 (N5053,  N4240);
not NOT1_1035 (N5054,  N4243);
not NOT1_1036 (N5055,  N4255);
not NOT1_1037 (N5056,  N4258);
nand NAND2_1038 (N5057,  N3819,  N4720);
not NOT1_1039 (N5058,  N4264);
nand NAND2_1040 (N5059,  N4264,  N4267);
and AND4_1041 (N5060,  N4724,  N4725,  N4269,  N4027);
and AND4_1042 (N5061,  N4726,  N4727,  N3827,  N4728);
and AND4_1043 (N5062,  N4729,  N4730,  N4731,  N4732);
and AND4_1044 (N5063,  N4733,  N4734,  N4735,  N4736);
and AND2_1045 (N5065,  N4357,  N4375);
and AND3_1046 (N5066,  N4364,  N4357,  N4379);
and AND2_1047 (N5067,  N4418,  N4436);
and AND3_1048 (N5068,  N4425,  N4418,  N4440);
not NOT1_1049 (N5069,  N4548);
nand NAND2_1050 (N5070,  N4548,  N2628);
not NOT1_1051 (N5071,  N4551);
nand NAND2_1052 (N5072,  N4551,  N2629);
not NOT1_1053 (N5073,  N4554);
nand NAND2_1054 (N5074,  N4554,  N2630);
not NOT1_1055 (N5075,  N4557);
nand NAND2_1056 (N5076,  N4557,  N2631);
not NOT1_1057 (N5077,  N4560);
nand NAND2_1058 (N5078,  N4560,  N2632);
not NOT1_1059 (N5079,  N4563);
nand NAND2_1060 (N5080,  N4563,  N2633);
not NOT1_1061 (N5081,  N4566);
nand NAND2_1062 (N5082,  N4566,  N2634);
not NOT1_1063 (N5083,  N4569);
nand NAND2_1064 (N5084,  N4569,  N2635);
not NOT1_1065 (N5085,  N4572);
nand NAND2_1066 (N5086,  N4572,  N2636);
not NOT1_1067 (N5087,  N4575);
nand NAND2_1068 (N5088,  N4578,  N2638);
not NOT1_1069 (N5089,  N4578);
nand NAND2_1070 (N5090,  N4581,  N2639);
not NOT1_1071 (N5091,  N4581);
nand NAND2_1072 (N5092,  N4584,  N2640);
not NOT1_1073 (N5093,  N4584);
nand NAND2_1074 (N5094,  N4587,  N2641);
not NOT1_1075 (N5095,  N4587);
nand NAND2_1076 (N5096,  N4590,  N2642);
not NOT1_1077 (N5097,  N4590);
nand NAND2_1078 (N5098,  N4593,  N2643);
not NOT1_1079 (N5099,  N4593);
nand NAND2_1080 (N5100,  N4596,  N2644);
not NOT1_1081 (N5101,  N4596);
nand NAND2_1082 (N5102,  N4599,  N2645);
not NOT1_1083 (N5103,  N4599);
nand NAND2_1084 (N5104,  N4602,  N2646);
not NOT1_1085 (N5105,  N4602);
not NOT1_1086 (N5106,  N4611);
nand NAND2_1087 (N5107,  N4611,  N2709);
not NOT1_1088 (N5108,  N4614);
nand NAND2_1089 (N5109,  N4614,  N2710);
not NOT1_1090 (N5110,  N4617);
nand NAND2_1091 (N5111,  N4617,  N2711);
nand NAND2_1092 (N5112,  N1890,  N4855);
not NOT1_1093 (N5113,  N4621);
nand NAND2_1094 (N5114,  N4621,  N2713);
not NOT1_1095 (N5115,  N4624);
nand NAND2_1096 (N5116,  N4624,  N2714);
and AND2_1097 (N5117,  N4364,  N4379);
and AND2_1098 (N5118,  N4364,  N4379);
and AND2_1099 (N5119,  N54,  N4405);
not NOT1_1100 (N5120,  N4627);
nand NAND2_1101 (N5121,  N4630,  N2716);
not NOT1_1102 (N5122,  N4630);
nand NAND2_1103 (N5123,  N4633,  N2717);
not NOT1_1104 (N5124,  N4633);
nand NAND2_1105 (N5125,  N1908,  N4909);
nand NAND2_1106 (N5126,  N4637,  N2719);
not NOT1_1107 (N5127,  N4637);
nand NAND2_1108 (N5128,  N4640,  N2720);
not NOT1_1109 (N5129,  N4640);
nand NAND2_1110 (N5130,  N4643,  N2721);
not NOT1_1111 (N5131,  N4643);
and AND2_1112 (N5132,  N4425,  N4440);
and AND2_1113 (N5133,  N4425,  N4440);
not NOT1_1114 (N5135,  N4649);
not NOT1_1115 (N5136,  N4652);
nand NAND2_1116 (N5137,  N4655,  N4521);
not NOT1_1117 (N5138,  N4655);
not NOT1_1118 (N5139,  N4658);
nand NAND2_1119 (N5140,  N4658,  N4947);
not NOT1_1120 (N5141,  N4674);
not NOT1_1121 (N5142,  N4677);
not NOT1_1122 (N5143,  N4680);
not NOT1_1123 (N5144,  N4683);
nand NAND2_1124 (N5145,  N4686,  N4523);
not NOT1_1125 (N5146,  N4686);
nor NOR2_1126 (N5147,  N4953,  N4196);
nor NOR2_1127 (N5148,  N4954,  N4955);
not NOT1_1128 (N5150,  N4524);
nand NAND2_1129 (N5153,  N4228,  N4965);
nand NAND2_1130 (N5154,  N4225,  N4966);
nand NAND2_1131 (N5155,  N4234,  N4967);
nand NAND2_1132 (N5156,  N4231,  N4968);
not NOT1_1133 (N5157,  N4532);
nand NAND2_1134 (N5160,  N4249,  N4972);
nand NAND2_1135 (N5161,  N4246,  N4973);
nand NAND2_1136 (N5162,  N3816,  N4974);
and AND3_1137 (N5163,  N4200,  N3793,  N4976);
and AND3_1138 (N5164,  N3789,  N4203,  N4977);
and AND3_1139 (N5165,  N4942,  N3147,  N3158);
not NOT1_1140 (N5166,  N4512);
buf BUFF1_1141 (N5169,  N4290);
not NOT1_1142 (N5172,  N4605);
buf BUFF1_1143 (N5173,  N4325);
not NOT1_1144 (N5176,  N4608);
buf BUFF1_1145 (N5177,  N4349);
buf BUFF1_1146 (N5180,  N4405);
buf BUFF1_1147 (N5183,  N4357);
buf BUFF1_1148 (N5186,  N4357);
buf BUFF1_1149 (N5189,  N4364);
buf BUFF1_1150 (N5192,  N4364);
buf BUFF1_1151 (N5195,  N4385);
not NOT1_1152 (N5198,  N4646);
buf BUFF1_1153 (N5199,  N4418);
buf BUFF1_1154 (N5202,  N4425);
buf BUFF1_1155 (N5205,  N4445);
buf BUFF1_1156 (N5208,  N4418);
buf BUFF1_1157 (N5211,  N4425);
buf BUFF1_1158 (N5214,  N4477);
buf BUFF1_1159 (N5217,  N4469);
buf BUFF1_1160 (N5220,  N4477);
not NOT1_1161 (N5223,  N4662);
not NOT1_1162 (N5224,  N4665);
not NOT1_1163 (N5225,  N4668);
not NOT1_1164 (N5226,  N4671);
not NOT1_1165 (N5227,  N4689);
not NOT1_1166 (N5228,  N4692);
not NOT1_1167 (N5229,  N4695);
not NOT1_1168 (N5230,  N4698);
nand NAND2_1169 (N5232,  N4240,  N5052);
nand NAND2_1170 (N5233,  N4237,  N5053);
nand NAND2_1171 (N5234,  N4258,  N5055);
nand NAND2_1172 (N5235,  N4255,  N5056);
nand NAND2_1173 (N5236,  N4721,  N5057);
nand NAND2_1174 (N5239,  N3824,  N5058);
and AND3_1175 (N5240,  N5060,  N5061,  N4270);
not NOT1_1176 (N5241,  N4939);
nand NAND2_1177 (N5242,  N1824,  N5069);
nand NAND2_1178 (N5243,  N1827,  N5071);
nand NAND2_1179 (N5244,  N1830,  N5073);
nand NAND2_1180 (N5245,  N1833,  N5075);
nand NAND2_1181 (N5246,  N1836,  N5077);
nand NAND2_1182 (N5247,  N1839,  N5079);
nand NAND2_1183 (N5248,  N1842,  N5081);
nand NAND2_1184 (N5249,  N1845,  N5083);
nand NAND2_1185 (N5250,  N1848,  N5085);
nand NAND2_1186 (N5252,  N1854,  N5089);
nand NAND2_1187 (N5253,  N1857,  N5091);
nand NAND2_1188 (N5254,  N1860,  N5093);
nand NAND2_1189 (N5255,  N1863,  N5095);
nand NAND2_1190 (N5256,  N1866,  N5097);
nand NAND2_1191 (N5257,  N1869,  N5099);
nand NAND2_1192 (N5258,  N1872,  N5101);
nand NAND2_1193 (N5259,  N1875,  N5103);
nand NAND2_1194 (N5260,  N1878,  N5105);
nand NAND2_1195 (N5261,  N1881,  N5106);
nand NAND2_1196 (N5262,  N1884,  N5108);
nand NAND2_1197 (N5263,  N1887,  N5110);
nand NAND2_1198 (N5264,  N5112,  N4856);
nand NAND2_1199 (N5274,  N1893,  N5113);
nand NAND2_1200 (N5275,  N1896,  N5115);
nand NAND2_1201 (N5282,  N1902,  N5122);
nand NAND2_1202 (N5283,  N1905,  N5124);
nand NAND2_1203 (N5284,  N4908,  N5125);
nand NAND2_1204 (N5298,  N1911,  N5127);
nand NAND2_1205 (N5299,  N1914,  N5129);
nand NAND2_1206 (N5300,  N1917,  N5131);
nand NAND2_1207 (N5303,  N4652,  N5135);
nand NAND2_1208 (N5304,  N4649,  N5136);
nand NAND2_1209 (N5305,  N4008,  N5138);
nand NAND2_1210 (N5306,  N4219,  N5139);
nand NAND2_1211 (N5307,  N4677,  N5141);
nand NAND2_1212 (N5308,  N4674,  N5142);
nand NAND2_1213 (N5309,  N4683,  N5143);
nand NAND2_1214 (N5310,  N4680,  N5144);
nand NAND2_1215 (N5311,  N4011,  N5146);
not NOT1_1216 (N5312,  N5049);
nand NAND2_1217 (N5315,  N5153,  N5154);
nand NAND2_1218 (N5319,  N5155,  N5156);
nand NAND2_1219 (N5324,  N5160,  N5161);
nand NAND2_1220 (N5328,  N5162,  N4975);
nor NOR2_1221 (N5331,  N5163,  N4978);
nor NOR2_1222 (N5332,  N5164,  N4979);
or OR2_1223 (N5346,  N4412,  N5119);
nand NAND2_1224 (N5363,  N4665,  N5223);
nand NAND2_1225 (N5364,  N4662,  N5224);
nand NAND2_1226 (N5365,  N4671,  N5225);
nand NAND2_1227 (N5366,  N4668,  N5226);
nand NAND2_1228 (N5367,  N4692,  N5227);
nand NAND2_1229 (N5368,  N4689,  N5228);
nand NAND2_1230 (N5369,  N4698,  N5229);
nand NAND2_1231 (N5370,  N4695,  N5230);
nand NAND2_1232 (N5371,  N5148,  N5147);
buf BUFF1_1233 (N5374,  N4939);
nand NAND2_1234 (N5377,  N5232,  N5233);
nand NAND2_1235 (N5382,  N5234,  N5235);
nand NAND2_1236 (N5385,  N5239,  N5059);
and AND3_1237 (N5388,  N5062,  N5063,  N5241);
nand NAND2_1238 (N5389,  N5242,  N5070);
nand NAND2_1239 (N5396,  N5243,  N5072);
nand NAND2_1240 (N5407,  N5244,  N5074);
nand NAND2_1241 (N5418,  N5245,  N5076);
nand NAND2_1242 (N5424,  N5246,  N5078);
nand NAND2_1243 (N5431,  N5247,  N5080);
nand NAND2_1244 (N5441,  N5248,  N5082);
nand NAND2_1245 (N5452,  N5249,  N5084);
nand NAND2_1246 (N5462,  N5250,  N5086);
not NOT1_1247 (N5469,  N5169);
nand NAND2_1248 (N5470,  N5088,  N5252);
nand NAND2_1249 (N5477,  N5090,  N5253);
nand NAND2_1250 (N5488,  N5092,  N5254);
nand NAND2_1251 (N5498,  N5094,  N5255);
nand NAND2_1252 (N5506,  N5096,  N5256);
nand NAND2_1253 (N5520,  N5098,  N5257);
nand NAND2_1254 (N5536,  N5100,  N5258);
nand NAND2_1255 (N5549,  N5102,  N5259);
nand NAND2_1256 (N5555,  N5104,  N5260);
nand NAND2_1257 (N5562,  N5261,  N5107);
nand NAND2_1258 (N5573,  N5262,  N5109);
nand NAND2_1259 (N5579,  N5263,  N5111);
nand NAND2_1260 (N5595,  N5274,  N5114);
nand NAND2_1261 (N5606,  N5275,  N5116);
nand NAND2_1262 (N5616,  N5180,  N2715);
not NOT1_1263 (N5617,  N5180);
not NOT1_1264 (N5618,  N5183);
not NOT1_1265 (N5619,  N5186);
not NOT1_1266 (N5620,  N5189);
not NOT1_1267 (N5621,  N5192);
not NOT1_1268 (N5622,  N5195);
nand NAND2_1269 (N5624,  N5121,  N5282);
nand NAND2_1270 (N5634,  N5123,  N5283);
nand NAND2_1271 (N5655,  N5126,  N5298);
nand NAND2_1272 (N5671,  N5128,  N5299);
nand NAND2_1273 (N5684,  N5130,  N5300);
not NOT1_1274 (N5690,  N5202);
not NOT1_1275 (N5691,  N5211);
nand NAND2_1276 (N5692,  N5303,  N5304);
nand NAND2_1277 (N5696,  N5137,  N5305);
nand NAND2_1278 (N5700,  N5306,  N5140);
nand NAND2_1279 (N5703,  N5307,  N5308);
nand NAND2_1280 (N5707,  N5309,  N5310);
nand NAND2_1281 (N5711,  N5145,  N5311);
and AND2_1282 (N5726,  N5166,  N4512);
not NOT1_1283 (N5727,  N5173);
not NOT1_1284 (N5728,  N5177);
not NOT1_1285 (N5730,  N5199);
not NOT1_1286 (N5731,  N5205);
not NOT1_1287 (N5732,  N5208);
not NOT1_1288 (N5733,  N5214);
not NOT1_1289 (N5734,  N5217);
not NOT1_1290 (N5735,  N5220);
nand NAND2_1291 (N5736,  N5365,  N5366);
nand NAND2_1292 (N5739,  N5363,  N5364);
nand NAND2_1293 (N5742,  N5369,  N5370);
nand NAND2_1294 (N5745,  N5367,  N5368);
not NOT1_1295 (N5755,  N5236);
nand NAND2_1296 (N5756,  N5332,  N5331);
and AND2_1297 (N5954,  N5264,  N4396);
nand NAND2_1298 (N5955,  N1899,  N5617);
not NOT1_1299 (N5956,  N5346);
and AND2_1300 (N6005,  N5284,  N4456);
and AND2_1301 (N6006,  N5284,  N4456);
not NOT1_1302 (N6023,  N5371);
nand NAND2_1303 (N6024,  N5371,  N5312);
not NOT1_1304 (N6025,  N5315);
not NOT1_1305 (N6028,  N5324);
buf BUFF1_1306 (N6031,  N5319);
buf BUFF1_1307 (N6034,  N5319);
buf BUFF1_1308 (N6037,  N5328);
buf BUFF1_1309 (N6040,  N5328);
not NOT1_1310 (N6044,  N5385);
or OR2_1311 (N6045,  N5166,  N5726);
buf BUFF1_1312 (N6048,  N5264);
buf BUFF1_1313 (N6051,  N5284);
buf BUFF1_1314 (N6054,  N5284);
not NOT1_1315 (N6065,  N5374);
nand NAND2_1316 (N6066,  N5374,  N5054);
not NOT1_1317 (N6067,  N5377);
not NOT1_1318 (N6068,  N5382);
nand NAND2_1319 (N6069,  N5382,  N5755);
and AND2_1320 (N6071,  N5470,  N4316);
and AND3_1321 (N6072,  N5477,  N5470,  N4320);
and AND4_1322 (N6073,  N5488,  N5470,  N4325,  N5477);
and AND4_1323 (N6074,  N5562,  N4357,  N4385,  N4364);
and AND2_1324 (N6075,  N5389,  N4280);
and AND3_1325 (N6076,  N5396,  N5389,  N4284);
and AND4_1326 (N6077,  N5407,  N5389,  N4290,  N5396);
and AND4_1327 (N6078,  N5624,  N4418,  N4445,  N4425);
not NOT1_1328 (N6079,  N5418);
and AND4_1329 (N6080,  N5396,  N5418,  N5407,  N5389);
and AND2_1330 (N6083,  N5396,  N4284);
and AND3_1331 (N6084,  N5407,  N4290,  N5396);
and AND3_1332 (N6085,  N5418,  N5407,  N5396);
and AND2_1333 (N6086,  N5396,  N4284);
and AND3_1334 (N6087,  N4290,  N5407,  N5396);
and AND2_1335 (N6088,  N5407,  N4290);
and AND2_1336 (N6089,  N5418,  N5407);
and AND2_1337 (N6090,  N5407,  N4290);
and AND5_1338 (N6091,  N5431,  N5462,  N5441,  N5424,  N5452);
and AND2_1339 (N6094,  N5424,  N4298);
and AND3_1340 (N6095,  N5431,  N5424,  N4301);
and AND4_1341 (N6096,  N5441,  N5424,  N4305,  N5431);
and AND5_1342 (N6097,  N5452,  N5441,  N5424,  N4310,  N5431);
and AND2_1343 (N6098,  N5431,  N4301);
and AND3_1344 (N6099,  N5441,  N4305,  N5431);
and AND4_1345 (N6100,  N5452,  N5441,  N4310,  N5431);
and AND5_1346 (N6101,  N4,  N5462,  N5441,  N5452,  N5431);
and AND2_1347 (N6102,  N4305,  N5441);
and AND3_1348 (N6103,  N5452,  N5441,  N4310);
and AND4_1349 (N6104,  N4,  N5462,  N5441,  N5452);
and AND2_1350 (N6105,  N5452,  N4310);
and AND3_1351 (N6106,  N4,  N5462,  N5452);
and AND2_1352 (N6107,  N4,  N5462);
and AND4_1353 (N6108,  N5549,  N5488,  N5477,  N5470);
and AND2_1354 (N6111,  N5477,  N4320);
and AND3_1355 (N6112,  N5488,  N4325,  N5477);
and AND3_1356 (N6113,  N5549,  N5488,  N5477);
and AND2_1357 (N6114,  N5477,  N4320);
and AND3_1358 (N6115,  N5488,  N4325,  N5477);
and AND2_1359 (N6116,  N5488,  N4325);
and AND5_1360 (N6117,  N5555,  N5536,  N5520,  N5506,  N5498);
and AND2_1361 (N6120,  N5498,  N4332);
and AND3_1362 (N6121,  N5506,  N5498,  N4336);
and AND4_1363 (N6122,  N5520,  N5498,  N4342,  N5506);
and AND5_1364 (N6123,  N5536,  N5520,  N5498,  N4349,  N5506);
and AND2_1365 (N6124,  N5506,  N4336);
and AND3_1366 (N6125,  N5520,  N4342,  N5506);
and AND4_1367 (N6126,  N5536,  N5520,  N4349,  N5506);
and AND4_1368 (N6127,  N5555,  N5520,  N5506,  N5536);
and AND2_1369 (N6128,  N5506,  N4336);
and AND3_1370 (N6129,  N5520,  N4342,  N5506);
and AND4_1371 (N6130,  N5536,  N5520,  N4349,  N5506);
and AND2_1372 (N6131,  N5520,  N4342);
and AND3_1373 (N6132,  N5536,  N5520,  N4349);
and AND3_1374 (N6133,  N5555,  N5520,  N5536);
and AND2_1375 (N6134,  N5520,  N4342);
and AND3_1376 (N6135,  N5536,  N5520,  N4349);
and AND2_1377 (N6136,  N5536,  N4349);
and AND2_1378 (N6137,  N5549,  N5488);
and AND2_1379 (N6138,  N5555,  N5536);
not NOT1_1380 (N6139,  N5573);
and AND4_1381 (N6140,  N4364,  N5573,  N5562,  N4357);
and AND3_1382 (N6143,  N5562,  N4385,  N4364);
and AND3_1383 (N6144,  N5573,  N5562,  N4364);
and AND3_1384 (N6145,  N4385,  N5562,  N4364);
and AND2_1385 (N6146,  N5562,  N4385);
and AND2_1386 (N6147,  N5573,  N5562);
and AND2_1387 (N6148,  N5562,  N4385);
and AND5_1388 (N6149,  N5264,  N4405,  N5595,  N5579,  N5606);
and AND2_1389 (N6152,  N5579,  N4067);
and AND3_1390 (N6153,  N5264,  N5579,  N4396);
and AND4_1391 (N6154,  N5595,  N5579,  N4400,  N5264);
and AND5_1392 (N6155,  N5606,  N5595,  N5579,  N4412,  N5264);
and AND3_1393 (N6156,  N5595,  N4400,  N5264);
and AND4_1394 (N6157,  N5606,  N5595,  N4412,  N5264);
and AND5_1395 (N6158,  N54,  N4405,  N5595,  N5606,  N5264);
and AND2_1396 (N6159,  N4400,  N5595);
and AND3_1397 (N6160,  N5606,  N5595,  N4412);
and AND4_1398 (N6161,  N54,  N4405,  N5595,  N5606);
and AND2_1399 (N6162,  N5606,  N4412);
and AND3_1400 (N6163,  N54,  N4405,  N5606);
nand NAND2_1401 (N6164,  N5616,  N5955);
and AND4_1402 (N6168,  N5684,  N5624,  N4425,  N4418);
and AND3_1403 (N6171,  N5624,  N4445,  N4425);
and AND3_1404 (N6172,  N5684,  N5624,  N4425);
and AND3_1405 (N6173,  N5624,  N4445,  N4425);
and AND2_1406 (N6174,  N5624,  N4445);
and AND5_1407 (N6175,  N4477,  N5671,  N5655,  N5284,  N5634);
and AND2_1408 (N6178,  N5634,  N4080);
and AND3_1409 (N6179,  N5284,  N5634,  N4456);
and AND4_1410 (N6180,  N5655,  N5634,  N4462,  N5284);
and AND5_1411 (N6181,  N5671,  N5655,  N5634,  N4469,  N5284);
and AND3_1412 (N6182,  N5655,  N4462,  N5284);
and AND4_1413 (N6183,  N5671,  N5655,  N4469,  N5284);
and AND4_1414 (N6184,  N4477,  N5655,  N5284,  N5671);
and AND3_1415 (N6185,  N5655,  N4462,  N5284);
and AND4_1416 (N6186,  N5671,  N5655,  N4469,  N5284);
and AND2_1417 (N6187,  N5655,  N4462);
and AND3_1418 (N6188,  N5671,  N5655,  N4469);
and AND3_1419 (N6189,  N4477,  N5655,  N5671);
and AND2_1420 (N6190,  N5655,  N4462);
and AND3_1421 (N6191,  N5671,  N5655,  N4469);
and AND2_1422 (N6192,  N5671,  N4469);
and AND2_1423 (N6193,  N5684,  N5624);
and AND2_1424 (N6194,  N4477,  N5671);
not NOT1_1425 (N6197,  N5692);
not NOT1_1426 (N6200,  N5696);
not NOT1_1427 (N6203,  N5703);
not NOT1_1428 (N6206,  N5707);
buf BUFF1_1429 (N6209,  N5700);
buf BUFF1_1430 (N6212,  N5700);
buf BUFF1_1431 (N6215,  N5711);
buf BUFF1_1432 (N6218,  N5711);
nand NAND2_1433 (N6221,  N5049,  N6023);
not NOT1_1434 (N6234,  N5756);
nand NAND2_1435 (N6235,  N5756,  N6044);
buf BUFF1_1436 (N6238,  N5462);
buf BUFF1_1437 (N6241,  N5389);
buf BUFF1_1438 (N6244,  N5389);
buf BUFF1_1439 (N6247,  N5396);
buf BUFF1_1440 (N6250,  N5396);
buf BUFF1_1441 (N6253,  N5407);
buf BUFF1_1442 (N6256,  N5407);
buf BUFF1_1443 (N6259,  N5424);
buf BUFF1_1444 (N6262,  N5431);
buf BUFF1_1445 (N6265,  N5441);
buf BUFF1_1446 (N6268,  N5452);
buf BUFF1_1447 (N6271,  N5549);
buf BUFF1_1448 (N6274,  N5488);
buf BUFF1_1449 (N6277,  N5470);
buf BUFF1_1450 (N6280,  N5477);
buf BUFF1_1451 (N6283,  N5549);
buf BUFF1_1452 (N6286,  N5488);
buf BUFF1_1453 (N6289,  N5470);
buf BUFF1_1454 (N6292,  N5477);
buf BUFF1_1455 (N6295,  N5555);
buf BUFF1_1456 (N6298,  N5536);
buf BUFF1_1457 (N6301,  N5498);
buf BUFF1_1458 (N6304,  N5520);
buf BUFF1_1459 (N6307,  N5506);
buf BUFF1_1460 (N6310,  N5506);
buf BUFF1_1461 (N6313,  N5555);
buf BUFF1_1462 (N6316,  N5536);
buf BUFF1_1463 (N6319,  N5498);
buf BUFF1_1464 (N6322,  N5520);
buf BUFF1_1465 (N6325,  N5562);
buf BUFF1_1466 (N6328,  N5562);
buf BUFF1_1467 (N6331,  N5579);
buf BUFF1_1468 (N6335,  N5595);
buf BUFF1_1469 (N6338,  N5606);
buf BUFF1_1470 (N6341,  N5684);
buf BUFF1_1471 (N6344,  N5624);
buf BUFF1_1472 (N6347,  N5684);
buf BUFF1_1473 (N6350,  N5624);
buf BUFF1_1474 (N6353,  N5671);
buf BUFF1_1475 (N6356,  N5634);
buf BUFF1_1476 (N6359,  N5655);
buf BUFF1_1477 (N6364,  N5671);
buf BUFF1_1478 (N6367,  N5634);
buf BUFF1_1479 (N6370,  N5655);
not NOT1_1480 (N6373,  N5736);
not NOT1_1481 (N6374,  N5739);
not NOT1_1482 (N6375,  N5742);
not NOT1_1483 (N6376,  N5745);
nand NAND2_1484 (N6377,  N4243,  N6065);
nand NAND2_1485 (N6378,  N5236,  N6068);
or OR4_1486 (N6382,  N4268,  N6071,  N6072,  N6073);
or OR4_1487 (N6386,  N3968,  N5065,  N5066,  N6074);
or OR4_1488 (N6388,  N4271,  N6075,  N6076,  N6077);
or OR4_1489 (N6392,  N3968,  N5067,  N5068,  N6078);
or OR5_1490 (N6397,  N4297,  N6094,  N6095,  N6096,  N6097);
or OR2_1491 (N6411,  N4320,  N6116);
or OR5_1492 (N6415,  N4331,  N6120,  N6121,  N6122,  N6123);
or OR2_1493 (N6419,  N4342,  N6136);
or OR5_1494 (N6427,  N4392,  N6152,  N6153,  N6154,  N6155);
not NOT1_1495 (N6434,  N6048);
or OR2_1496 (N6437,  N4440,  N6174);
or OR5_1497 (N6441,  N4451,  N6178,  N6179,  N6180,  N6181);
or OR2_1498 (N6445,  N4462,  N6192);
not NOT1_1499 (N6448,  N6051);
not NOT1_1500 (N6449,  N6054);
nand NAND2_1501 (N6466,  N6221,  N6024);
not NOT1_1502 (N6469,  N6031);
not NOT1_1503 (N6470,  N6034);
not NOT1_1504 (N6471,  N6037);
not NOT1_1505 (N6472,  N6040);
and AND3_1506 (N6473,  N5315,  N4524,  N6031);
and AND3_1507 (N6474,  N6025,  N5150,  N6034);
and AND3_1508 (N6475,  N5324,  N4532,  N6037);
and AND3_1509 (N6476,  N6028,  N5157,  N6040);
nand NAND2_1510 (N6477,  N5385,  N6234);
nand NAND2_1511 (N6478,  N6045,  N132);
or OR4_1512 (N6482,  N4280,  N6083,  N6084,  N6085);
nor NOR3_1513 (N6486,  N4280,  N6086,  N6087);
or OR3_1514 (N6490,  N4284,  N6088,  N6089);
nor NOR2_1515 (N6494,  N4284,  N6090);
or OR5_1516 (N6500,  N4298,  N6098,  N6099,  N6100,  N6101);
or OR4_1517 (N6504,  N4301,  N6102,  N6103,  N6104);
or OR3_1518 (N6508,  N4305,  N6105,  N6106);
or OR2_1519 (N6512,  N4310,  N6107);
or OR4_1520 (N6516,  N4316,  N6111,  N6112,  N6113);
nor NOR3_1521 (N6526,  N4316,  N6114,  N6115);
or OR4_1522 (N6536,  N4336,  N6131,  N6132,  N6133);
or OR5_1523 (N6539,  N4332,  N6124,  N6125,  N6126,  N6127);
nor NOR3_1524 (N6553,  N4336,  N6134,  N6135);
nor NOR4_1525 (N6556,  N4332,  N6128,  N6129,  N6130);
or OR4_1526 (N6566,  N4375,  N5117,  N6143,  N6144);
nor NOR3_1527 (N6569,  N4375,  N5118,  N6145);
or OR3_1528 (N6572,  N4379,  N6146,  N6147);
nor NOR2_1529 (N6575,  N4379,  N6148);
or OR5_1530 (N6580,  N4067,  N5954,  N6156,  N6157,  N6158);
or OR4_1531 (N6584,  N4396,  N6159,  N6160,  N6161);
or OR3_1532 (N6587,  N4400,  N6162,  N6163);
or OR4_1533 (N6592,  N4436,  N5132,  N6171,  N6172);
nor NOR3_1534 (N6599,  N4436,  N5133,  N6173);
or OR4_1535 (N6606,  N4456,  N6187,  N6188,  N6189);
or OR5_1536 (N6609,  N4080,  N6005,  N6182,  N6183,  N6184);
nor NOR3_1537 (N6619,  N4456,  N6190,  N6191);
nor NOR4_1538 (N6622,  N4080,  N6006,  N6185,  N6186);
nand NAND2_1539 (N6630,  N5739,  N6373);
nand NAND2_1540 (N6631,  N5736,  N6374);
nand NAND2_1541 (N6632,  N5745,  N6375);
nand NAND2_1542 (N6633,  N5742,  N6376);
nand NAND2_1543 (N6634,  N6377,  N6066);
nand NAND2_1544 (N6637,  N6069,  N6378);
not NOT1_1545 (N6640,  N6164);
and AND2_1546 (N6641,  N6108,  N6117);
and AND2_1547 (N6643,  N6140,  N6149);
and AND2_1548 (N6646,  N6168,  N6175);
and AND2_1549 (N6648,  N6080,  N6091);
nand NAND2_1550 (N6650,  N6238,  N2637);
not NOT1_1551 (N6651,  N6238);
not NOT1_1552 (N6653,  N6241);
not NOT1_1553 (N6655,  N6244);
not NOT1_1554 (N6657,  N6247);
not NOT1_1555 (N6659,  N6250);
nand NAND2_1556 (N6660,  N6253,  N5087);
not NOT1_1557 (N6661,  N6253);
nand NAND2_1558 (N6662,  N6256,  N5469);
not NOT1_1559 (N6663,  N6256);
and AND2_1560 (N6664,  N6091,  N4);
not NOT1_1561 (N6666,  N6259);
not NOT1_1562 (N6668,  N6262);
not NOT1_1563 (N6670,  N6265);
not NOT1_1564 (N6672,  N6268);
not NOT1_1565 (N6675,  N6117);
not NOT1_1566 (N6680,  N6280);
not NOT1_1567 (N6681,  N6292);
not NOT1_1568 (N6682,  N6307);
not NOT1_1569 (N6683,  N6310);
nand NAND2_1570 (N6689,  N6325,  N5120);
not NOT1_1571 (N6690,  N6325);
nand NAND2_1572 (N6691,  N6328,  N5622);
not NOT1_1573 (N6692,  N6328);
and AND2_1574 (N6693,  N6149,  N54);
not NOT1_1575 (N6695,  N6331);
not NOT1_1576 (N6698,  N6335);
nand NAND2_1577 (N6699,  N6338,  N5956);
not NOT1_1578 (N6700,  N6338);
not NOT1_1579 (N6703,  N6175);
not NOT1_1580 (N6708,  N6209);
not NOT1_1581 (N6709,  N6212);
not NOT1_1582 (N6710,  N6215);
not NOT1_1583 (N6711,  N6218);
and AND3_1584 (N6712,  N5696,  N5692,  N6209);
and AND3_1585 (N6713,  N6200,  N6197,  N6212);
and AND3_1586 (N6714,  N5707,  N5703,  N6215);
and AND3_1587 (N6715,  N6206,  N6203,  N6218);
buf BUFF1_1588 (N6716,  N6466);
and AND3_1589 (N6718,  N6164,  N1777,  N3130);
and AND3_1590 (N6719,  N5150,  N5315,  N6469);
and AND3_1591 (N6720,  N4524,  N6025,  N6470);
and AND3_1592 (N6721,  N5157,  N5324,  N6471);
and AND3_1593 (N6722,  N4532,  N6028,  N6472);
nand NAND2_1594 (N6724,  N6477,  N6235);
not NOT1_1595 (N6739,  N6271);
not NOT1_1596 (N6740,  N6274);
not NOT1_1597 (N6741,  N6277);
not NOT1_1598 (N6744,  N6283);
not NOT1_1599 (N6745,  N6286);
not NOT1_1600 (N6746,  N6289);
not NOT1_1601 (N6751,  N6295);
not NOT1_1602 (N6752,  N6298);
not NOT1_1603 (N6753,  N6301);
not NOT1_1604 (N6754,  N6304);
not NOT1_1605 (N6755,  N6322);
not NOT1_1606 (N6760,  N6313);
not NOT1_1607 (N6761,  N6316);
not NOT1_1608 (N6762,  N6319);
not NOT1_1609 (N6772,  N6341);
not NOT1_1610 (N6773,  N6344);
not NOT1_1611 (N6776,  N6347);
not NOT1_1612 (N6777,  N6350);
not NOT1_1613 (N6782,  N6353);
not NOT1_1614 (N6783,  N6356);
not NOT1_1615 (N6784,  N6359);
not NOT1_1616 (N6785,  N6370);
not NOT1_1617 (N6790,  N6364);
not NOT1_1618 (N6791,  N6367);
nand NAND2_1619 (N6792,  N6630,  N6631);
nand NAND2_1620 (N6795,  N6632,  N6633);
and AND2_1621 (N6801,  N6108,  N6415);
and AND2_1622 (N6802,  N6427,  N6140);
and AND2_1623 (N6803,  N6397,  N6080);
and AND2_1624 (N6804,  N6168,  N6441);
not NOT1_1625 (N6805,  N6466);
nand NAND2_1626 (N6806,  N1851,  N6651);
not NOT1_1627 (N6807,  N6482);
nand NAND2_1628 (N6808,  N6482,  N6653);
not NOT1_1629 (N6809,  N6486);
nand NAND2_1630 (N6810,  N6486,  N6655);
not NOT1_1631 (N6811,  N6490);
nand NAND2_1632 (N6812,  N6490,  N6657);
not NOT1_1633 (N6813,  N6494);
nand NAND2_1634 (N6814,  N6494,  N6659);
nand NAND2_1635 (N6815,  N4575,  N6661);
nand NAND2_1636 (N6816,  N5169,  N6663);
or OR2_1637 (N6817,  N6397,  N6664);
not NOT1_1638 (N6823,  N6500);
nand NAND2_1639 (N6824,  N6500,  N6666);
not NOT1_1640 (N6825,  N6504);
nand NAND2_1641 (N6826,  N6504,  N6668);
not NOT1_1642 (N6827,  N6508);
nand NAND2_1643 (N6828,  N6508,  N6670);
not NOT1_1644 (N6829,  N6512);
nand NAND2_1645 (N6830,  N6512,  N6672);
not NOT1_1646 (N6831,  N6415);
not NOT1_1647 (N6834,  N6566);
nand NAND2_1648 (N6835,  N6566,  N5618);
not NOT1_1649 (N6836,  N6569);
nand NAND2_1650 (N6837,  N6569,  N5619);
not NOT1_1651 (N6838,  N6572);
nand NAND2_1652 (N6839,  N6572,  N5620);
not NOT1_1653 (N6840,  N6575);
nand NAND2_1654 (N6841,  N6575,  N5621);
nand NAND2_1655 (N6842,  N4627,  N6690);
nand NAND2_1656 (N6843,  N5195,  N6692);
or OR2_1657 (N6844,  N6427,  N6693);
not NOT1_1658 (N6850,  N6580);
nand NAND2_1659 (N6851,  N6580,  N6695);
not NOT1_1660 (N6852,  N6584);
nand NAND2_1661 (N6853,  N6584,  N6434);
not NOT1_1662 (N6854,  N6587);
nand NAND2_1663 (N6855,  N6587,  N6698);
nand NAND2_1664 (N6856,  N5346,  N6700);
not NOT1_1665 (N6857,  N6441);
and AND3_1666 (N6860,  N6197,  N5696,  N6708);
and AND3_1667 (N6861,  N5692,  N6200,  N6709);
and AND3_1668 (N6862,  N6203,  N5707,  N6710);
and AND3_1669 (N6863,  N5703,  N6206,  N6711);
or OR3_1670 (N6866,  N4197,  N6718,  N3785);
nor NOR2_1671 (N6872,  N6719,  N6473);
nor NOR2_1672 (N6873,  N6720,  N6474);
nor NOR2_1673 (N6874,  N6721,  N6475);
nor NOR2_1674 (N6875,  N6722,  N6476);
not NOT1_1675 (N6876,  N6637);
buf BUFF1_1676 (N6877,  N6724);
and AND2_1677 (N6879,  N6045,  N6478);
and AND2_1678 (N6880,  N6478,  N132);
or OR2_1679 (N6881,  N6411,  N6137);
not NOT1_1680 (N6884,  N6516);
not NOT1_1681 (N6885,  N6411);
not NOT1_1682 (N6888,  N6526);
not NOT1_1683 (N6889,  N6536);
nand NAND2_1684 (N6890,  N6536,  N5176);
or OR2_1685 (N6891,  N6419,  N6138);
not NOT1_1686 (N6894,  N6539);
not NOT1_1687 (N6895,  N6553);
nand NAND2_1688 (N6896,  N6553,  N5728);
not NOT1_1689 (N6897,  N6419);
not NOT1_1690 (N6900,  N6556);
or OR2_1691 (N6901,  N6437,  N6193);
not NOT1_1692 (N6904,  N6592);
not NOT1_1693 (N6905,  N6437);
not NOT1_1694 (N6908,  N6599);
or OR2_1695 (N6909,  N6445,  N6194);
not NOT1_1696 (N6912,  N6606);
not NOT1_1697 (N6913,  N6609);
not NOT1_1698 (N6914,  N6619);
nand NAND2_1699 (N6915,  N6619,  N5734);
not NOT1_1700 (N6916,  N6445);
not NOT1_1701 (N6919,  N6622);
not NOT1_1702 (N6922,  N6634);
nand NAND2_1703 (N6923,  N6634,  N6067);
or OR2_1704 (N6924,  N6382,  N6801);
or OR2_1705 (N6925,  N6386,  N6802);
or OR2_1706 (N6926,  N6388,  N6803);
or OR2_1707 (N6927,  N6392,  N6804);
not NOT1_1708 (N6930,  N6724);
nand NAND2_1709 (N6932,  N6650,  N6806);
nand NAND2_1710 (N6935,  N6241,  N6807);
nand NAND2_1711 (N6936,  N6244,  N6809);
nand NAND2_1712 (N6937,  N6247,  N6811);
nand NAND2_1713 (N6938,  N6250,  N6813);
nand NAND2_1714 (N6939,  N6660,  N6815);
nand NAND2_1715 (N6940,  N6662,  N6816);
nand NAND2_1716 (N6946,  N6259,  N6823);
nand NAND2_1717 (N6947,  N6262,  N6825);
nand NAND2_1718 (N6948,  N6265,  N6827);
nand NAND2_1719 (N6949,  N6268,  N6829);
nand NAND2_1720 (N6953,  N5183,  N6834);
nand NAND2_1721 (N6954,  N5186,  N6836);
nand NAND2_1722 (N6955,  N5189,  N6838);
nand NAND2_1723 (N6956,  N5192,  N6840);
nand NAND2_1724 (N6957,  N6689,  N6842);
nand NAND2_1725 (N6958,  N6691,  N6843);
nand NAND2_1726 (N6964,  N6331,  N6850);
nand NAND2_1727 (N6965,  N6048,  N6852);
nand NAND2_1728 (N6966,  N6335,  N6854);
nand NAND2_1729 (N6967,  N6699,  N6856);
nor NOR2_1730 (N6973,  N6860,  N6712);
nor NOR2_1731 (N6974,  N6861,  N6713);
nor NOR2_1732 (N6975,  N6862,  N6714);
nor NOR2_1733 (N6976,  N6863,  N6715);
not NOT1_1734 (N6977,  N6792);
not NOT1_1735 (N6978,  N6795);
or OR2_1736 (N6979,  N6879,  N6880);
nand NAND2_1737 (N6987,  N4608,  N6889);
nand NAND2_1738 (N6990,  N5177,  N6895);
nand NAND2_1739 (N6999,  N5217,  N6914);
nand NAND2_1740 (N7002,  N5377,  N6922);
nand NAND2_1741 (N7003,  N6873,  N6872);
nand NAND2_1742 (N7006,  N6875,  N6874);
and AND3_1743 (N7011,  N6866,  N2681,  N2692);
and AND3_1744 (N7012,  N6866,  N2756,  N2767);
and AND3_1745 (N7013,  N6866,  N2779,  N2790);
not NOT1_1746 (N7015,  N6866);
and AND3_1747 (N7016,  N6866,  N2801,  N2812);
nand NAND2_1748 (N7018,  N6935,  N6808);
nand NAND2_1749 (N7019,  N6936,  N6810);
nand NAND2_1750 (N7020,  N6937,  N6812);
nand NAND2_1751 (N7021,  N6938,  N6814);
not NOT1_1752 (N7022,  N6939);
not NOT1_1753 (N7023,  N6817);
nand NAND2_1754 (N7028,  N6946,  N6824);
nand NAND2_1755 (N7031,  N6947,  N6826);
nand NAND2_1756 (N7034,  N6948,  N6828);
nand NAND2_1757 (N7037,  N6949,  N6830);
and AND2_1758 (N7040,  N6817,  N6079);
and AND2_1759 (N7041,  N6831,  N6675);
nand NAND2_1760 (N7044,  N6953,  N6835);
nand NAND2_1761 (N7045,  N6954,  N6837);
nand NAND2_1762 (N7046,  N6955,  N6839);
nand NAND2_1763 (N7047,  N6956,  N6841);
not NOT1_1764 (N7048,  N6957);
not NOT1_1765 (N7049,  N6844);
nand NAND2_1766 (N7054,  N6964,  N6851);
nand NAND2_1767 (N7057,  N6965,  N6853);
nand NAND2_1768 (N7060,  N6966,  N6855);
and AND2_1769 (N7064,  N6844,  N6139);
and AND2_1770 (N7065,  N6857,  N6703);
not NOT1_1771 (N7072,  N6881);
nand NAND2_1772 (N7073,  N6881,  N5172);
not NOT1_1773 (N7074,  N6885);
nand NAND2_1774 (N7075,  N6885,  N5727);
nand NAND2_1775 (N7076,  N6890,  N6987);
not NOT1_1776 (N7079,  N6891);
nand NAND2_1777 (N7080,  N6896,  N6990);
not NOT1_1778 (N7083,  N6897);
not NOT1_1779 (N7084,  N6901);
nand NAND2_1780 (N7085,  N6901,  N5198);
not NOT1_1781 (N7086,  N6905);
nand NAND2_1782 (N7087,  N6905,  N5731);
not NOT1_1783 (N7088,  N6909);
nand NAND2_1784 (N7089,  N6909,  N6912);
nand NAND2_1785 (N7090,  N6915,  N6999);
not NOT1_1786 (N7093,  N6916);
nand NAND2_1787 (N7094,  N6974,  N6973);
nand NAND2_1788 (N7097,  N6976,  N6975);
nand NAND2_1789 (N7101,  N7002,  N6923);
not NOT1_1790 (N7105,  N6932);
not NOT1_1791 (N7110,  N6967);
and AND3_1792 (N7114,  N6979,  N603,  N1755);
not NOT1_1793 (N7115,  N7019);
not NOT1_1794 (N7116,  N7021);
and AND2_1795 (N7125,  N6817,  N7018);
and AND2_1796 (N7126,  N6817,  N7020);
and AND2_1797 (N7127,  N6817,  N7022);
not NOT1_1798 (N7130,  N7045);
not NOT1_1799 (N7131,  N7047);
and AND2_1800 (N7139,  N6844,  N7044);
and AND2_1801 (N7140,  N6844,  N7046);
and AND2_1802 (N7141,  N6844,  N7048);
and AND3_1803 (N7146,  N6932,  N1761,  N3108);
and AND3_1804 (N7147,  N6967,  N1777,  N3130);
not NOT1_1805 (N7149,  N7003);
not NOT1_1806 (N7150,  N7006);
nand NAND2_1807 (N7151,  N7006,  N6876);
nand NAND2_1808 (N7152,  N4605,  N7072);
nand NAND2_1809 (N7153,  N5173,  N7074);
nand NAND2_1810 (N7158,  N4646,  N7084);
nand NAND2_1811 (N7159,  N5205,  N7086);
nand NAND2_1812 (N7160,  N6606,  N7088);
not NOT1_1813 (N7166,  N7037);
not NOT1_1814 (N7167,  N7034);
not NOT1_1815 (N7168,  N7031);
not NOT1_1816 (N7169,  N7028);
not NOT1_1817 (N7170,  N7060);
not NOT1_1818 (N7171,  N7057);
not NOT1_1819 (N7172,  N7054);
and AND2_1820 (N7173,  N7115,  N7023);
and AND2_1821 (N7174,  N7116,  N7023);
and AND2_1822 (N7175,  N6940,  N7023);
and AND2_1823 (N7176,  N5418,  N7023);
not NOT1_1824 (N7177,  N7041);
and AND2_1825 (N7178,  N7130,  N7049);
and AND2_1826 (N7179,  N7131,  N7049);
and AND2_1827 (N7180,  N6958,  N7049);
and AND2_1828 (N7181,  N5573,  N7049);
not NOT1_1829 (N7182,  N7065);
not NOT1_1830 (N7183,  N7094);
nand NAND2_1831 (N7184,  N7094,  N6977);
not NOT1_1832 (N7185,  N7097);
nand NAND2_1833 (N7186,  N7097,  N6978);
and AND3_1834 (N7187,  N7037,  N1761,  N3108);
and AND3_1835 (N7188,  N7034,  N1761,  N3108);
and AND3_1836 (N7189,  N7031,  N1761,  N3108);
or OR3_1837 (N7190,  N4956,  N7146,  N3781);
and AND3_1838 (N7196,  N7060,  N1777,  N3130);
and AND3_1839 (N7197,  N7057,  N1777,  N3130);
or OR3_1840 (N7198,  N4960,  N7147,  N3786);
nand NAND2_1841 (N7204,  N7101,  N7149);
not NOT1_1842 (N7205,  N7101);
nand NAND2_1843 (N7206,  N6637,  N7150);
and AND3_1844 (N7207,  N7028,  N1793,  N3158);
and AND3_1845 (N7208,  N7054,  N1807,  N3180);
nand NAND2_1846 (N7209,  N7073,  N7152);
nand NAND2_1847 (N7212,  N7075,  N7153);
not NOT1_1848 (N7215,  N7076);
nand NAND2_1849 (N7216,  N7076,  N7079);
not NOT1_1850 (N7217,  N7080);
nand NAND2_1851 (N7218,  N7080,  N7083);
nand NAND2_1852 (N7219,  N7085,  N7158);
nand NAND2_1853 (N7222,  N7087,  N7159);
nand NAND2_1854 (N7225,  N7089,  N7160);
not NOT1_1855 (N7228,  N7090);
nand NAND2_1856 (N7229,  N7090,  N7093);
or OR2_1857 (N7236,  N7173,  N7125);
or OR2_1858 (N7239,  N7174,  N7126);
or OR2_1859 (N7242,  N7175,  N7127);
or OR2_1860 (N7245,  N7176,  N7040);
or OR2_1861 (N7250,  N7178,  N7139);
or OR2_1862 (N7257,  N7179,  N7140);
or OR2_1863 (N7260,  N7180,  N7141);
or OR2_1864 (N7263,  N7181,  N7064);
nand NAND2_1865 (N7268,  N6792,  N7183);
nand NAND2_1866 (N7269,  N6795,  N7185);
or OR3_1867 (N7270,  N4957,  N7187,  N3782);
or OR3_1868 (N7276,  N4958,  N7188,  N3783);
or OR3_1869 (N7282,  N4959,  N7189,  N3784);
or OR3_1870 (N7288,  N4961,  N7196,  N3787);
or OR3_1871 (N7294,  N3998,  N7197,  N3788);
nand NAND2_1872 (N7300,  N7003,  N7205);
nand NAND2_1873 (N7301,  N7206,  N7151);
or OR3_1874 (N7304,  N4980,  N7207,  N3800);
or OR3_1875 (N7310,  N4984,  N7208,  N3805);
nand NAND2_1876 (N7320,  N6891,  N7215);
nand NAND2_1877 (N7321,  N6897,  N7217);
nand NAND2_1878 (N7328,  N6916,  N7228);
and AND3_1879 (N7338,  N7190,  N1185,  N2692);
and AND3_1880 (N7339,  N7198,  N2681,  N2692);
and AND3_1881 (N7340,  N7190,  N1247,  N2767);
and AND3_1882 (N7341,  N7198,  N2756,  N2767);
and AND3_1883 (N7342,  N7190,  N1327,  N2790);
and AND3_1884 (N7349,  N7198,  N2779,  N2790);
and AND3_1885 (N7357,  N7198,  N2801,  N2812);
not NOT1_1886 (N7363,  N7198);
and AND3_1887 (N7364,  N7190,  N1351,  N2812);
not NOT1_1888 (N7365,  N7190);
nand NAND2_1889 (N7394,  N7268,  N7184);
nand NAND2_1890 (N7397,  N7269,  N7186);
nand NAND2_1891 (N7402,  N7204,  N7300);
not NOT1_1892 (N7405,  N7209);
nand NAND2_1893 (N7406,  N7209,  N6884);
not NOT1_1894 (N7407,  N7212);
nand NAND2_1895 (N7408,  N7212,  N6888);
nand NAND2_1896 (N7409,  N7320,  N7216);
nand NAND2_1897 (N7412,  N7321,  N7218);
not NOT1_1898 (N7415,  N7219);
nand NAND2_1899 (N7416,  N7219,  N6904);
not NOT1_1900 (N7417,  N7222);
nand NAND2_1901 (N7418,  N7222,  N6908);
not NOT1_1902 (N7419,  N7225);
nand NAND2_1903 (N7420,  N7225,  N6913);
nand NAND2_1904 (N7421,  N7328,  N7229);
not NOT1_1905 (N7424,  N7245);
not NOT1_1906 (N7425,  N7242);
not NOT1_1907 (N7426,  N7239);
not NOT1_1908 (N7427,  N7236);
not NOT1_1909 (N7428,  N7263);
not NOT1_1910 (N7429,  N7260);
not NOT1_1911 (N7430,  N7257);
not NOT1_1912 (N7431,  N7250);
not NOT1_1913 (N7432,  N7250);
and AND3_1914 (N7433,  N7310,  N2653,  N2664);
and AND3_1915 (N7434,  N7304,  N1161,  N2664);
or OR4_1916 (N7435,  N7011,  N7338,  N3621,  N2591);
and AND3_1917 (N7436,  N7270,  N1185,  N2692);
and AND3_1918 (N7437,  N7288,  N2681,  N2692);
and AND3_1919 (N7438,  N7276,  N1185,  N2692);
and AND3_1920 (N7439,  N7294,  N2681,  N2692);
and AND3_1921 (N7440,  N7282,  N1185,  N2692);
and AND3_1922 (N7441,  N7310,  N2728,  N2739);
and AND3_1923 (N7442,  N7304,  N1223,  N2739);
or OR4_1924 (N7443,  N7012,  N7340,  N3632,  N2600);
and AND3_1925 (N7444,  N7270,  N1247,  N2767);
and AND3_1926 (N7445,  N7288,  N2756,  N2767);
and AND3_1927 (N7446,  N7276,  N1247,  N2767);
and AND3_1928 (N7447,  N7294,  N2756,  N2767);
and AND3_1929 (N7448,  N7282,  N1247,  N2767);
or OR4_1930 (N7449,  N7013,  N7342,  N3641,  N2605);
and AND3_1931 (N7450,  N7310,  N3041,  N3052);
and AND3_1932 (N7451,  N7304,  N1697,  N3052);
and AND3_1933 (N7452,  N7294,  N2779,  N2790);
and AND3_1934 (N7453,  N7282,  N1327,  N2790);
and AND3_1935 (N7454,  N7288,  N2779,  N2790);
and AND3_1936 (N7455,  N7276,  N1327,  N2790);
and AND3_1937 (N7456,  N7270,  N1327,  N2790);
and AND3_1938 (N7457,  N7310,  N3075,  N3086);
and AND3_1939 (N7458,  N7304,  N1731,  N3086);
and AND3_1940 (N7459,  N7294,  N2801,  N2812);
and AND3_1941 (N7460,  N7282,  N1351,  N2812);
and AND3_1942 (N7461,  N7288,  N2801,  N2812);
and AND3_1943 (N7462,  N7276,  N1351,  N2812);
and AND3_1944 (N7463,  N7270,  N1351,  N2812);
and AND3_1945 (N7464,  N7250,  N603,  N599);
not NOT1_1946 (N7465,  N7310);
not NOT1_1947 (N7466,  N7294);
not NOT1_1948 (N7467,  N7288);
not NOT1_1949 (N7468,  N7301);
or OR4_1950 (N7469,  N7016,  N7364,  N3660,  N2626);
not NOT1_1951 (N7470,  N7304);
not NOT1_1952 (N7471,  N7282);
not NOT1_1953 (N7472,  N7276);
not NOT1_1954 (N7473,  N7270);
buf BUFF1_1955 (N7474,  N7394);
buf BUFF1_1956 (N7476,  N7397);
and AND2_1957 (N7479,  N7301,  N3068);
and AND3_1958 (N7481,  N7245,  N1793,  N3158);
and AND3_1959 (N7482,  N7242,  N1793,  N3158);
and AND3_1960 (N7483,  N7239,  N1793,  N3158);
and AND3_1961 (N7484,  N7236,  N1793,  N3158);
and AND3_1962 (N7485,  N7263,  N1807,  N3180);
and AND3_1963 (N7486,  N7260,  N1807,  N3180);
and AND3_1964 (N7487,  N7257,  N1807,  N3180);
and AND3_1965 (N7488,  N7250,  N1807,  N3180);
nand NAND2_1966 (N7489,  N6979,  N7250);
nand NAND2_1967 (N7492,  N6516,  N7405);
nand NAND2_1968 (N7493,  N6526,  N7407);
nand NAND2_1969 (N7498,  N6592,  N7415);
nand NAND2_1970 (N7499,  N6599,  N7417);
nand NAND2_1971 (N7500,  N6609,  N7419);
and AND9_1972 (N7503,  N7105,  N7166,  N7167,  N7168,  N7169,  N7424,  N7425,  N7426,  N7427);
and AND9_1973 (N7504,  N6640,  N7110,  N7170,  N7171,  N7172,  N7428,  N7429,  N7430,  N7431);
or OR4_1974 (N7505,  N7433,  N7434,  N3616,  N2585);
and AND2_1975 (N7506,  N7435,  N2675);
or OR4_1976 (N7507,  N7339,  N7436,  N3622,  N2592);
or OR4_1977 (N7508,  N7437,  N7438,  N3623,  N2593);
or OR4_1978 (N7509,  N7439,  N7440,  N3624,  N2594);
or OR4_1979 (N7510,  N7441,  N7442,  N3627,  N2595);
and AND2_1980 (N7511,  N7443,  N2750);
or OR4_1981 (N7512,  N7341,  N7444,  N3633,  N2601);
or OR4_1982 (N7513,  N7445,  N7446,  N3634,  N2602);
or OR4_1983 (N7514,  N7447,  N7448,  N3635,  N2603);
or OR4_1984 (N7515,  N7450,  N7451,  N3646,  N2610);
or OR4_1985 (N7516,  N7452,  N7453,  N3647,  N2611);
or OR4_1986 (N7517,  N7454,  N7455,  N3648,  N2612);
or OR4_1987 (N7518,  N7349,  N7456,  N3649,  N2613);
or OR4_1988 (N7519,  N7457,  N7458,  N3654,  N2618);
or OR4_1989 (N7520,  N7459,  N7460,  N3655,  N2619);
or OR4_1990 (N7521,  N7461,  N7462,  N3656,  N2620);
or OR4_1991 (N7522,  N7357,  N7463,  N3657,  N2621);
or OR4_1992 (N7525,  N4741,  N7114,  N2624,  N7464);
and AND3_1993 (N7526,  N7468,  N3119,  N3130);
not NOT1_1994 (N7527,  N7394);
not NOT1_1995 (N7528,  N7397);
not NOT1_1996 (N7529,  N7402);
and AND2_1997 (N7530,  N7402,  N3068);
or OR3_1998 (N7531,  N4981,  N7481,  N3801);
or OR3_1999 (N7537,  N4982,  N7482,  N3802);
or OR3_2000 (N7543,  N4983,  N7483,  N3803);
or OR3_2001 (N7549,  N5165,  N7484,  N3804);
or OR3_2002 (N7555,  N4985,  N7485,  N3806);
or OR3_2003 (N7561,  N4986,  N7486,  N3807);
or OR3_2004 (N7567,  N4547,  N7487,  N3808);
or OR3_2005 (N7573,  N4987,  N7488,  N3809);
nand NAND2_2006 (N7579,  N7492,  N7406);
nand NAND2_2007 (N7582,  N7493,  N7408);
not NOT1_2008 (N7585,  N7409);
nand NAND2_2009 (N7586,  N7409,  N6894);
not NOT1_2010 (N7587,  N7412);
nand NAND2_2011 (N7588,  N7412,  N6900);
nand NAND2_2012 (N7589,  N7498,  N7416);
nand NAND2_2013 (N7592,  N7499,  N7418);
nand NAND2_2014 (N7595,  N7500,  N7420);
not NOT1_2015 (N7598,  N7421);
nand NAND2_2016 (N7599,  N7421,  N6919);
and AND2_2017 (N7600,  N7505,  N2647);
and AND2_2018 (N7601,  N7507,  N2675);
and AND2_2019 (N7602,  N7508,  N2675);
and AND2_2020 (N7603,  N7509,  N2675);
and AND2_2021 (N7604,  N7510,  N2722);
and AND2_2022 (N7605,  N7512,  N2750);
and AND2_2023 (N7606,  N7513,  N2750);
and AND2_2024 (N7607,  N7514,  N2750);
and AND2_2025 (N7624,  N6979,  N7489);
and AND2_2026 (N7625,  N7489,  N7250);
and AND2_2027 (N7626,  N1149,  N7525);
and AND5_2028 (N7631,  N562,  N7527,  N7528,  N6805,  N6930);
and AND3_2029 (N7636,  N7529,  N3097,  N3108);
nand NAND2_2030 (N7657,  N6539,  N7585);
nand NAND2_2031 (N7658,  N6556,  N7587);
nand NAND2_2032 (N7665,  N6622,  N7598);
and AND3_2033 (N7666,  N7555,  N2653,  N2664);
and AND3_2034 (N7667,  N7531,  N1161,  N2664);
and AND3_2035 (N7668,  N7561,  N2653,  N2664);
and AND3_2036 (N7669,  N7537,  N1161,  N2664);
and AND3_2037 (N7670,  N7567,  N2653,  N2664);
and AND3_2038 (N7671,  N7543,  N1161,  N2664);
and AND3_2039 (N7672,  N7573,  N2653,  N2664);
and AND3_2040 (N7673,  N7549,  N1161,  N2664);
and AND3_2041 (N7674,  N7555,  N2728,  N2739);
and AND3_2042 (N7675,  N7531,  N1223,  N2739);
and AND3_2043 (N7676,  N7561,  N2728,  N2739);
and AND3_2044 (N7677,  N7537,  N1223,  N2739);
and AND3_2045 (N7678,  N7567,  N2728,  N2739);
and AND3_2046 (N7679,  N7543,  N1223,  N2739);
and AND3_2047 (N7680,  N7573,  N2728,  N2739);
and AND3_2048 (N7681,  N7549,  N1223,  N2739);
and AND3_2049 (N7682,  N7573,  N3075,  N3086);
and AND3_2050 (N7683,  N7549,  N1731,  N3086);
and AND3_2051 (N7684,  N7573,  N3041,  N3052);
and AND3_2052 (N7685,  N7549,  N1697,  N3052);
and AND3_2053 (N7686,  N7567,  N3041,  N3052);
and AND3_2054 (N7687,  N7543,  N1697,  N3052);
and AND3_2055 (N7688,  N7561,  N3041,  N3052);
and AND3_2056 (N7689,  N7537,  N1697,  N3052);
and AND3_2057 (N7690,  N7555,  N3041,  N3052);
and AND3_2058 (N7691,  N7531,  N1697,  N3052);
and AND3_2059 (N7692,  N7567,  N3075,  N3086);
and AND3_2060 (N7693,  N7543,  N1731,  N3086);
and AND3_2061 (N7694,  N7561,  N3075,  N3086);
and AND3_2062 (N7695,  N7537,  N1731,  N3086);
and AND3_2063 (N7696,  N7555,  N3075,  N3086);
and AND3_2064 (N7697,  N7531,  N1731,  N3086);
or OR2_2065 (N7698,  N7624,  N7625);
not NOT1_2066 (N7699,  N7573);
not NOT1_2067 (N7700,  N7567);
not NOT1_2068 (N7701,  N7561);
not NOT1_2069 (N7702,  N7555);
and AND3_2070 (N7703,  N1156,  N7631,  N245);
not NOT1_2071 (N7704,  N7549);
not NOT1_2072 (N7705,  N7543);
not NOT1_2073 (N7706,  N7537);
not NOT1_2074 (N7707,  N7531);
not NOT1_2075 (N7708,  N7579);
nand NAND2_2076 (N7709,  N7579,  N6739);
not NOT1_2077 (N7710,  N7582);
nand NAND2_2078 (N7711,  N7582,  N6744);
nand NAND2_2079 (N7712,  N7657,  N7586);
nand NAND2_2080 (N7715,  N7658,  N7588);
not NOT1_2081 (N7718,  N7589);
nand NAND2_2082 (N7719,  N7589,  N6772);
not NOT1_2083 (N7720,  N7592);
nand NAND2_2084 (N7721,  N7592,  N6776);
not NOT1_2085 (N7722,  N7595);
nand NAND2_2086 (N7723,  N7595,  N5733);
nand NAND2_2087 (N7724,  N7665,  N7599);
or OR4_2088 (N7727,  N7666,  N7667,  N3617,  N2586);
or OR4_2089 (N7728,  N7668,  N7669,  N3618,  N2587);
or OR4_2090 (N7729,  N7670,  N7671,  N3619,  N2588);
or OR4_2091 (N7730,  N7672,  N7673,  N3620,  N2589);
or OR4_2092 (N7731,  N7674,  N7675,  N3628,  N2596);
or OR4_2093 (N7732,  N7676,  N7677,  N3629,  N2597);
or OR4_2094 (N7733,  N7678,  N7679,  N3630,  N2598);
or OR4_2095 (N7734,  N7680,  N7681,  N3631,  N2599);
or OR4_2096 (N7735,  N7682,  N7683,  N3638,  N2604);
or OR4_2097 (N7736,  N7684,  N7685,  N3642,  N2606);
or OR4_2098 (N7737,  N7686,  N7687,  N3643,  N2607);
or OR4_2099 (N7738,  N7688,  N7689,  N3644,  N2608);
or OR4_2100 (N7739,  N7690,  N7691,  N3645,  N2609);
or OR4_2101 (N7740,  N7692,  N7693,  N3651,  N2615);
or OR4_2102 (N7741,  N7694,  N7695,  N3652,  N2616);
or OR4_2103 (N7742,  N7696,  N7697,  N3653,  N2617);
nand NAND2_2104 (N7743,  N6271,  N7708);
nand NAND2_2105 (N7744,  N6283,  N7710);
nand NAND2_2106 (N7749,  N6341,  N7718);
nand NAND2_2107 (N7750,  N6347,  N7720);
nand NAND2_2108 (N7751,  N5214,  N7722);
and AND2_2109 (N7754,  N7727,  N2647);
and AND2_2110 (N7755,  N7728,  N2647);
and AND2_2111 (N7756,  N7729,  N2647);
and AND2_2112 (N7757,  N7730,  N2647);
and AND2_2113 (N7758,  N7731,  N2722);
and AND2_2114 (N7759,  N7732,  N2722);
and AND2_2115 (N7760,  N7733,  N2722);
and AND2_2116 (N7761,  N7734,  N2722);
nand NAND2_2117 (N7762,  N7743,  N7709);
nand NAND2_2118 (N7765,  N7744,  N7711);
not NOT1_2119 (N7768,  N7712);
nand NAND2_2120 (N7769,  N7712,  N6751);
not NOT1_2121 (N7770,  N7715);
nand NAND2_2122 (N7771,  N7715,  N6760);
nand NAND2_2123 (N7772,  N7749,  N7719);
nand NAND2_2124 (N7775,  N7750,  N7721);
nand NAND2_2125 (N7778,  N7751,  N7723);
not NOT1_2126 (N7781,  N7724);
nand NAND2_2127 (N7782,  N7724,  N5735);
nand NAND2_2128 (N7787,  N6295,  N7768);
nand NAND2_2129 (N7788,  N6313,  N7770);
nand NAND2_2130 (N7795,  N5220,  N7781);
not NOT1_2131 (N7796,  N7762);
nand NAND2_2132 (N7797,  N7762,  N6740);
not NOT1_2133 (N7798,  N7765);
nand NAND2_2134 (N7799,  N7765,  N6745);
nand NAND2_2135 (N7800,  N7787,  N7769);
nand NAND2_2136 (N7803,  N7788,  N7771);
not NOT1_2137 (N7806,  N7772);
nand NAND2_2138 (N7807,  N7772,  N6773);
not NOT1_2139 (N7808,  N7775);
nand NAND2_2140 (N7809,  N7775,  N6777);
not NOT1_2141 (N7810,  N7778);
nand NAND2_2142 (N7811,  N7778,  N6782);
nand NAND2_2143 (N7812,  N7795,  N7782);
nand NAND2_2144 (N7815,  N6274,  N7796);
nand NAND2_2145 (N7816,  N6286,  N7798);
nand NAND2_2146 (N7821,  N6344,  N7806);
nand NAND2_2147 (N7822,  N6350,  N7808);
nand NAND2_2148 (N7823,  N6353,  N7810);
nand NAND2_2149 (N7826,  N7815,  N7797);
nand NAND2_2150 (N7829,  N7816,  N7799);
not NOT1_2151 (N7832,  N7800);
nand NAND2_2152 (N7833,  N7800,  N6752);
not NOT1_2153 (N7834,  N7803);
nand NAND2_2154 (N7835,  N7803,  N6761);
nand NAND2_2155 (N7836,  N7821,  N7807);
nand NAND2_2156 (N7839,  N7822,  N7809);
nand NAND2_2157 (N7842,  N7823,  N7811);
not NOT1_2158 (N7845,  N7812);
nand NAND2_2159 (N7846,  N7812,  N6790);
nand NAND2_2160 (N7851,  N6298,  N7832);
nand NAND2_2161 (N7852,  N6316,  N7834);
nand NAND2_2162 (N7859,  N6364,  N7845);
not NOT1_2163 (N7860,  N7826);
nand NAND2_2164 (N7861,  N7826,  N6741);
not NOT1_2165 (N7862,  N7829);
nand NAND2_2166 (N7863,  N7829,  N6746);
nand NAND2_2167 (N7864,  N7851,  N7833);
nand NAND2_2168 (N7867,  N7852,  N7835);
not NOT1_2169 (N7870,  N7836);
nand NAND2_2170 (N7871,  N7836,  N5730);
not NOT1_2171 (N7872,  N7839);
nand NAND2_2172 (N7873,  N7839,  N5732);
not NOT1_2173 (N7874,  N7842);
nand NAND2_2174 (N7875,  N7842,  N6783);
nand NAND2_2175 (N7876,  N7859,  N7846);
nand NAND2_2176 (N7879,  N6277,  N7860);
nand NAND2_2177 (N7880,  N6289,  N7862);
nand NAND2_2178 (N7885,  N5199,  N7870);
nand NAND2_2179 (N7886,  N5208,  N7872);
nand NAND2_2180 (N7887,  N6356,  N7874);
nand NAND2_2181 (N7890,  N7879,  N7861);
nand NAND2_2182 (N7893,  N7880,  N7863);
not NOT1_2183 (N7896,  N7864);
nand NAND2_2184 (N7897,  N7864,  N6753);
not NOT1_2185 (N7898,  N7867);
nand NAND2_2186 (N7899,  N7867,  N6762);
nand NAND2_2187 (N7900,  N7885,  N7871);
nand NAND2_2188 (N7903,  N7886,  N7873);
nand NAND2_2189 (N7906,  N7887,  N7875);
not NOT1_2190 (N7909,  N7876);
nand NAND2_2191 (N7910,  N7876,  N6791);
nand NAND2_2192 (N7917,  N6301,  N7896);
nand NAND2_2193 (N7918,  N6319,  N7898);
nand NAND2_2194 (N7923,  N6367,  N7909);
not NOT1_2195 (N7924,  N7890);
nand NAND2_2196 (N7925,  N7890,  N6680);
not NOT1_2197 (N7926,  N7893);
nand NAND2_2198 (N7927,  N7893,  N6681);
not NOT1_2199 (N7928,  N7900);
nand NAND2_2200 (N7929,  N7900,  N5690);
not NOT1_2201 (N7930,  N7903);
nand NAND2_2202 (N7931,  N7903,  N5691);
nand NAND2_2203 (N7932,  N7917,  N7897);
nand NAND2_2204 (N7935,  N7918,  N7899);
not NOT1_2205 (N7938,  N7906);
nand NAND2_2206 (N7939,  N7906,  N6784);
nand NAND2_2207 (N7940,  N7923,  N7910);
nand NAND2_2208 (N7943,  N6280,  N7924);
nand NAND2_2209 (N7944,  N6292,  N7926);
nand NAND2_2210 (N7945,  N5202,  N7928);
nand NAND2_2211 (N7946,  N5211,  N7930);
nand NAND2_2212 (N7951,  N6359,  N7938);
nand NAND2_2213 (N7954,  N7943,  N7925);
nand NAND2_2214 (N7957,  N7944,  N7927);
nand NAND2_2215 (N7960,  N7945,  N7929);
nand NAND2_2216 (N7963,  N7946,  N7931);
not NOT1_2217 (N7966,  N7932);
nand NAND2_2218 (N7967,  N7932,  N6754);
not NOT1_2219 (N7968,  N7935);
nand NAND2_2220 (N7969,  N7935,  N6755);
nand NAND2_2221 (N7970,  N7951,  N7939);
not NOT1_2222 (N7973,  N7940);
nand NAND2_2223 (N7974,  N7940,  N6785);
nand NAND2_2224 (N7984,  N6304,  N7966);
nand NAND2_2225 (N7985,  N6322,  N7968);
nand NAND2_2226 (N7987,  N6370,  N7973);
and AND3_2227 (N7988,  N7957,  N6831,  N1157);
and AND3_2228 (N7989,  N7954,  N6415,  N1157);
and AND3_2229 (N7990,  N7957,  N7041,  N566);
and AND3_2230 (N7991,  N7954,  N7177,  N566);
not NOT1_2231 (N7992,  N7970);
nand NAND2_2232 (N7993,  N7970,  N6448);
and AND3_2233 (N7994,  N7963,  N6857,  N1219);
and AND3_2234 (N7995,  N7960,  N6441,  N1219);
and AND3_2235 (N7996,  N7963,  N7065,  N583);
and AND3_2236 (N7997,  N7960,  N7182,  N583);
nand NAND2_2237 (N7998,  N7984,  N7967);
nand NAND2_2238 (N8001,  N7985,  N7969);
nand NAND2_2239 (N8004,  N7987,  N7974);
nand NAND2_2240 (N8009,  N6051,  N7992);
or OR4_2241 (N8013,  N7988,  N7989,  N7990,  N7991);
or OR4_2242 (N8017,  N7994,  N7995,  N7996,  N7997);
not NOT1_2243 (N8020,  N7998);
nand NAND2_2244 (N8021,  N7998,  N6682);
not NOT1_2245 (N8022,  N8001);
nand NAND2_2246 (N8023,  N8001,  N6683);
nand NAND2_2247 (N8025,  N8009,  N7993);
not NOT1_2248 (N8026,  N8004);
nand NAND2_2249 (N8027,  N8004,  N6449);
nand NAND2_2250 (N8031,  N6307,  N8020);
nand NAND2_2251 (N8032,  N6310,  N8022);
not NOT1_2252 (N8033,  N8013);
nand NAND2_2253 (N8034,  N6054,  N8026);
and AND2_2254 (N8035,  N583,  N8025);
not NOT1_2255 (N8036,  N8017);
nand NAND2_2256 (N8037,  N8031,  N8021);
nand NAND2_2257 (N8038,  N8032,  N8023);
nand NAND2_2258 (N8039,  N8034,  N8027);
not NOT1_2259 (N8040,  N8038);
and AND2_2260 (N8041,  N566,  N8037);
not NOT1_2261 (N8042,  N8039);
and AND2_2262 (N8043,  N8040,  N1157);
and AND2_2263 (N8044,  N8042,  N1219);
or OR2_2264 (N8045,  N8043,  N8041);
or OR2_2265 (N8048,  N8044,  N8035);
nand NAND2_2266 (N8055,  N8045,  N8033);
not NOT1_2267 (N8056,  N8045);
nand NAND2_2268 (N8057,  N8048,  N8036);
not NOT1_2269 (N8058,  N8048);
nand NAND2_2270 (N8059,  N8013,  N8056);
nand NAND2_2271 (N8060,  N8017,  N8058);
nand NAND2_2272 (N8061,  N8055,  N8059);
nand NAND2_2273 (N8064,  N8057,  N8060);
and AND3_2274 (N8071,  N8064,  N1777,  N3130);
and AND3_2275 (N8072,  N8061,  N1761,  N3108);
not NOT1_2276 (N8073,  N8061);
not NOT1_2277 (N8074,  N8064);
or OR4_2278 (N8075,  N7526,  N8071,  N3659,  N2625);
or OR4_2279 (N8076,  N7636,  N8072,  N3661,  N2627);
and AND2_2280 (N8077,  N8073,  N1727);
and AND2_2281 (N8078,  N8074,  N1727);
or OR2_2282 (N8079,  N7530,  N8077);
or OR2_2283 (N8082,  N7479,  N8078);
and AND2_2284 (N8089,  N8079,  N3063);
and AND2_2285 (N8090,  N8082,  N3063);
and AND2_2286 (N8091,  N8079,  N3063);
and AND2_2287 (N8092,  N8082,  N3063);
or OR2_2288 (N8093,  N8089,  N3071);
or OR2_2289 (N8096,  N8090,  N3072);
or OR2_2290 (N8099,  N8091,  N3073);
or OR2_2291 (N8102,  N8092,  N3074);
and AND3_2292 (N8113,  N8102,  N2779,  N2790);
and AND3_2293 (N8114,  N8099,  N1327,  N2790);
and AND3_2294 (N8115,  N8102,  N2801,  N2812);
and AND3_2295 (N8116,  N8099,  N1351,  N2812);
and AND3_2296 (N8117,  N8096,  N2681,  N2692);
and AND3_2297 (N8118,  N8093,  N1185,  N2692);
and AND3_2298 (N8119,  N8096,  N2756,  N2767);
and AND3_2299 (N8120,  N8093,  N1247,  N2767);
or OR4_2300 (N8121,  N8117,  N8118,  N3662,  N2703);
or OR4_2301 (N8122,  N8119,  N8120,  N3663,  N2778);
or OR4_2302 (N8123,  N8113,  N8114,  N3650,  N2614);
or OR4_2303 (N8124,  N8115,  N8116,  N3658,  N2622);
and AND2_2304 (N8125,  N8121,  N2675);
and AND2_2305 (N8126,  N8122,  N2750);
not NOT1_2306 (N8127,  N8125);
not NOT1_2307 (N8128,  N8126);

endmodule
