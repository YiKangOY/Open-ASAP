module sk16 (in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, );
input in0;
input in1;
input in2;
input in3;
input in4;
input in5;
input in6;
input in7;
input in8;
input in9;
input in10;
input in11;
input in12;
input in13;
input in14;
input in15;
input in16;
input in17;
input in18;
input in19;
input in20;
input in21;
input in22;
input in23;
input in24;
input in25;
input in26;
input in27;
input in28;
input in29;
input in30;
input in31;
output out0;
output out1;
output out2;
output out3;
output out4;
output out5;
output out6;
output out7;
output out8;
output out9;
output out10;
output out11;
output out12;
output out13;
output out14;
output out15;
output out16;
wire var0;
wire var1;
wire var2;
wire var3;
wire var4;
wire var5;
wire var6;
wire var7;
wire var8;
wire var9;
wire var10;
wire var11;
wire var12;
wire var13;
wire var14;
wire var15;
wire var16;
wire var17;
wire var18;
wire var19;
wire var20;
wire var21;
wire var22;
wire var23;
wire var24;
wire var25;
wire var26;
wire var27;
wire var28;
wire var29;
wire var30;
wire var31;
wire var32;
wire var33;
wire var34;
wire var35;
wire var36;
wire var37;
wire var38;
wire var39;
wire var40;
wire var41;
wire var42;
wire var43;
wire var44;
wire var45;
wire var46;
wire var47;
wire var48;
wire var49;
wire var50;
wire var51;
wire var52;
wire var53;
wire var54;
wire var55;
wire var56;
wire var57;
wire var58;
wire var59;
wire var60;
wire var61;
wire var62;
wire var63;
wire var64;
wire var65;
wire var66;
wire var67;
wire var68;
wire var69;
wire var70;
wire var71;
wire var72;
wire var73;
wire var74;
wire var75;
wire var76;
wire var77;
wire var78;
wire var79;
wire var80;
wire var81;
wire var82;
wire var83;
wire var84;
wire var85;
wire var86;
wire var87;
wire var88;
wire var89;
wire var90;
wire var91;
wire var92;
wire var93;
wire var94;
wire var95;
wire var96;
wire var97;
wire var98;
wire var99;
wire var100;
wire var101;
wire var102;
wire var103;
wire var104;
wire var105;
wire var106;
wire var107;
wire var108;
wire var109;
wire var110;
wire var111;
wire var112;
wire var113;
wire var114;
wire var115;
wire var116;
wire var117;
wire var118;
wire var119;
wire var120;
wire var121;
wire var122;
wire var123;
wire var124;
wire var125;
wire var126;
wire var127;
assign var0 = in31 & in15;
assign var1 = in30 & in14;
assign var2 = in29 & in13;
assign var3 = in28 & in12;
assign var4 = in27 & in11;
assign var5 = in26 & in10;
assign var6 = in25 & in9;
assign var7 = in24 & in8;
assign var8 = in23 & in7;
assign var9 = in22 & in6;
assign var10 = in21 & in5;
assign var11 = in20 & in4;
assign var12 = in19 & in3;
assign var13 = in18 & in2;
assign var14 = in17 & in1;
assign var15 = in16 & in0;
assign var16 = in31 ^ in15;
assign var17 = in30 ^ in14;
assign var18 = in29 ^ in13;
assign var19 = in28 ^ in12;
assign var20 = in27 ^ in11;
assign var21 = in26 ^ in10;
assign var22 = in25 ^ in9;
assign var23 = in24 ^ in8;
assign var24 = in23 ^ in7;
assign var25 = in22 ^ in6;
assign var26 = in21 ^ in5;
assign var27 = in20 ^ in4;
assign var28 = in19 ^ in3;
assign var29 = in18 ^ in2;
assign var30 = in17 ^ in1;
assign var31 = in16 ^ in0;
assign var32 = var31 & var14;
assign var33 = var15 | var32;
assign var34 = var31 & var30;
assign var35 = var29 & var12;
assign var36 = var13 | var35;
assign var37 = var29 & var28;
assign var38 = var27 & var10;
assign var39 = var11 | var38;
assign var40 = var27 & var26;
assign var41 = var25 & var8;
assign var42 = var9 | var41;
assign var43 = var25 & var24;
assign var44 = var23 & var6;
assign var45 = var7 | var44;
assign var46 = var23 & var22;
assign var47 = var21 & var4;
assign var48 = var5 | var47;
assign var49 = var21 & var20;
assign var50 = var19 & var2;
assign var51 = var3 | var50;
assign var52 = var19 & var18;
assign var53 = var17 & var0;
assign var54 = var1 | var53;
assign var55 = var34 & var36;
assign var56 = var33 | var55;
assign var57 = var34 & var37;
assign var58 = var30 & var36;
assign var59 = var14 | var58;
assign var60 = var30 & var37;
assign var61 = var40 & var42;
assign var62 = var39 | var61;
assign var63 = var40 & var43;
assign var64 = var26 & var42;
assign var65 = var10 | var64;
assign var66 = var26 & var43;
assign var67 = var46 & var48;
assign var68 = var45 | var67;
assign var69 = var46 & var49;
assign var70 = var22 & var48;
assign var71 = var6 | var70;
assign var72 = var22 & var49;
assign var73 = var52 & var54;
assign var74 = var51 | var73;
assign var75 = var18 & var54;
assign var76 = var2 | var75;
assign var77 = var57 & var62;
assign var78 = var56 | var77;
assign var79 = var57 & var63;
assign var80 = var60 & var62;
assign var81 = var59 | var80;
assign var82 = var60 & var63;
assign var83 = var37 & var62;
assign var84 = var36 | var83;
assign var85 = var37 & var63;
assign var86 = var28 & var62;
assign var87 = var12 | var86;
assign var88 = var28 & var63;
assign var89 = var69 & var74;
assign var90 = var68 | var89;
assign var91 = var72 & var74;
assign var92 = var71 | var91;
assign var93 = var49 & var74;
assign var94 = var48 | var93;
assign var95 = var20 & var74;
assign var96 = var4 | var95;
assign var97 = var79 & var90;
assign var98 = var78 | var97;
assign var99 = var82 & var90;
assign var100 = var81 | var99;
assign var101 = var85 & var90;
assign var102 = var84 | var101;
assign var103 = var88 & var90;
assign var104 = var87 | var103;
assign var105 = var63 & var90;
assign var106 = var62 | var105;
assign var107 = var66 & var90;
assign var108 = var65 | var107;
assign var109 = var43 & var90;
assign var110 = var42 | var109;
assign var111 = var24 & var90;
assign var112 = var8 | var111;
assign var113 = var17 ^ var0;
assign var114 = var18 ^ var54;
assign var115 = var19 ^ var76;
assign var116 = var20 ^ var74;
assign var117 = var21 ^ var96;
assign var118 = var22 ^ var94;
assign var119 = var23 ^ var92;
assign var120 = var24 ^ var90;
assign var121 = var25 ^ var112;
assign var122 = var26 ^ var110;
assign var123 = var27 ^ var108;
assign var124 = var28 ^ var106;
assign var125 = var29 ^ var104;
assign var126 = var30 ^ var102;
assign var127 = var31 ^ var100;
assign out0 = var98;
assign out1 = var127;
assign out2 = var126;
assign out3 = var125;
assign out4 = var124;
assign out5 = var123;
assign out6 = var122;
assign out7 = var121;
assign out8 = var120;
assign out9 = var119;
assign out10 = var118;
assign out11 = var117;
assign out12 = var116;
assign out13 = var115;
assign out14 = var114;
assign out15 = var113;
assign out16 = var16;
endmodule 
