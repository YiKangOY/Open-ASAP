module hc64 (in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, in100, in101, in102, in103, in104, in105, in106, in107, in108, in109, in110, in111, in112, in113, in114, in115, in116, in117, in118, in119, in120, in121, in122, in123, in124, in125, in126, in127, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, out30, out31, out32, out33, out34, out35, out36, out37, out38, out39, out40, out41, out42, out43, out44, out45, out46, out47, out48, out49, out50, out51, out52, out53, out54, out55, out56, out57, out58, out59, out60, out61, out62, out63, out64, );
input in0;
input in1;
input in2;
input in3;
input in4;
input in5;
input in6;
input in7;
input in8;
input in9;
input in10;
input in11;
input in12;
input in13;
input in14;
input in15;
input in16;
input in17;
input in18;
input in19;
input in20;
input in21;
input in22;
input in23;
input in24;
input in25;
input in26;
input in27;
input in28;
input in29;
input in30;
input in31;
input in32;
input in33;
input in34;
input in35;
input in36;
input in37;
input in38;
input in39;
input in40;
input in41;
input in42;
input in43;
input in44;
input in45;
input in46;
input in47;
input in48;
input in49;
input in50;
input in51;
input in52;
input in53;
input in54;
input in55;
input in56;
input in57;
input in58;
input in59;
input in60;
input in61;
input in62;
input in63;
input in64;
input in65;
input in66;
input in67;
input in68;
input in69;
input in70;
input in71;
input in72;
input in73;
input in74;
input in75;
input in76;
input in77;
input in78;
input in79;
input in80;
input in81;
input in82;
input in83;
input in84;
input in85;
input in86;
input in87;
input in88;
input in89;
input in90;
input in91;
input in92;
input in93;
input in94;
input in95;
input in96;
input in97;
input in98;
input in99;
input in100;
input in101;
input in102;
input in103;
input in104;
input in105;
input in106;
input in107;
input in108;
input in109;
input in110;
input in111;
input in112;
input in113;
input in114;
input in115;
input in116;
input in117;
input in118;
input in119;
input in120;
input in121;
input in122;
input in123;
input in124;
input in125;
input in126;
input in127;
output out0;
output out1;
output out2;
output out3;
output out4;
output out5;
output out6;
output out7;
output out8;
output out9;
output out10;
output out11;
output out12;
output out13;
output out14;
output out15;
output out16;
output out17;
output out18;
output out19;
output out20;
output out21;
output out22;
output out23;
output out24;
output out25;
output out26;
output out27;
output out28;
output out29;
output out30;
output out31;
output out32;
output out33;
output out34;
output out35;
output out36;
output out37;
output out38;
output out39;
output out40;
output out41;
output out42;
output out43;
output out44;
output out45;
output out46;
output out47;
output out48;
output out49;
output out50;
output out51;
output out52;
output out53;
output out54;
output out55;
output out56;
output out57;
output out58;
output out59;
output out60;
output out61;
output out62;
output out63;
output out64;
wire var0;
wire var1;
wire var2;
wire var3;
wire var4;
wire var5;
wire var6;
wire var7;
wire var8;
wire var9;
wire var10;
wire var11;
wire var12;
wire var13;
wire var14;
wire var15;
wire var16;
wire var17;
wire var18;
wire var19;
wire var20;
wire var21;
wire var22;
wire var23;
wire var24;
wire var25;
wire var26;
wire var27;
wire var28;
wire var29;
wire var30;
wire var31;
wire var32;
wire var33;
wire var34;
wire var35;
wire var36;
wire var37;
wire var38;
wire var39;
wire var40;
wire var41;
wire var42;
wire var43;
wire var44;
wire var45;
wire var46;
wire var47;
wire var48;
wire var49;
wire var50;
wire var51;
wire var52;
wire var53;
wire var54;
wire var55;
wire var56;
wire var57;
wire var58;
wire var59;
wire var60;
wire var61;
wire var62;
wire var63;
wire var64;
wire var65;
wire var66;
wire var67;
wire var68;
wire var69;
wire var70;
wire var71;
wire var72;
wire var73;
wire var74;
wire var75;
wire var76;
wire var77;
wire var78;
wire var79;
wire var80;
wire var81;
wire var82;
wire var83;
wire var84;
wire var85;
wire var86;
wire var87;
wire var88;
wire var89;
wire var90;
wire var91;
wire var92;
wire var93;
wire var94;
wire var95;
wire var96;
wire var97;
wire var98;
wire var99;
wire var100;
wire var101;
wire var102;
wire var103;
wire var104;
wire var105;
wire var106;
wire var107;
wire var108;
wire var109;
wire var110;
wire var111;
wire var112;
wire var113;
wire var114;
wire var115;
wire var116;
wire var117;
wire var118;
wire var119;
wire var120;
wire var121;
wire var122;
wire var123;
wire var124;
wire var125;
wire var126;
wire var127;
wire var128;
wire var129;
wire var130;
wire var131;
wire var132;
wire var133;
wire var134;
wire var135;
wire var136;
wire var137;
wire var138;
wire var139;
wire var140;
wire var141;
wire var142;
wire var143;
wire var144;
wire var145;
wire var146;
wire var147;
wire var148;
wire var149;
wire var150;
wire var151;
wire var152;
wire var153;
wire var154;
wire var155;
wire var156;
wire var157;
wire var158;
wire var159;
wire var160;
wire var161;
wire var162;
wire var163;
wire var164;
wire var165;
wire var166;
wire var167;
wire var168;
wire var169;
wire var170;
wire var171;
wire var172;
wire var173;
wire var174;
wire var175;
wire var176;
wire var177;
wire var178;
wire var179;
wire var180;
wire var181;
wire var182;
wire var183;
wire var184;
wire var185;
wire var186;
wire var187;
wire var188;
wire var189;
wire var190;
wire var191;
wire var192;
wire var193;
wire var194;
wire var195;
wire var196;
wire var197;
wire var198;
wire var199;
wire var200;
wire var201;
wire var202;
wire var203;
wire var204;
wire var205;
wire var206;
wire var207;
wire var208;
wire var209;
wire var210;
wire var211;
wire var212;
wire var213;
wire var214;
wire var215;
wire var216;
wire var217;
wire var218;
wire var219;
wire var220;
wire var221;
wire var222;
wire var223;
wire var224;
wire var225;
wire var226;
wire var227;
wire var228;
wire var229;
wire var230;
wire var231;
wire var232;
wire var233;
wire var234;
wire var235;
wire var236;
wire var237;
wire var238;
wire var239;
wire var240;
wire var241;
wire var242;
wire var243;
wire var244;
wire var245;
wire var246;
wire var247;
wire var248;
wire var249;
wire var250;
wire var251;
wire var252;
wire var253;
wire var254;
wire var255;
wire var256;
wire var257;
wire var258;
wire var259;
wire var260;
wire var261;
wire var262;
wire var263;
wire var264;
wire var265;
wire var266;
wire var267;
wire var268;
wire var269;
wire var270;
wire var271;
wire var272;
wire var273;
wire var274;
wire var275;
wire var276;
wire var277;
wire var278;
wire var279;
wire var280;
wire var281;
wire var282;
wire var283;
wire var284;
wire var285;
wire var286;
wire var287;
wire var288;
wire var289;
wire var290;
wire var291;
wire var292;
wire var293;
wire var294;
wire var295;
wire var296;
wire var297;
wire var298;
wire var299;
wire var300;
wire var301;
wire var302;
wire var303;
wire var304;
wire var305;
wire var306;
wire var307;
wire var308;
wire var309;
wire var310;
wire var311;
wire var312;
wire var313;
wire var314;
wire var315;
wire var316;
wire var317;
wire var318;
wire var319;
wire var320;
wire var321;
wire var322;
wire var323;
wire var324;
wire var325;
wire var326;
wire var327;
wire var328;
wire var329;
wire var330;
wire var331;
wire var332;
wire var333;
wire var334;
wire var335;
wire var336;
wire var337;
wire var338;
wire var339;
wire var340;
wire var341;
wire var342;
wire var343;
wire var344;
wire var345;
wire var346;
wire var347;
wire var348;
wire var349;
wire var350;
wire var351;
wire var352;
wire var353;
wire var354;
wire var355;
wire var356;
wire var357;
wire var358;
wire var359;
wire var360;
wire var361;
wire var362;
wire var363;
wire var364;
wire var365;
wire var366;
wire var367;
wire var368;
wire var369;
wire var370;
wire var371;
wire var372;
wire var373;
wire var374;
wire var375;
wire var376;
wire var377;
wire var378;
wire var379;
wire var380;
wire var381;
wire var382;
wire var383;
wire var384;
wire var385;
wire var386;
wire var387;
wire var388;
wire var389;
wire var390;
wire var391;
wire var392;
wire var393;
wire var394;
wire var395;
wire var396;
wire var397;
wire var398;
wire var399;
wire var400;
wire var401;
wire var402;
wire var403;
wire var404;
wire var405;
wire var406;
wire var407;
wire var408;
wire var409;
wire var410;
wire var411;
wire var412;
wire var413;
wire var414;
wire var415;
wire var416;
wire var417;
wire var418;
wire var419;
wire var420;
wire var421;
wire var422;
wire var423;
wire var424;
wire var425;
wire var426;
wire var427;
wire var428;
wire var429;
wire var430;
wire var431;
wire var432;
wire var433;
wire var434;
wire var435;
wire var436;
wire var437;
wire var438;
wire var439;
wire var440;
wire var441;
wire var442;
wire var443;
wire var444;
wire var445;
wire var446;
wire var447;
wire var448;
wire var449;
wire var450;
wire var451;
wire var452;
wire var453;
wire var454;
wire var455;
wire var456;
wire var457;
wire var458;
wire var459;
wire var460;
wire var461;
wire var462;
wire var463;
wire var464;
wire var465;
wire var466;
wire var467;
wire var468;
wire var469;
wire var470;
wire var471;
wire var472;
wire var473;
wire var474;
wire var475;
wire var476;
wire var477;
wire var478;
wire var479;
wire var480;
wire var481;
wire var482;
wire var483;
wire var484;
wire var485;
wire var486;
wire var487;
wire var488;
wire var489;
wire var490;
wire var491;
wire var492;
wire var493;
wire var494;
wire var495;
wire var496;
wire var497;
wire var498;
wire var499;
wire var500;
wire var501;
wire var502;
wire var503;
wire var504;
wire var505;
wire var506;
wire var507;
wire var508;
wire var509;
wire var510;
wire var511;
wire var512;
wire var513;
wire var514;
wire var515;
wire var516;
wire var517;
wire var518;
wire var519;
wire var520;
wire var521;
wire var522;
wire var523;
wire var524;
wire var525;
wire var526;
wire var527;
wire var528;
wire var529;
wire var530;
wire var531;
wire var532;
wire var533;
wire var534;
wire var535;
wire var536;
wire var537;
wire var538;
wire var539;
wire var540;
wire var541;
wire var542;
wire var543;
wire var544;
wire var545;
wire var546;
wire var547;
wire var548;
wire var549;
wire var550;
wire var551;
wire var552;
wire var553;
wire var554;
wire var555;
wire var556;
wire var557;
wire var558;
wire var559;
wire var560;
wire var561;
wire var562;
wire var563;
wire var564;
wire var565;
wire var566;
wire var567;
wire var568;
wire var569;
wire var570;
wire var571;
wire var572;
wire var573;
wire var574;
wire var575;
wire var576;
wire var577;
wire var578;
wire var579;
wire var580;
wire var581;
wire var582;
wire var583;
wire var584;
wire var585;
wire var586;
wire var587;
wire var588;
wire var589;
wire var590;
wire var591;
wire var592;
wire var593;
wire var594;
wire var595;
wire var596;
wire var597;
wire var598;
wire var599;
wire var600;
wire var601;
wire var602;
wire var603;
wire var604;
wire var605;
wire var606;
wire var607;
wire var608;
wire var609;
wire var610;
wire var611;
wire var612;
wire var613;
wire var614;
wire var615;
wire var616;
wire var617;
wire var618;
wire var619;
wire var620;
wire var621;
wire var622;
wire var623;
wire var624;
wire var625;
wire var626;
wire var627;
wire var628;
wire var629;
wire var630;
wire var631;
wire var632;
wire var633;
wire var634;
wire var635;
wire var636;
wire var637;
wire var638;
wire var639;
wire var640;
wire var641;
wire var642;
wire var643;
wire var644;
wire var645;
wire var646;
wire var647;
wire var648;
wire var649;
wire var650;
wire var651;
wire var652;
wire var653;
wire var654;
wire var655;
wire var656;
wire var657;
wire var658;
wire var659;
wire var660;
wire var661;
wire var662;
wire var663;
wire var664;
wire var665;
wire var666;
wire var667;
wire var668;
wire var669;
wire var670;
wire var671;
wire var672;
wire var673;
wire var674;
wire var675;
wire var676;
wire var677;
wire var678;
wire var679;
wire var680;
wire var681;
wire var682;
wire var683;
wire var684;
wire var685;
wire var686;
wire var687;
wire var688;
wire var689;
wire var690;
wire var691;
wire var692;
wire var693;
wire var694;
wire var695;
wire var696;
wire var697;
wire var698;
wire var699;
wire var700;
wire var701;
wire var702;
wire var703;
wire var704;
wire var705;
wire var706;
wire var707;
wire var708;
wire var709;
wire var710;
wire var711;
wire var712;
wire var713;
wire var714;
wire var715;
wire var716;
wire var717;
wire var718;
wire var719;
wire var720;
wire var721;
wire var722;
wire var723;
wire var724;
wire var725;
wire var726;
wire var727;
wire var728;
wire var729;
wire var730;
wire var731;
wire var732;
wire var733;
wire var734;
assign var0 = in127 & in63;
assign var1 = in126 & in62;
assign var2 = in125 & in61;
assign var3 = in124 & in60;
assign var4 = in123 & in59;
assign var5 = in122 & in58;
assign var6 = in121 & in57;
assign var7 = in120 & in56;
assign var8 = in119 & in55;
assign var9 = in118 & in54;
assign var10 = in117 & in53;
assign var11 = in116 & in52;
assign var12 = in115 & in51;
assign var13 = in114 & in50;
assign var14 = in113 & in49;
assign var15 = in112 & in48;
assign var16 = in111 & in47;
assign var17 = in110 & in46;
assign var18 = in109 & in45;
assign var19 = in108 & in44;
assign var20 = in107 & in43;
assign var21 = in106 & in42;
assign var22 = in105 & in41;
assign var23 = in104 & in40;
assign var24 = in103 & in39;
assign var25 = in102 & in38;
assign var26 = in101 & in37;
assign var27 = in100 & in36;
assign var28 = in99 & in35;
assign var29 = in98 & in34;
assign var30 = in97 & in33;
assign var31 = in96 & in32;
assign var32 = in95 & in31;
assign var33 = in94 & in30;
assign var34 = in93 & in29;
assign var35 = in92 & in28;
assign var36 = in91 & in27;
assign var37 = in90 & in26;
assign var38 = in89 & in25;
assign var39 = in88 & in24;
assign var40 = in87 & in23;
assign var41 = in86 & in22;
assign var42 = in85 & in21;
assign var43 = in84 & in20;
assign var44 = in83 & in19;
assign var45 = in82 & in18;
assign var46 = in81 & in17;
assign var47 = in80 & in16;
assign var48 = in79 & in15;
assign var49 = in78 & in14;
assign var50 = in77 & in13;
assign var51 = in76 & in12;
assign var52 = in75 & in11;
assign var53 = in74 & in10;
assign var54 = in73 & in9;
assign var55 = in72 & in8;
assign var56 = in71 & in7;
assign var57 = in70 & in6;
assign var58 = in69 & in5;
assign var59 = in68 & in4;
assign var60 = in67 & in3;
assign var61 = in66 & in2;
assign var62 = in65 & in1;
assign var63 = in64 & in0;
assign var64 = in127 ^ in63;
assign var65 = in126 ^ in62;
assign var66 = in125 ^ in61;
assign var67 = in124 ^ in60;
assign var68 = in123 ^ in59;
assign var69 = in122 ^ in58;
assign var70 = in121 ^ in57;
assign var71 = in120 ^ in56;
assign var72 = in119 ^ in55;
assign var73 = in118 ^ in54;
assign var74 = in117 ^ in53;
assign var75 = in116 ^ in52;
assign var76 = in115 ^ in51;
assign var77 = in114 ^ in50;
assign var78 = in113 ^ in49;
assign var79 = in112 ^ in48;
assign var80 = in111 ^ in47;
assign var81 = in110 ^ in46;
assign var82 = in109 ^ in45;
assign var83 = in108 ^ in44;
assign var84 = in107 ^ in43;
assign var85 = in106 ^ in42;
assign var86 = in105 ^ in41;
assign var87 = in104 ^ in40;
assign var88 = in103 ^ in39;
assign var89 = in102 ^ in38;
assign var90 = in101 ^ in37;
assign var91 = in100 ^ in36;
assign var92 = in99 ^ in35;
assign var93 = in98 ^ in34;
assign var94 = in97 ^ in33;
assign var95 = in96 ^ in32;
assign var96 = in95 ^ in31;
assign var97 = in94 ^ in30;
assign var98 = in93 ^ in29;
assign var99 = in92 ^ in28;
assign var100 = in91 ^ in27;
assign var101 = in90 ^ in26;
assign var102 = in89 ^ in25;
assign var103 = in88 ^ in24;
assign var104 = in87 ^ in23;
assign var105 = in86 ^ in22;
assign var106 = in85 ^ in21;
assign var107 = in84 ^ in20;
assign var108 = in83 ^ in19;
assign var109 = in82 ^ in18;
assign var110 = in81 ^ in17;
assign var111 = in80 ^ in16;
assign var112 = in79 ^ in15;
assign var113 = in78 ^ in14;
assign var114 = in77 ^ in13;
assign var115 = in76 ^ in12;
assign var116 = in75 ^ in11;
assign var117 = in74 ^ in10;
assign var118 = in73 ^ in9;
assign var119 = in72 ^ in8;
assign var120 = in71 ^ in7;
assign var121 = in70 ^ in6;
assign var122 = in69 ^ in5;
assign var123 = in68 ^ in4;
assign var124 = in67 ^ in3;
assign var125 = in66 ^ in2;
assign var126 = in65 ^ in1;
assign var127 = in64 ^ in0;
assign var128 = var127 & var62;
assign var129 = var63 | var128;
assign var130 = var127 & var126;
assign var131 = var125 & var60;
assign var132 = var61 | var131;
assign var133 = var125 & var124;
assign var134 = var123 & var58;
assign var135 = var59 | var134;
assign var136 = var123 & var122;
assign var137 = var121 & var56;
assign var138 = var57 | var137;
assign var139 = var121 & var120;
assign var140 = var119 & var54;
assign var141 = var55 | var140;
assign var142 = var119 & var118;
assign var143 = var117 & var52;
assign var144 = var53 | var143;
assign var145 = var117 & var116;
assign var146 = var115 & var50;
assign var147 = var51 | var146;
assign var148 = var115 & var114;
assign var149 = var113 & var48;
assign var150 = var49 | var149;
assign var151 = var113 & var112;
assign var152 = var111 & var46;
assign var153 = var47 | var152;
assign var154 = var111 & var110;
assign var155 = var109 & var44;
assign var156 = var45 | var155;
assign var157 = var109 & var108;
assign var158 = var107 & var42;
assign var159 = var43 | var158;
assign var160 = var107 & var106;
assign var161 = var105 & var40;
assign var162 = var41 | var161;
assign var163 = var105 & var104;
assign var164 = var103 & var38;
assign var165 = var39 | var164;
assign var166 = var103 & var102;
assign var167 = var101 & var36;
assign var168 = var37 | var167;
assign var169 = var101 & var100;
assign var170 = var99 & var34;
assign var171 = var35 | var170;
assign var172 = var99 & var98;
assign var173 = var97 & var32;
assign var174 = var33 | var173;
assign var175 = var97 & var96;
assign var176 = var95 & var30;
assign var177 = var31 | var176;
assign var178 = var95 & var94;
assign var179 = var93 & var28;
assign var180 = var29 | var179;
assign var181 = var93 & var92;
assign var182 = var91 & var26;
assign var183 = var27 | var182;
assign var184 = var91 & var90;
assign var185 = var89 & var24;
assign var186 = var25 | var185;
assign var187 = var89 & var88;
assign var188 = var87 & var22;
assign var189 = var23 | var188;
assign var190 = var87 & var86;
assign var191 = var85 & var20;
assign var192 = var21 | var191;
assign var193 = var85 & var84;
assign var194 = var83 & var18;
assign var195 = var19 | var194;
assign var196 = var83 & var82;
assign var197 = var81 & var16;
assign var198 = var17 | var197;
assign var199 = var81 & var80;
assign var200 = var79 & var14;
assign var201 = var15 | var200;
assign var202 = var79 & var78;
assign var203 = var77 & var12;
assign var204 = var13 | var203;
assign var205 = var77 & var76;
assign var206 = var75 & var10;
assign var207 = var11 | var206;
assign var208 = var75 & var74;
assign var209 = var73 & var8;
assign var210 = var9 | var209;
assign var211 = var73 & var72;
assign var212 = var71 & var6;
assign var213 = var7 | var212;
assign var214 = var71 & var70;
assign var215 = var69 & var4;
assign var216 = var5 | var215;
assign var217 = var69 & var68;
assign var218 = var67 & var2;
assign var219 = var3 | var218;
assign var220 = var67 & var66;
assign var221 = var65 & var0;
assign var222 = var1 | var221;
assign var223 = var130 & var132;
assign var224 = var129 | var223;
assign var225 = var130 & var133;
assign var226 = var133 & var135;
assign var227 = var132 | var226;
assign var228 = var133 & var136;
assign var229 = var136 & var138;
assign var230 = var135 | var229;
assign var231 = var136 & var139;
assign var232 = var139 & var141;
assign var233 = var138 | var232;
assign var234 = var139 & var142;
assign var235 = var142 & var144;
assign var236 = var141 | var235;
assign var237 = var142 & var145;
assign var238 = var145 & var147;
assign var239 = var144 | var238;
assign var240 = var145 & var148;
assign var241 = var148 & var150;
assign var242 = var147 | var241;
assign var243 = var148 & var151;
assign var244 = var151 & var153;
assign var245 = var150 | var244;
assign var246 = var151 & var154;
assign var247 = var154 & var156;
assign var248 = var153 | var247;
assign var249 = var154 & var157;
assign var250 = var157 & var159;
assign var251 = var156 | var250;
assign var252 = var157 & var160;
assign var253 = var160 & var162;
assign var254 = var159 | var253;
assign var255 = var160 & var163;
assign var256 = var163 & var165;
assign var257 = var162 | var256;
assign var258 = var163 & var166;
assign var259 = var166 & var168;
assign var260 = var165 | var259;
assign var261 = var166 & var169;
assign var262 = var169 & var171;
assign var263 = var168 | var262;
assign var264 = var169 & var172;
assign var265 = var172 & var174;
assign var266 = var171 | var265;
assign var267 = var172 & var175;
assign var268 = var175 & var177;
assign var269 = var174 | var268;
assign var270 = var175 & var178;
assign var271 = var178 & var180;
assign var272 = var177 | var271;
assign var273 = var178 & var181;
assign var274 = var181 & var183;
assign var275 = var180 | var274;
assign var276 = var181 & var184;
assign var277 = var184 & var186;
assign var278 = var183 | var277;
assign var279 = var184 & var187;
assign var280 = var187 & var189;
assign var281 = var186 | var280;
assign var282 = var187 & var190;
assign var283 = var190 & var192;
assign var284 = var189 | var283;
assign var285 = var190 & var193;
assign var286 = var193 & var195;
assign var287 = var192 | var286;
assign var288 = var193 & var196;
assign var289 = var196 & var198;
assign var290 = var195 | var289;
assign var291 = var196 & var199;
assign var292 = var199 & var201;
assign var293 = var198 | var292;
assign var294 = var199 & var202;
assign var295 = var202 & var204;
assign var296 = var201 | var295;
assign var297 = var202 & var205;
assign var298 = var205 & var207;
assign var299 = var204 | var298;
assign var300 = var205 & var208;
assign var301 = var208 & var210;
assign var302 = var207 | var301;
assign var303 = var208 & var211;
assign var304 = var211 & var213;
assign var305 = var210 | var304;
assign var306 = var211 & var214;
assign var307 = var214 & var216;
assign var308 = var213 | var307;
assign var309 = var214 & var217;
assign var310 = var217 & var219;
assign var311 = var216 | var310;
assign var312 = var217 & var220;
assign var313 = var220 & var222;
assign var314 = var219 | var313;
assign var315 = var225 & var230;
assign var316 = var224 | var315;
assign var317 = var225 & var231;
assign var318 = var228 & var233;
assign var319 = var227 | var318;
assign var320 = var228 & var234;
assign var321 = var231 & var236;
assign var322 = var230 | var321;
assign var323 = var231 & var237;
assign var324 = var234 & var239;
assign var325 = var233 | var324;
assign var326 = var234 & var240;
assign var327 = var237 & var242;
assign var328 = var236 | var327;
assign var329 = var237 & var243;
assign var330 = var240 & var245;
assign var331 = var239 | var330;
assign var332 = var240 & var246;
assign var333 = var243 & var248;
assign var334 = var242 | var333;
assign var335 = var243 & var249;
assign var336 = var246 & var251;
assign var337 = var245 | var336;
assign var338 = var246 & var252;
assign var339 = var249 & var254;
assign var340 = var248 | var339;
assign var341 = var249 & var255;
assign var342 = var252 & var257;
assign var343 = var251 | var342;
assign var344 = var252 & var258;
assign var345 = var255 & var260;
assign var346 = var254 | var345;
assign var347 = var255 & var261;
assign var348 = var258 & var263;
assign var349 = var257 | var348;
assign var350 = var258 & var264;
assign var351 = var261 & var266;
assign var352 = var260 | var351;
assign var353 = var261 & var267;
assign var354 = var264 & var269;
assign var355 = var263 | var354;
assign var356 = var264 & var270;
assign var357 = var267 & var272;
assign var358 = var266 | var357;
assign var359 = var267 & var273;
assign var360 = var270 & var275;
assign var361 = var269 | var360;
assign var362 = var270 & var276;
assign var363 = var273 & var278;
assign var364 = var272 | var363;
assign var365 = var273 & var279;
assign var366 = var276 & var281;
assign var367 = var275 | var366;
assign var368 = var276 & var282;
assign var369 = var279 & var284;
assign var370 = var278 | var369;
assign var371 = var279 & var285;
assign var372 = var282 & var287;
assign var373 = var281 | var372;
assign var374 = var282 & var288;
assign var375 = var285 & var290;
assign var376 = var284 | var375;
assign var377 = var285 & var291;
assign var378 = var288 & var293;
assign var379 = var287 | var378;
assign var380 = var288 & var294;
assign var381 = var291 & var296;
assign var382 = var290 | var381;
assign var383 = var291 & var297;
assign var384 = var294 & var299;
assign var385 = var293 | var384;
assign var386 = var294 & var300;
assign var387 = var297 & var302;
assign var388 = var296 | var387;
assign var389 = var297 & var303;
assign var390 = var300 & var305;
assign var391 = var299 | var390;
assign var392 = var300 & var306;
assign var393 = var303 & var308;
assign var394 = var302 | var393;
assign var395 = var303 & var309;
assign var396 = var306 & var311;
assign var397 = var305 | var396;
assign var398 = var306 & var312;
assign var399 = var309 & var314;
assign var400 = var308 | var399;
assign var401 = var312 & var222;
assign var402 = var311 | var401;
assign var403 = var317 & var328;
assign var404 = var316 | var403;
assign var405 = var317 & var329;
assign var406 = var320 & var331;
assign var407 = var319 | var406;
assign var408 = var320 & var332;
assign var409 = var323 & var334;
assign var410 = var322 | var409;
assign var411 = var323 & var335;
assign var412 = var326 & var337;
assign var413 = var325 | var412;
assign var414 = var326 & var338;
assign var415 = var329 & var340;
assign var416 = var328 | var415;
assign var417 = var329 & var341;
assign var418 = var332 & var343;
assign var419 = var331 | var418;
assign var420 = var332 & var344;
assign var421 = var335 & var346;
assign var422 = var334 | var421;
assign var423 = var335 & var347;
assign var424 = var338 & var349;
assign var425 = var337 | var424;
assign var426 = var338 & var350;
assign var427 = var341 & var352;
assign var428 = var340 | var427;
assign var429 = var341 & var353;
assign var430 = var344 & var355;
assign var431 = var343 | var430;
assign var432 = var344 & var356;
assign var433 = var347 & var358;
assign var434 = var346 | var433;
assign var435 = var347 & var359;
assign var436 = var350 & var361;
assign var437 = var349 | var436;
assign var438 = var350 & var362;
assign var439 = var353 & var364;
assign var440 = var352 | var439;
assign var441 = var353 & var365;
assign var442 = var356 & var367;
assign var443 = var355 | var442;
assign var444 = var356 & var368;
assign var445 = var359 & var370;
assign var446 = var358 | var445;
assign var447 = var359 & var371;
assign var448 = var362 & var373;
assign var449 = var361 | var448;
assign var450 = var362 & var374;
assign var451 = var365 & var376;
assign var452 = var364 | var451;
assign var453 = var365 & var377;
assign var454 = var368 & var379;
assign var455 = var367 | var454;
assign var456 = var368 & var380;
assign var457 = var371 & var382;
assign var458 = var370 | var457;
assign var459 = var371 & var383;
assign var460 = var374 & var385;
assign var461 = var373 | var460;
assign var462 = var374 & var386;
assign var463 = var377 & var388;
assign var464 = var376 | var463;
assign var465 = var377 & var389;
assign var466 = var380 & var391;
assign var467 = var379 | var466;
assign var468 = var380 & var392;
assign var469 = var383 & var394;
assign var470 = var382 | var469;
assign var471 = var383 & var395;
assign var472 = var386 & var397;
assign var473 = var385 | var472;
assign var474 = var386 & var398;
assign var475 = var389 & var400;
assign var476 = var388 | var475;
assign var477 = var392 & var402;
assign var478 = var391 | var477;
assign var479 = var395 & var314;
assign var480 = var394 | var479;
assign var481 = var398 & var222;
assign var482 = var397 | var481;
assign var483 = var405 & var428;
assign var484 = var404 | var483;
assign var485 = var405 & var429;
assign var486 = var408 & var431;
assign var487 = var407 | var486;
assign var488 = var408 & var432;
assign var489 = var411 & var434;
assign var490 = var410 | var489;
assign var491 = var411 & var435;
assign var492 = var414 & var437;
assign var493 = var413 | var492;
assign var494 = var414 & var438;
assign var495 = var417 & var440;
assign var496 = var416 | var495;
assign var497 = var417 & var441;
assign var498 = var420 & var443;
assign var499 = var419 | var498;
assign var500 = var420 & var444;
assign var501 = var423 & var446;
assign var502 = var422 | var501;
assign var503 = var423 & var447;
assign var504 = var426 & var449;
assign var505 = var425 | var504;
assign var506 = var426 & var450;
assign var507 = var429 & var452;
assign var508 = var428 | var507;
assign var509 = var429 & var453;
assign var510 = var432 & var455;
assign var511 = var431 | var510;
assign var512 = var432 & var456;
assign var513 = var435 & var458;
assign var514 = var434 | var513;
assign var515 = var435 & var459;
assign var516 = var438 & var461;
assign var517 = var437 | var516;
assign var518 = var438 & var462;
assign var519 = var441 & var464;
assign var520 = var440 | var519;
assign var521 = var441 & var465;
assign var522 = var444 & var467;
assign var523 = var443 | var522;
assign var524 = var444 & var468;
assign var525 = var447 & var470;
assign var526 = var446 | var525;
assign var527 = var447 & var471;
assign var528 = var450 & var473;
assign var529 = var449 | var528;
assign var530 = var450 & var474;
assign var531 = var453 & var476;
assign var532 = var452 | var531;
assign var533 = var456 & var478;
assign var534 = var455 | var533;
assign var535 = var459 & var480;
assign var536 = var458 | var535;
assign var537 = var462 & var482;
assign var538 = var461 | var537;
assign var539 = var465 & var400;
assign var540 = var464 | var539;
assign var541 = var468 & var402;
assign var542 = var467 | var541;
assign var543 = var471 & var314;
assign var544 = var470 | var543;
assign var545 = var474 & var222;
assign var546 = var473 | var545;
assign var547 = var485 & var532;
assign var548 = var484 | var547;
assign var549 = var488 & var534;
assign var550 = var487 | var549;
assign var551 = var491 & var536;
assign var552 = var490 | var551;
assign var553 = var494 & var538;
assign var554 = var493 | var553;
assign var555 = var497 & var540;
assign var556 = var496 | var555;
assign var557 = var500 & var542;
assign var558 = var499 | var557;
assign var559 = var503 & var544;
assign var560 = var502 | var559;
assign var561 = var506 & var546;
assign var562 = var505 | var561;
assign var563 = var509 & var476;
assign var564 = var508 | var563;
assign var565 = var512 & var478;
assign var566 = var511 | var565;
assign var567 = var515 & var480;
assign var568 = var514 | var567;
assign var569 = var518 & var482;
assign var570 = var517 | var569;
assign var571 = var521 & var400;
assign var572 = var520 | var571;
assign var573 = var524 & var402;
assign var574 = var523 | var573;
assign var575 = var527 & var314;
assign var576 = var526 | var575;
assign var577 = var530 & var222;
assign var578 = var529 | var577;
assign var579 = var126 & var550;
assign var580 = var62 | var579;
assign var581 = var126 & var488;
assign var582 = var124 & var552;
assign var583 = var60 | var582;
assign var584 = var124 & var491;
assign var585 = var122 & var554;
assign var586 = var58 | var585;
assign var587 = var122 & var494;
assign var588 = var120 & var556;
assign var589 = var56 | var588;
assign var590 = var120 & var497;
assign var591 = var118 & var558;
assign var592 = var54 | var591;
assign var593 = var118 & var500;
assign var594 = var116 & var560;
assign var595 = var52 | var594;
assign var596 = var116 & var503;
assign var597 = var114 & var562;
assign var598 = var50 | var597;
assign var599 = var114 & var506;
assign var600 = var112 & var564;
assign var601 = var48 | var600;
assign var602 = var112 & var509;
assign var603 = var110 & var566;
assign var604 = var46 | var603;
assign var605 = var110 & var512;
assign var606 = var108 & var568;
assign var607 = var44 | var606;
assign var608 = var108 & var515;
assign var609 = var106 & var570;
assign var610 = var42 | var609;
assign var611 = var106 & var518;
assign var612 = var104 & var572;
assign var613 = var40 | var612;
assign var614 = var104 & var521;
assign var615 = var102 & var574;
assign var616 = var38 | var615;
assign var617 = var102 & var524;
assign var618 = var100 & var576;
assign var619 = var36 | var618;
assign var620 = var100 & var527;
assign var621 = var98 & var578;
assign var622 = var34 | var621;
assign var623 = var98 & var530;
assign var624 = var96 & var532;
assign var625 = var32 | var624;
assign var626 = var96 & var453;
assign var627 = var94 & var534;
assign var628 = var30 | var627;
assign var629 = var94 & var456;
assign var630 = var92 & var536;
assign var631 = var28 | var630;
assign var632 = var92 & var459;
assign var633 = var90 & var538;
assign var634 = var26 | var633;
assign var635 = var90 & var462;
assign var636 = var88 & var540;
assign var637 = var24 | var636;
assign var638 = var88 & var465;
assign var639 = var86 & var542;
assign var640 = var22 | var639;
assign var641 = var86 & var468;
assign var642 = var84 & var544;
assign var643 = var20 | var642;
assign var644 = var84 & var471;
assign var645 = var82 & var546;
assign var646 = var18 | var645;
assign var647 = var82 & var474;
assign var648 = var80 & var476;
assign var649 = var16 | var648;
assign var650 = var80 & var389;
assign var651 = var78 & var478;
assign var652 = var14 | var651;
assign var653 = var78 & var392;
assign var654 = var76 & var480;
assign var655 = var12 | var654;
assign var656 = var76 & var395;
assign var657 = var74 & var482;
assign var658 = var10 | var657;
assign var659 = var74 & var398;
assign var660 = var72 & var400;
assign var661 = var8 | var660;
assign var662 = var72 & var309;
assign var663 = var70 & var402;
assign var664 = var6 | var663;
assign var665 = var70 & var312;
assign var666 = var68 & var314;
assign var667 = var4 | var666;
assign var668 = var68 & var220;
assign var669 = var66 & var222;
assign var670 = var2 | var669;
assign var671 = var66 & var65;
assign var672 = var65 ^ var0;
assign var673 = var66 ^ var222;
assign var674 = var67 ^ var670;
assign var675 = var68 ^ var314;
assign var676 = var69 ^ var667;
assign var677 = var70 ^ var402;
assign var678 = var71 ^ var664;
assign var679 = var72 ^ var400;
assign var680 = var73 ^ var661;
assign var681 = var74 ^ var482;
assign var682 = var75 ^ var658;
assign var683 = var76 ^ var480;
assign var684 = var77 ^ var655;
assign var685 = var78 ^ var478;
assign var686 = var79 ^ var652;
assign var687 = var80 ^ var476;
assign var688 = var81 ^ var649;
assign var689 = var82 ^ var546;
assign var690 = var83 ^ var646;
assign var691 = var84 ^ var544;
assign var692 = var85 ^ var643;
assign var693 = var86 ^ var542;
assign var694 = var87 ^ var640;
assign var695 = var88 ^ var540;
assign var696 = var89 ^ var637;
assign var697 = var90 ^ var538;
assign var698 = var91 ^ var634;
assign var699 = var92 ^ var536;
assign var700 = var93 ^ var631;
assign var701 = var94 ^ var534;
assign var702 = var95 ^ var628;
assign var703 = var96 ^ var532;
assign var704 = var97 ^ var625;
assign var705 = var98 ^ var578;
assign var706 = var99 ^ var622;
assign var707 = var100 ^ var576;
assign var708 = var101 ^ var619;
assign var709 = var102 ^ var574;
assign var710 = var103 ^ var616;
assign var711 = var104 ^ var572;
assign var712 = var105 ^ var613;
assign var713 = var106 ^ var570;
assign var714 = var107 ^ var610;
assign var715 = var108 ^ var568;
assign var716 = var109 ^ var607;
assign var717 = var110 ^ var566;
assign var718 = var111 ^ var604;
assign var719 = var112 ^ var564;
assign var720 = var113 ^ var601;
assign var721 = var114 ^ var562;
assign var722 = var115 ^ var598;
assign var723 = var116 ^ var560;
assign var724 = var117 ^ var595;
assign var725 = var118 ^ var558;
assign var726 = var119 ^ var592;
assign var727 = var120 ^ var556;
assign var728 = var121 ^ var589;
assign var729 = var122 ^ var554;
assign var730 = var123 ^ var586;
assign var731 = var124 ^ var552;
assign var732 = var125 ^ var583;
assign var733 = var126 ^ var550;
assign var734 = var127 ^ var580;
assign out0 = var548;
assign out1 = var734;
assign out2 = var733;
assign out3 = var732;
assign out4 = var731;
assign out5 = var730;
assign out6 = var729;
assign out7 = var728;
assign out8 = var727;
assign out9 = var726;
assign out10 = var725;
assign out11 = var724;
assign out12 = var723;
assign out13 = var722;
assign out14 = var721;
assign out15 = var720;
assign out16 = var719;
assign out17 = var718;
assign out18 = var717;
assign out19 = var716;
assign out20 = var715;
assign out21 = var714;
assign out22 = var713;
assign out23 = var712;
assign out24 = var711;
assign out25 = var710;
assign out26 = var709;
assign out27 = var708;
assign out28 = var707;
assign out29 = var706;
assign out30 = var705;
assign out31 = var704;
assign out32 = var703;
assign out33 = var702;
assign out34 = var701;
assign out35 = var700;
assign out36 = var699;
assign out37 = var698;
assign out38 = var697;
assign out39 = var696;
assign out40 = var695;
assign out41 = var694;
assign out42 = var693;
assign out43 = var692;
assign out44 = var691;
assign out45 = var690;
assign out46 = var689;
assign out47 = var688;
assign out48 = var687;
assign out49 = var686;
assign out50 = var685;
assign out51 = var684;
assign out52 = var683;
assign out53 = var682;
assign out54 = var681;
assign out55 = var680;
assign out56 = var679;
assign out57 = var678;
assign out58 = var677;
assign out59 = var676;
assign out60 = var675;
assign out61 = var674;
assign out62 = var673;
assign out63 = var672;
assign out64 = var64;
endmodule 
