module bk64 (in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, in100, in101, in102, in103, in104, in105, in106, in107, in108, in109, in110, in111, in112, in113, in114, in115, in116, in117, in118, in119, in120, in121, in122, in123, in124, in125, in126, in127, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, out30, out31, out32, out33, out34, out35, out36, out37, out38, out39, out40, out41, out42, out43, out44, out45, out46, out47, out48, out49, out50, out51, out52, out53, out54, out55, out56, out57, out58, out59, out60, out61, out62, out63, out64, );
input in0;
input in1;
input in2;
input in3;
input in4;
input in5;
input in6;
input in7;
input in8;
input in9;
input in10;
input in11;
input in12;
input in13;
input in14;
input in15;
input in16;
input in17;
input in18;
input in19;
input in20;
input in21;
input in22;
input in23;
input in24;
input in25;
input in26;
input in27;
input in28;
input in29;
input in30;
input in31;
input in32;
input in33;
input in34;
input in35;
input in36;
input in37;
input in38;
input in39;
input in40;
input in41;
input in42;
input in43;
input in44;
input in45;
input in46;
input in47;
input in48;
input in49;
input in50;
input in51;
input in52;
input in53;
input in54;
input in55;
input in56;
input in57;
input in58;
input in59;
input in60;
input in61;
input in62;
input in63;
input in64;
input in65;
input in66;
input in67;
input in68;
input in69;
input in70;
input in71;
input in72;
input in73;
input in74;
input in75;
input in76;
input in77;
input in78;
input in79;
input in80;
input in81;
input in82;
input in83;
input in84;
input in85;
input in86;
input in87;
input in88;
input in89;
input in90;
input in91;
input in92;
input in93;
input in94;
input in95;
input in96;
input in97;
input in98;
input in99;
input in100;
input in101;
input in102;
input in103;
input in104;
input in105;
input in106;
input in107;
input in108;
input in109;
input in110;
input in111;
input in112;
input in113;
input in114;
input in115;
input in116;
input in117;
input in118;
input in119;
input in120;
input in121;
input in122;
input in123;
input in124;
input in125;
input in126;
input in127;
output out0;
output out1;
output out2;
output out3;
output out4;
output out5;
output out6;
output out7;
output out8;
output out9;
output out10;
output out11;
output out12;
output out13;
output out14;
output out15;
output out16;
output out17;
output out18;
output out19;
output out20;
output out21;
output out22;
output out23;
output out24;
output out25;
output out26;
output out27;
output out28;
output out29;
output out30;
output out31;
output out32;
output out33;
output out34;
output out35;
output out36;
output out37;
output out38;
output out39;
output out40;
output out41;
output out42;
output out43;
output out44;
output out45;
output out46;
output out47;
output out48;
output out49;
output out50;
output out51;
output out52;
output out53;
output out54;
output out55;
output out56;
output out57;
output out58;
output out59;
output out60;
output out61;
output out62;
output out63;
output out64;
wire var0;
wire var1;
wire var2;
wire var3;
wire var4;
wire var5;
wire var6;
wire var7;
wire var8;
wire var9;
wire var10;
wire var11;
wire var12;
wire var13;
wire var14;
wire var15;
wire var16;
wire var17;
wire var18;
wire var19;
wire var20;
wire var21;
wire var22;
wire var23;
wire var24;
wire var25;
wire var26;
wire var27;
wire var28;
wire var29;
wire var30;
wire var31;
wire var32;
wire var33;
wire var34;
wire var35;
wire var36;
wire var37;
wire var38;
wire var39;
wire var40;
wire var41;
wire var42;
wire var43;
wire var44;
wire var45;
wire var46;
wire var47;
wire var48;
wire var49;
wire var50;
wire var51;
wire var52;
wire var53;
wire var54;
wire var55;
wire var56;
wire var57;
wire var58;
wire var59;
wire var60;
wire var61;
wire var62;
wire var63;
wire var64;
wire var65;
wire var66;
wire var67;
wire var68;
wire var69;
wire var70;
wire var71;
wire var72;
wire var73;
wire var74;
wire var75;
wire var76;
wire var77;
wire var78;
wire var79;
wire var80;
wire var81;
wire var82;
wire var83;
wire var84;
wire var85;
wire var86;
wire var87;
wire var88;
wire var89;
wire var90;
wire var91;
wire var92;
wire var93;
wire var94;
wire var95;
wire var96;
wire var97;
wire var98;
wire var99;
wire var100;
wire var101;
wire var102;
wire var103;
wire var104;
wire var105;
wire var106;
wire var107;
wire var108;
wire var109;
wire var110;
wire var111;
wire var112;
wire var113;
wire var114;
wire var115;
wire var116;
wire var117;
wire var118;
wire var119;
wire var120;
wire var121;
wire var122;
wire var123;
wire var124;
wire var125;
wire var126;
wire var127;
wire var128;
wire var129;
wire var130;
wire var131;
wire var132;
wire var133;
wire var134;
wire var135;
wire var136;
wire var137;
wire var138;
wire var139;
wire var140;
wire var141;
wire var142;
wire var143;
wire var144;
wire var145;
wire var146;
wire var147;
wire var148;
wire var149;
wire var150;
wire var151;
wire var152;
wire var153;
wire var154;
wire var155;
wire var156;
wire var157;
wire var158;
wire var159;
wire var160;
wire var161;
wire var162;
wire var163;
wire var164;
wire var165;
wire var166;
wire var167;
wire var168;
wire var169;
wire var170;
wire var171;
wire var172;
wire var173;
wire var174;
wire var175;
wire var176;
wire var177;
wire var178;
wire var179;
wire var180;
wire var181;
wire var182;
wire var183;
wire var184;
wire var185;
wire var186;
wire var187;
wire var188;
wire var189;
wire var190;
wire var191;
wire var192;
wire var193;
wire var194;
wire var195;
wire var196;
wire var197;
wire var198;
wire var199;
wire var200;
wire var201;
wire var202;
wire var203;
wire var204;
wire var205;
wire var206;
wire var207;
wire var208;
wire var209;
wire var210;
wire var211;
wire var212;
wire var213;
wire var214;
wire var215;
wire var216;
wire var217;
wire var218;
wire var219;
wire var220;
wire var221;
wire var222;
wire var223;
wire var224;
wire var225;
wire var226;
wire var227;
wire var228;
wire var229;
wire var230;
wire var231;
wire var232;
wire var233;
wire var234;
wire var235;
wire var236;
wire var237;
wire var238;
wire var239;
wire var240;
wire var241;
wire var242;
wire var243;
wire var244;
wire var245;
wire var246;
wire var247;
wire var248;
wire var249;
wire var250;
wire var251;
wire var252;
wire var253;
wire var254;
wire var255;
wire var256;
wire var257;
wire var258;
wire var259;
wire var260;
wire var261;
wire var262;
wire var263;
wire var264;
wire var265;
wire var266;
wire var267;
wire var268;
wire var269;
wire var270;
wire var271;
wire var272;
wire var273;
wire var274;
wire var275;
wire var276;
wire var277;
wire var278;
wire var279;
wire var280;
wire var281;
wire var282;
wire var283;
wire var284;
wire var285;
wire var286;
wire var287;
wire var288;
wire var289;
wire var290;
wire var291;
wire var292;
wire var293;
wire var294;
wire var295;
wire var296;
wire var297;
wire var298;
wire var299;
wire var300;
wire var301;
wire var302;
wire var303;
wire var304;
wire var305;
wire var306;
wire var307;
wire var308;
wire var309;
wire var310;
wire var311;
wire var312;
wire var313;
wire var314;
wire var315;
wire var316;
wire var317;
wire var318;
wire var319;
wire var320;
wire var321;
wire var322;
wire var323;
wire var324;
wire var325;
wire var326;
wire var327;
wire var328;
wire var329;
wire var330;
wire var331;
wire var332;
wire var333;
wire var334;
wire var335;
wire var336;
wire var337;
wire var338;
wire var339;
wire var340;
wire var341;
wire var342;
wire var343;
wire var344;
wire var345;
wire var346;
wire var347;
wire var348;
wire var349;
wire var350;
wire var351;
wire var352;
wire var353;
wire var354;
wire var355;
wire var356;
wire var357;
wire var358;
wire var359;
wire var360;
wire var361;
wire var362;
wire var363;
wire var364;
wire var365;
wire var366;
wire var367;
wire var368;
wire var369;
wire var370;
wire var371;
wire var372;
wire var373;
wire var374;
wire var375;
wire var376;
wire var377;
wire var378;
wire var379;
wire var380;
wire var381;
wire var382;
wire var383;
wire var384;
wire var385;
wire var386;
wire var387;
wire var388;
wire var389;
wire var390;
wire var391;
wire var392;
wire var393;
wire var394;
wire var395;
wire var396;
wire var397;
wire var398;
wire var399;
wire var400;
wire var401;
wire var402;
wire var403;
wire var404;
wire var405;
wire var406;
wire var407;
wire var408;
wire var409;
wire var410;
wire var411;
wire var412;
wire var413;
wire var414;
wire var415;
wire var416;
wire var417;
wire var418;
wire var419;
wire var420;
wire var421;
wire var422;
wire var423;
wire var424;
wire var425;
wire var426;
wire var427;
wire var428;
wire var429;
wire var430;
wire var431;
wire var432;
wire var433;
wire var434;
wire var435;
wire var436;
wire var437;
wire var438;
wire var439;
wire var440;
wire var441;
wire var442;
wire var443;
wire var444;
wire var445;
wire var446;
wire var447;
wire var448;
wire var449;
wire var450;
wire var451;
wire var452;
wire var453;
wire var454;
wire var455;
wire var456;
wire var457;
wire var458;
wire var459;
wire var460;
wire var461;
wire var462;
wire var463;
wire var464;
wire var465;
wire var466;
wire var467;
wire var468;
wire var469;
wire var470;
wire var471;
wire var472;
wire var473;
wire var474;
wire var475;
wire var476;
wire var477;
wire var478;
wire var479;
wire var480;
wire var481;
wire var482;
wire var483;
wire var484;
wire var485;
wire var486;
wire var487;
wire var488;
wire var489;
wire var490;
wire var491;
wire var492;
wire var493;
wire var494;
wire var495;
wire var496;
wire var497;
wire var498;
wire var499;
wire var500;
wire var501;
wire var502;
wire var503;
wire var504;
wire var505;
wire var506;
wire var507;
wire var508;
wire var509;
wire var510;
wire var511;
wire var512;
wire var513;
wire var514;
wire var515;
wire var516;
wire var517;
wire var518;
assign var0 = in127 & in63;
assign var1 = in126 & in62;
assign var2 = in125 & in61;
assign var3 = in124 & in60;
assign var4 = in123 & in59;
assign var5 = in122 & in58;
assign var6 = in121 & in57;
assign var7 = in120 & in56;
assign var8 = in119 & in55;
assign var9 = in118 & in54;
assign var10 = in117 & in53;
assign var11 = in116 & in52;
assign var12 = in115 & in51;
assign var13 = in114 & in50;
assign var14 = in113 & in49;
assign var15 = in112 & in48;
assign var16 = in111 & in47;
assign var17 = in110 & in46;
assign var18 = in109 & in45;
assign var19 = in108 & in44;
assign var20 = in107 & in43;
assign var21 = in106 & in42;
assign var22 = in105 & in41;
assign var23 = in104 & in40;
assign var24 = in103 & in39;
assign var25 = in102 & in38;
assign var26 = in101 & in37;
assign var27 = in100 & in36;
assign var28 = in99 & in35;
assign var29 = in98 & in34;
assign var30 = in97 & in33;
assign var31 = in96 & in32;
assign var32 = in95 & in31;
assign var33 = in94 & in30;
assign var34 = in93 & in29;
assign var35 = in92 & in28;
assign var36 = in91 & in27;
assign var37 = in90 & in26;
assign var38 = in89 & in25;
assign var39 = in88 & in24;
assign var40 = in87 & in23;
assign var41 = in86 & in22;
assign var42 = in85 & in21;
assign var43 = in84 & in20;
assign var44 = in83 & in19;
assign var45 = in82 & in18;
assign var46 = in81 & in17;
assign var47 = in80 & in16;
assign var48 = in79 & in15;
assign var49 = in78 & in14;
assign var50 = in77 & in13;
assign var51 = in76 & in12;
assign var52 = in75 & in11;
assign var53 = in74 & in10;
assign var54 = in73 & in9;
assign var55 = in72 & in8;
assign var56 = in71 & in7;
assign var57 = in70 & in6;
assign var58 = in69 & in5;
assign var59 = in68 & in4;
assign var60 = in67 & in3;
assign var61 = in66 & in2;
assign var62 = in65 & in1;
assign var63 = in64 & in0;
assign var64 = in127 ^ in63;
assign var65 = in126 ^ in62;
assign var66 = in125 ^ in61;
assign var67 = in124 ^ in60;
assign var68 = in123 ^ in59;
assign var69 = in122 ^ in58;
assign var70 = in121 ^ in57;
assign var71 = in120 ^ in56;
assign var72 = in119 ^ in55;
assign var73 = in118 ^ in54;
assign var74 = in117 ^ in53;
assign var75 = in116 ^ in52;
assign var76 = in115 ^ in51;
assign var77 = in114 ^ in50;
assign var78 = in113 ^ in49;
assign var79 = in112 ^ in48;
assign var80 = in111 ^ in47;
assign var81 = in110 ^ in46;
assign var82 = in109 ^ in45;
assign var83 = in108 ^ in44;
assign var84 = in107 ^ in43;
assign var85 = in106 ^ in42;
assign var86 = in105 ^ in41;
assign var87 = in104 ^ in40;
assign var88 = in103 ^ in39;
assign var89 = in102 ^ in38;
assign var90 = in101 ^ in37;
assign var91 = in100 ^ in36;
assign var92 = in99 ^ in35;
assign var93 = in98 ^ in34;
assign var94 = in97 ^ in33;
assign var95 = in96 ^ in32;
assign var96 = in95 ^ in31;
assign var97 = in94 ^ in30;
assign var98 = in93 ^ in29;
assign var99 = in92 ^ in28;
assign var100 = in91 ^ in27;
assign var101 = in90 ^ in26;
assign var102 = in89 ^ in25;
assign var103 = in88 ^ in24;
assign var104 = in87 ^ in23;
assign var105 = in86 ^ in22;
assign var106 = in85 ^ in21;
assign var107 = in84 ^ in20;
assign var108 = in83 ^ in19;
assign var109 = in82 ^ in18;
assign var110 = in81 ^ in17;
assign var111 = in80 ^ in16;
assign var112 = in79 ^ in15;
assign var113 = in78 ^ in14;
assign var114 = in77 ^ in13;
assign var115 = in76 ^ in12;
assign var116 = in75 ^ in11;
assign var117 = in74 ^ in10;
assign var118 = in73 ^ in9;
assign var119 = in72 ^ in8;
assign var120 = in71 ^ in7;
assign var121 = in70 ^ in6;
assign var122 = in69 ^ in5;
assign var123 = in68 ^ in4;
assign var124 = in67 ^ in3;
assign var125 = in66 ^ in2;
assign var126 = in65 ^ in1;
assign var127 = in64 ^ in0;
assign var128 = var127 & var62;
assign var129 = var63 | var128;
assign var130 = var127 & var126;
assign var131 = var125 & var60;
assign var132 = var61 | var131;
assign var133 = var125 & var124;
assign var134 = var123 & var58;
assign var135 = var59 | var134;
assign var136 = var123 & var122;
assign var137 = var121 & var56;
assign var138 = var57 | var137;
assign var139 = var121 & var120;
assign var140 = var119 & var54;
assign var141 = var55 | var140;
assign var142 = var119 & var118;
assign var143 = var117 & var52;
assign var144 = var53 | var143;
assign var145 = var117 & var116;
assign var146 = var115 & var50;
assign var147 = var51 | var146;
assign var148 = var115 & var114;
assign var149 = var113 & var48;
assign var150 = var49 | var149;
assign var151 = var113 & var112;
assign var152 = var111 & var46;
assign var153 = var47 | var152;
assign var154 = var111 & var110;
assign var155 = var109 & var44;
assign var156 = var45 | var155;
assign var157 = var109 & var108;
assign var158 = var107 & var42;
assign var159 = var43 | var158;
assign var160 = var107 & var106;
assign var161 = var105 & var40;
assign var162 = var41 | var161;
assign var163 = var105 & var104;
assign var164 = var103 & var38;
assign var165 = var39 | var164;
assign var166 = var103 & var102;
assign var167 = var101 & var36;
assign var168 = var37 | var167;
assign var169 = var101 & var100;
assign var170 = var99 & var34;
assign var171 = var35 | var170;
assign var172 = var99 & var98;
assign var173 = var97 & var32;
assign var174 = var33 | var173;
assign var175 = var97 & var96;
assign var176 = var95 & var30;
assign var177 = var31 | var176;
assign var178 = var95 & var94;
assign var179 = var93 & var28;
assign var180 = var29 | var179;
assign var181 = var93 & var92;
assign var182 = var91 & var26;
assign var183 = var27 | var182;
assign var184 = var91 & var90;
assign var185 = var89 & var24;
assign var186 = var25 | var185;
assign var187 = var89 & var88;
assign var188 = var87 & var22;
assign var189 = var23 | var188;
assign var190 = var87 & var86;
assign var191 = var85 & var20;
assign var192 = var21 | var191;
assign var193 = var85 & var84;
assign var194 = var83 & var18;
assign var195 = var19 | var194;
assign var196 = var83 & var82;
assign var197 = var81 & var16;
assign var198 = var17 | var197;
assign var199 = var81 & var80;
assign var200 = var79 & var14;
assign var201 = var15 | var200;
assign var202 = var79 & var78;
assign var203 = var77 & var12;
assign var204 = var13 | var203;
assign var205 = var77 & var76;
assign var206 = var75 & var10;
assign var207 = var11 | var206;
assign var208 = var75 & var74;
assign var209 = var73 & var8;
assign var210 = var9 | var209;
assign var211 = var73 & var72;
assign var212 = var71 & var6;
assign var213 = var7 | var212;
assign var214 = var71 & var70;
assign var215 = var69 & var4;
assign var216 = var5 | var215;
assign var217 = var69 & var68;
assign var218 = var67 & var2;
assign var219 = var3 | var218;
assign var220 = var67 & var66;
assign var221 = var65 & var0;
assign var222 = var1 | var221;
assign var223 = var130 & var132;
assign var224 = var129 | var223;
assign var225 = var130 & var133;
assign var226 = var136 & var138;
assign var227 = var135 | var226;
assign var228 = var136 & var139;
assign var229 = var142 & var144;
assign var230 = var141 | var229;
assign var231 = var142 & var145;
assign var232 = var148 & var150;
assign var233 = var147 | var232;
assign var234 = var148 & var151;
assign var235 = var154 & var156;
assign var236 = var153 | var235;
assign var237 = var154 & var157;
assign var238 = var160 & var162;
assign var239 = var159 | var238;
assign var240 = var160 & var163;
assign var241 = var166 & var168;
assign var242 = var165 | var241;
assign var243 = var166 & var169;
assign var244 = var172 & var174;
assign var245 = var171 | var244;
assign var246 = var172 & var175;
assign var247 = var178 & var180;
assign var248 = var177 | var247;
assign var249 = var178 & var181;
assign var250 = var184 & var186;
assign var251 = var183 | var250;
assign var252 = var184 & var187;
assign var253 = var190 & var192;
assign var254 = var189 | var253;
assign var255 = var190 & var193;
assign var256 = var196 & var198;
assign var257 = var195 | var256;
assign var258 = var196 & var199;
assign var259 = var202 & var204;
assign var260 = var201 | var259;
assign var261 = var202 & var205;
assign var262 = var208 & var210;
assign var263 = var207 | var262;
assign var264 = var208 & var211;
assign var265 = var214 & var216;
assign var266 = var213 | var265;
assign var267 = var214 & var217;
assign var268 = var220 & var222;
assign var269 = var219 | var268;
assign var270 = var225 & var227;
assign var271 = var224 | var270;
assign var272 = var225 & var228;
assign var273 = var231 & var233;
assign var274 = var230 | var273;
assign var275 = var231 & var234;
assign var276 = var237 & var239;
assign var277 = var236 | var276;
assign var278 = var237 & var240;
assign var279 = var243 & var245;
assign var280 = var242 | var279;
assign var281 = var243 & var246;
assign var282 = var249 & var251;
assign var283 = var248 | var282;
assign var284 = var249 & var252;
assign var285 = var255 & var257;
assign var286 = var254 | var285;
assign var287 = var255 & var258;
assign var288 = var261 & var263;
assign var289 = var260 | var288;
assign var290 = var261 & var264;
assign var291 = var267 & var269;
assign var292 = var266 | var291;
assign var293 = var272 & var274;
assign var294 = var271 | var293;
assign var295 = var272 & var275;
assign var296 = var278 & var280;
assign var297 = var277 | var296;
assign var298 = var278 & var281;
assign var299 = var284 & var286;
assign var300 = var283 | var299;
assign var301 = var284 & var287;
assign var302 = var290 & var292;
assign var303 = var289 | var302;
assign var304 = var295 & var297;
assign var305 = var294 | var304;
assign var306 = var295 & var298;
assign var307 = var301 & var303;
assign var308 = var300 | var307;
assign var309 = var306 & var308;
assign var310 = var305 | var309;
assign var311 = var298 & var308;
assign var312 = var297 | var311;
assign var313 = var275 & var312;
assign var314 = var274 | var313;
assign var315 = var281 & var308;
assign var316 = var280 | var315;
assign var317 = var287 & var303;
assign var318 = var286 | var317;
assign var319 = var228 & var314;
assign var320 = var227 | var319;
assign var321 = var234 & var312;
assign var322 = var233 | var321;
assign var323 = var240 & var316;
assign var324 = var239 | var323;
assign var325 = var246 & var308;
assign var326 = var245 | var325;
assign var327 = var252 & var318;
assign var328 = var251 | var327;
assign var329 = var258 & var303;
assign var330 = var257 | var329;
assign var331 = var264 & var292;
assign var332 = var263 | var331;
assign var333 = var133 & var320;
assign var334 = var132 | var333;
assign var335 = var139 & var314;
assign var336 = var138 | var335;
assign var337 = var145 & var322;
assign var338 = var144 | var337;
assign var339 = var151 & var312;
assign var340 = var150 | var339;
assign var341 = var157 & var324;
assign var342 = var156 | var341;
assign var343 = var163 & var316;
assign var344 = var162 | var343;
assign var345 = var169 & var326;
assign var346 = var168 | var345;
assign var347 = var175 & var308;
assign var348 = var174 | var347;
assign var349 = var181 & var328;
assign var350 = var180 | var349;
assign var351 = var187 & var318;
assign var352 = var186 | var351;
assign var353 = var193 & var330;
assign var354 = var192 | var353;
assign var355 = var199 & var303;
assign var356 = var198 | var355;
assign var357 = var205 & var332;
assign var358 = var204 | var357;
assign var359 = var211 & var292;
assign var360 = var210 | var359;
assign var361 = var217 & var269;
assign var362 = var216 | var361;
assign var363 = var126 & var334;
assign var364 = var62 | var363;
assign var365 = var126 & var133;
assign var366 = var124 & var320;
assign var367 = var60 | var366;
assign var368 = var124 & var228;
assign var369 = var122 & var336;
assign var370 = var58 | var369;
assign var371 = var122 & var139;
assign var372 = var120 & var314;
assign var373 = var56 | var372;
assign var374 = var120 & var275;
assign var375 = var118 & var338;
assign var376 = var54 | var375;
assign var377 = var118 & var145;
assign var378 = var116 & var322;
assign var379 = var52 | var378;
assign var380 = var116 & var234;
assign var381 = var114 & var340;
assign var382 = var50 | var381;
assign var383 = var114 & var151;
assign var384 = var112 & var312;
assign var385 = var48 | var384;
assign var386 = var112 & var298;
assign var387 = var110 & var342;
assign var388 = var46 | var387;
assign var389 = var110 & var157;
assign var390 = var108 & var324;
assign var391 = var44 | var390;
assign var392 = var108 & var240;
assign var393 = var106 & var344;
assign var394 = var42 | var393;
assign var395 = var106 & var163;
assign var396 = var104 & var316;
assign var397 = var40 | var396;
assign var398 = var104 & var281;
assign var399 = var102 & var346;
assign var400 = var38 | var399;
assign var401 = var102 & var169;
assign var402 = var100 & var326;
assign var403 = var36 | var402;
assign var404 = var100 & var246;
assign var405 = var98 & var348;
assign var406 = var34 | var405;
assign var407 = var98 & var175;
assign var408 = var96 & var308;
assign var409 = var32 | var408;
assign var410 = var96 & var301;
assign var411 = var94 & var350;
assign var412 = var30 | var411;
assign var413 = var94 & var181;
assign var414 = var92 & var328;
assign var415 = var28 | var414;
assign var416 = var92 & var252;
assign var417 = var90 & var352;
assign var418 = var26 | var417;
assign var419 = var90 & var187;
assign var420 = var88 & var318;
assign var421 = var24 | var420;
assign var422 = var88 & var287;
assign var423 = var86 & var354;
assign var424 = var22 | var423;
assign var425 = var86 & var193;
assign var426 = var84 & var330;
assign var427 = var20 | var426;
assign var428 = var84 & var258;
assign var429 = var82 & var356;
assign var430 = var18 | var429;
assign var431 = var82 & var199;
assign var432 = var80 & var303;
assign var433 = var16 | var432;
assign var434 = var80 & var290;
assign var435 = var78 & var358;
assign var436 = var14 | var435;
assign var437 = var78 & var205;
assign var438 = var76 & var332;
assign var439 = var12 | var438;
assign var440 = var76 & var264;
assign var441 = var74 & var360;
assign var442 = var10 | var441;
assign var443 = var74 & var211;
assign var444 = var72 & var292;
assign var445 = var8 | var444;
assign var446 = var72 & var267;
assign var447 = var70 & var362;
assign var448 = var6 | var447;
assign var449 = var70 & var217;
assign var450 = var68 & var269;
assign var451 = var4 | var450;
assign var452 = var68 & var220;
assign var453 = var66 & var222;
assign var454 = var2 | var453;
assign var455 = var66 & var65;
assign var456 = var65 ^ var0;
assign var457 = var66 ^ var222;
assign var458 = var67 ^ var454;
assign var459 = var68 ^ var269;
assign var460 = var69 ^ var451;
assign var461 = var70 ^ var362;
assign var462 = var71 ^ var448;
assign var463 = var72 ^ var292;
assign var464 = var73 ^ var445;
assign var465 = var74 ^ var360;
assign var466 = var75 ^ var442;
assign var467 = var76 ^ var332;
assign var468 = var77 ^ var439;
assign var469 = var78 ^ var358;
assign var470 = var79 ^ var436;
assign var471 = var80 ^ var303;
assign var472 = var81 ^ var433;
assign var473 = var82 ^ var356;
assign var474 = var83 ^ var430;
assign var475 = var84 ^ var330;
assign var476 = var85 ^ var427;
assign var477 = var86 ^ var354;
assign var478 = var87 ^ var424;
assign var479 = var88 ^ var318;
assign var480 = var89 ^ var421;
assign var481 = var90 ^ var352;
assign var482 = var91 ^ var418;
assign var483 = var92 ^ var328;
assign var484 = var93 ^ var415;
assign var485 = var94 ^ var350;
assign var486 = var95 ^ var412;
assign var487 = var96 ^ var308;
assign var488 = var97 ^ var409;
assign var489 = var98 ^ var348;
assign var490 = var99 ^ var406;
assign var491 = var100 ^ var326;
assign var492 = var101 ^ var403;
assign var493 = var102 ^ var346;
assign var494 = var103 ^ var400;
assign var495 = var104 ^ var316;
assign var496 = var105 ^ var397;
assign var497 = var106 ^ var344;
assign var498 = var107 ^ var394;
assign var499 = var108 ^ var324;
assign var500 = var109 ^ var391;
assign var501 = var110 ^ var342;
assign var502 = var111 ^ var388;
assign var503 = var112 ^ var312;
assign var504 = var113 ^ var385;
assign var505 = var114 ^ var340;
assign var506 = var115 ^ var382;
assign var507 = var116 ^ var322;
assign var508 = var117 ^ var379;
assign var509 = var118 ^ var338;
assign var510 = var119 ^ var376;
assign var511 = var120 ^ var314;
assign var512 = var121 ^ var373;
assign var513 = var122 ^ var336;
assign var514 = var123 ^ var370;
assign var515 = var124 ^ var320;
assign var516 = var125 ^ var367;
assign var517 = var126 ^ var334;
assign var518 = var127 ^ var364;
assign out0 = var310;
assign out1 = var518;
assign out2 = var517;
assign out3 = var516;
assign out4 = var515;
assign out5 = var514;
assign out6 = var513;
assign out7 = var512;
assign out8 = var511;
assign out9 = var510;
assign out10 = var509;
assign out11 = var508;
assign out12 = var507;
assign out13 = var506;
assign out14 = var505;
assign out15 = var504;
assign out16 = var503;
assign out17 = var502;
assign out18 = var501;
assign out19 = var500;
assign out20 = var499;
assign out21 = var498;
assign out22 = var497;
assign out23 = var496;
assign out24 = var495;
assign out25 = var494;
assign out26 = var493;
assign out27 = var492;
assign out28 = var491;
assign out29 = var490;
assign out30 = var489;
assign out31 = var488;
assign out32 = var487;
assign out33 = var486;
assign out34 = var485;
assign out35 = var484;
assign out36 = var483;
assign out37 = var482;
assign out38 = var481;
assign out39 = var480;
assign out40 = var479;
assign out41 = var478;
assign out42 = var477;
assign out43 = var476;
assign out44 = var475;
assign out45 = var474;
assign out46 = var473;
assign out47 = var472;
assign out48 = var471;
assign out49 = var470;
assign out50 = var469;
assign out51 = var468;
assign out52 = var467;
assign out53 = var466;
assign out54 = var465;
assign out55 = var464;
assign out56 = var463;
assign out57 = var462;
assign out58 = var461;
assign out59 = var460;
assign out60 = var459;
assign out61 = var458;
assign out62 = var457;
assign out63 = var456;
assign out64 = var64;
endmodule 
