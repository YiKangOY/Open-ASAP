module PartialProd(
  input  [31:0] io_multiplicand,
  input  [31:0] io_multiplier,
  output [31:0] io_outs_0,
  output [31:0] io_outs_1,
  output [31:0] io_outs_2,
  output [31:0] io_outs_3,
  output [31:0] io_outs_4,
  output [31:0] io_outs_5,
  output [31:0] io_outs_6,
  output [31:0] io_outs_7,
  output [31:0] io_outs_8,
  output [31:0] io_outs_9,
  output [31:0] io_outs_10,
  output [31:0] io_outs_11,
  output [31:0] io_outs_12,
  output [31:0] io_outs_13,
  output [31:0] io_outs_14,
  output [31:0] io_outs_15,
  output [31:0] io_outs_16,
  output [31:0] io_outs_17,
  output [31:0] io_outs_18,
  output [31:0] io_outs_19,
  output [31:0] io_outs_20,
  output [31:0] io_outs_21,
  output [31:0] io_outs_22,
  output [31:0] io_outs_23,
  output [31:0] io_outs_24,
  output [31:0] io_outs_25,
  output [31:0] io_outs_26,
  output [31:0] io_outs_27,
  output [31:0] io_outs_28,
  output [31:0] io_outs_29,
  output [31:0] io_outs_30,
  output [31:0] io_outs_31
);
  wire  _T_34 = io_multiplicand[0] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_37 = io_multiplicand[1] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_40 = io_multiplicand[2] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_43 = io_multiplicand[3] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_46 = io_multiplicand[4] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_49 = io_multiplicand[5] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_52 = io_multiplicand[6] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_55 = io_multiplicand[7] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_58 = io_multiplicand[8] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_61 = io_multiplicand[9] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_64 = io_multiplicand[10] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_67 = io_multiplicand[11] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_70 = io_multiplicand[12] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_73 = io_multiplicand[13] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_76 = io_multiplicand[14] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_79 = io_multiplicand[15] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_82 = io_multiplicand[16] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_85 = io_multiplicand[17] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_88 = io_multiplicand[18] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_91 = io_multiplicand[19] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_94 = io_multiplicand[20] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_97 = io_multiplicand[21] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_100 = io_multiplicand[22] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_103 = io_multiplicand[23] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_106 = io_multiplicand[24] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_109 = io_multiplicand[25] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_112 = io_multiplicand[26] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_115 = io_multiplicand[27] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_118 = io_multiplicand[28] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_121 = io_multiplicand[29] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_124 = io_multiplicand[30] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_127 = io_multiplicand[31] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire [9:0] _T_136 = {_T_127,_T_124,_T_121,_T_118,_T_115,_T_112,_T_109,_T_106,_T_103,_T_100}; // @[Cat.scala 29:58]
  wire [18:0] _T_145 = {_T_136,_T_97,_T_94,_T_91,_T_88,_T_85,_T_82,_T_79,_T_76,_T_73}; // @[Cat.scala 29:58]
  wire [27:0] _T_154 = {_T_145,_T_70,_T_67,_T_64,_T_61,_T_58,_T_55,_T_52,_T_49,_T_46}; // @[Cat.scala 29:58]
  wire [30:0] _T_157 = {_T_154,_T_43,_T_40,_T_37}; // @[Cat.scala 29:58]
  wire  _T_193 = io_multiplicand[0] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_196 = io_multiplicand[1] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_199 = io_multiplicand[2] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_202 = io_multiplicand[3] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_205 = io_multiplicand[4] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_208 = io_multiplicand[5] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_211 = io_multiplicand[6] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_214 = io_multiplicand[7] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_217 = io_multiplicand[8] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_220 = io_multiplicand[9] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_223 = io_multiplicand[10] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_226 = io_multiplicand[11] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_229 = io_multiplicand[12] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_232 = io_multiplicand[13] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_235 = io_multiplicand[14] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_238 = io_multiplicand[15] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_241 = io_multiplicand[16] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_244 = io_multiplicand[17] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_247 = io_multiplicand[18] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_250 = io_multiplicand[19] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_253 = io_multiplicand[20] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_256 = io_multiplicand[21] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_259 = io_multiplicand[22] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_262 = io_multiplicand[23] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_265 = io_multiplicand[24] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_268 = io_multiplicand[25] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_271 = io_multiplicand[26] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_274 = io_multiplicand[27] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_277 = io_multiplicand[28] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_280 = io_multiplicand[29] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_283 = io_multiplicand[30] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_286 = io_multiplicand[31] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire [9:0] _T_295 = {_T_286,_T_283,_T_280,_T_277,_T_274,_T_271,_T_268,_T_265,_T_262,_T_259}; // @[Cat.scala 29:58]
  wire [18:0] _T_304 = {_T_295,_T_256,_T_253,_T_250,_T_247,_T_244,_T_241,_T_238,_T_235,_T_232}; // @[Cat.scala 29:58]
  wire [27:0] _T_313 = {_T_304,_T_229,_T_226,_T_223,_T_220,_T_217,_T_214,_T_211,_T_208,_T_205}; // @[Cat.scala 29:58]
  wire [30:0] _T_316 = {_T_313,_T_202,_T_199,_T_196}; // @[Cat.scala 29:58]
  wire  _T_352 = io_multiplicand[0] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_355 = io_multiplicand[1] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_358 = io_multiplicand[2] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_361 = io_multiplicand[3] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_364 = io_multiplicand[4] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_367 = io_multiplicand[5] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_370 = io_multiplicand[6] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_373 = io_multiplicand[7] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_376 = io_multiplicand[8] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_379 = io_multiplicand[9] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_382 = io_multiplicand[10] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_385 = io_multiplicand[11] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_388 = io_multiplicand[12] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_391 = io_multiplicand[13] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_394 = io_multiplicand[14] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_397 = io_multiplicand[15] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_400 = io_multiplicand[16] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_403 = io_multiplicand[17] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_406 = io_multiplicand[18] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_409 = io_multiplicand[19] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_412 = io_multiplicand[20] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_415 = io_multiplicand[21] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_418 = io_multiplicand[22] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_421 = io_multiplicand[23] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_424 = io_multiplicand[24] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_427 = io_multiplicand[25] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_430 = io_multiplicand[26] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_433 = io_multiplicand[27] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_436 = io_multiplicand[28] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_439 = io_multiplicand[29] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_442 = io_multiplicand[30] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_445 = io_multiplicand[31] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire [9:0] _T_454 = {_T_445,_T_442,_T_439,_T_436,_T_433,_T_430,_T_427,_T_424,_T_421,_T_418}; // @[Cat.scala 29:58]
  wire [18:0] _T_463 = {_T_454,_T_415,_T_412,_T_409,_T_406,_T_403,_T_400,_T_397,_T_394,_T_391}; // @[Cat.scala 29:58]
  wire [27:0] _T_472 = {_T_463,_T_388,_T_385,_T_382,_T_379,_T_376,_T_373,_T_370,_T_367,_T_364}; // @[Cat.scala 29:58]
  wire [30:0] _T_475 = {_T_472,_T_361,_T_358,_T_355}; // @[Cat.scala 29:58]
  wire  _T_511 = io_multiplicand[0] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_514 = io_multiplicand[1] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_517 = io_multiplicand[2] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_520 = io_multiplicand[3] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_523 = io_multiplicand[4] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_526 = io_multiplicand[5] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_529 = io_multiplicand[6] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_532 = io_multiplicand[7] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_535 = io_multiplicand[8] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_538 = io_multiplicand[9] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_541 = io_multiplicand[10] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_544 = io_multiplicand[11] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_547 = io_multiplicand[12] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_550 = io_multiplicand[13] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_553 = io_multiplicand[14] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_556 = io_multiplicand[15] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_559 = io_multiplicand[16] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_562 = io_multiplicand[17] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_565 = io_multiplicand[18] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_568 = io_multiplicand[19] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_571 = io_multiplicand[20] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_574 = io_multiplicand[21] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_577 = io_multiplicand[22] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_580 = io_multiplicand[23] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_583 = io_multiplicand[24] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_586 = io_multiplicand[25] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_589 = io_multiplicand[26] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_592 = io_multiplicand[27] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_595 = io_multiplicand[28] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_598 = io_multiplicand[29] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_601 = io_multiplicand[30] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_604 = io_multiplicand[31] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire [9:0] _T_613 = {_T_604,_T_601,_T_598,_T_595,_T_592,_T_589,_T_586,_T_583,_T_580,_T_577}; // @[Cat.scala 29:58]
  wire [18:0] _T_622 = {_T_613,_T_574,_T_571,_T_568,_T_565,_T_562,_T_559,_T_556,_T_553,_T_550}; // @[Cat.scala 29:58]
  wire [27:0] _T_631 = {_T_622,_T_547,_T_544,_T_541,_T_538,_T_535,_T_532,_T_529,_T_526,_T_523}; // @[Cat.scala 29:58]
  wire [30:0] _T_634 = {_T_631,_T_520,_T_517,_T_514}; // @[Cat.scala 29:58]
  wire  _T_670 = io_multiplicand[0] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_673 = io_multiplicand[1] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_676 = io_multiplicand[2] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_679 = io_multiplicand[3] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_682 = io_multiplicand[4] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_685 = io_multiplicand[5] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_688 = io_multiplicand[6] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_691 = io_multiplicand[7] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_694 = io_multiplicand[8] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_697 = io_multiplicand[9] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_700 = io_multiplicand[10] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_703 = io_multiplicand[11] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_706 = io_multiplicand[12] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_709 = io_multiplicand[13] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_712 = io_multiplicand[14] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_715 = io_multiplicand[15] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_718 = io_multiplicand[16] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_721 = io_multiplicand[17] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_724 = io_multiplicand[18] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_727 = io_multiplicand[19] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_730 = io_multiplicand[20] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_733 = io_multiplicand[21] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_736 = io_multiplicand[22] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_739 = io_multiplicand[23] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_742 = io_multiplicand[24] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_745 = io_multiplicand[25] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_748 = io_multiplicand[26] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_751 = io_multiplicand[27] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_754 = io_multiplicand[28] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_757 = io_multiplicand[29] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_760 = io_multiplicand[30] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_763 = io_multiplicand[31] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire [9:0] _T_772 = {_T_763,_T_760,_T_757,_T_754,_T_751,_T_748,_T_745,_T_742,_T_739,_T_736}; // @[Cat.scala 29:58]
  wire [18:0] _T_781 = {_T_772,_T_733,_T_730,_T_727,_T_724,_T_721,_T_718,_T_715,_T_712,_T_709}; // @[Cat.scala 29:58]
  wire [27:0] _T_790 = {_T_781,_T_706,_T_703,_T_700,_T_697,_T_694,_T_691,_T_688,_T_685,_T_682}; // @[Cat.scala 29:58]
  wire [30:0] _T_793 = {_T_790,_T_679,_T_676,_T_673}; // @[Cat.scala 29:58]
  wire  _T_829 = io_multiplicand[0] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_832 = io_multiplicand[1] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_835 = io_multiplicand[2] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_838 = io_multiplicand[3] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_841 = io_multiplicand[4] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_844 = io_multiplicand[5] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_847 = io_multiplicand[6] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_850 = io_multiplicand[7] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_853 = io_multiplicand[8] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_856 = io_multiplicand[9] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_859 = io_multiplicand[10] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_862 = io_multiplicand[11] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_865 = io_multiplicand[12] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_868 = io_multiplicand[13] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_871 = io_multiplicand[14] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_874 = io_multiplicand[15] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_877 = io_multiplicand[16] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_880 = io_multiplicand[17] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_883 = io_multiplicand[18] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_886 = io_multiplicand[19] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_889 = io_multiplicand[20] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_892 = io_multiplicand[21] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_895 = io_multiplicand[22] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_898 = io_multiplicand[23] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_901 = io_multiplicand[24] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_904 = io_multiplicand[25] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_907 = io_multiplicand[26] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_910 = io_multiplicand[27] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_913 = io_multiplicand[28] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_916 = io_multiplicand[29] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_919 = io_multiplicand[30] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_922 = io_multiplicand[31] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire [9:0] _T_931 = {_T_922,_T_919,_T_916,_T_913,_T_910,_T_907,_T_904,_T_901,_T_898,_T_895}; // @[Cat.scala 29:58]
  wire [18:0] _T_940 = {_T_931,_T_892,_T_889,_T_886,_T_883,_T_880,_T_877,_T_874,_T_871,_T_868}; // @[Cat.scala 29:58]
  wire [27:0] _T_949 = {_T_940,_T_865,_T_862,_T_859,_T_856,_T_853,_T_850,_T_847,_T_844,_T_841}; // @[Cat.scala 29:58]
  wire [30:0] _T_952 = {_T_949,_T_838,_T_835,_T_832}; // @[Cat.scala 29:58]
  wire  _T_988 = io_multiplicand[0] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_991 = io_multiplicand[1] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_994 = io_multiplicand[2] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_997 = io_multiplicand[3] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1000 = io_multiplicand[4] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1003 = io_multiplicand[5] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1006 = io_multiplicand[6] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1009 = io_multiplicand[7] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1012 = io_multiplicand[8] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1015 = io_multiplicand[9] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1018 = io_multiplicand[10] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1021 = io_multiplicand[11] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1024 = io_multiplicand[12] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1027 = io_multiplicand[13] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1030 = io_multiplicand[14] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1033 = io_multiplicand[15] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1036 = io_multiplicand[16] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1039 = io_multiplicand[17] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1042 = io_multiplicand[18] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1045 = io_multiplicand[19] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1048 = io_multiplicand[20] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1051 = io_multiplicand[21] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1054 = io_multiplicand[22] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1057 = io_multiplicand[23] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1060 = io_multiplicand[24] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1063 = io_multiplicand[25] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1066 = io_multiplicand[26] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1069 = io_multiplicand[27] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1072 = io_multiplicand[28] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1075 = io_multiplicand[29] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1078 = io_multiplicand[30] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1081 = io_multiplicand[31] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1090 = {_T_1081,_T_1078,_T_1075,_T_1072,_T_1069,_T_1066,_T_1063,_T_1060,_T_1057,_T_1054}; // @[Cat.scala 29:58]
  wire [18:0] _T_1099 = {_T_1090,_T_1051,_T_1048,_T_1045,_T_1042,_T_1039,_T_1036,_T_1033,_T_1030,_T_1027}; // @[Cat.scala 29:58]
  wire [27:0] _T_1108 = {_T_1099,_T_1024,_T_1021,_T_1018,_T_1015,_T_1012,_T_1009,_T_1006,_T_1003,_T_1000}; // @[Cat.scala 29:58]
  wire [30:0] _T_1111 = {_T_1108,_T_997,_T_994,_T_991}; // @[Cat.scala 29:58]
  wire  _T_1147 = io_multiplicand[0] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1150 = io_multiplicand[1] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1153 = io_multiplicand[2] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1156 = io_multiplicand[3] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1159 = io_multiplicand[4] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1162 = io_multiplicand[5] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1165 = io_multiplicand[6] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1168 = io_multiplicand[7] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1171 = io_multiplicand[8] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1174 = io_multiplicand[9] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1177 = io_multiplicand[10] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1180 = io_multiplicand[11] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1183 = io_multiplicand[12] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1186 = io_multiplicand[13] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1189 = io_multiplicand[14] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1192 = io_multiplicand[15] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1195 = io_multiplicand[16] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1198 = io_multiplicand[17] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1201 = io_multiplicand[18] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1204 = io_multiplicand[19] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1207 = io_multiplicand[20] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1210 = io_multiplicand[21] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1213 = io_multiplicand[22] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1216 = io_multiplicand[23] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1219 = io_multiplicand[24] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1222 = io_multiplicand[25] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1225 = io_multiplicand[26] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1228 = io_multiplicand[27] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1231 = io_multiplicand[28] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1234 = io_multiplicand[29] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1237 = io_multiplicand[30] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_1240 = io_multiplicand[31] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1249 = {_T_1240,_T_1237,_T_1234,_T_1231,_T_1228,_T_1225,_T_1222,_T_1219,_T_1216,_T_1213}; // @[Cat.scala 29:58]
  wire [18:0] _T_1258 = {_T_1249,_T_1210,_T_1207,_T_1204,_T_1201,_T_1198,_T_1195,_T_1192,_T_1189,_T_1186}; // @[Cat.scala 29:58]
  wire [27:0] _T_1267 = {_T_1258,_T_1183,_T_1180,_T_1177,_T_1174,_T_1171,_T_1168,_T_1165,_T_1162,_T_1159}; // @[Cat.scala 29:58]
  wire [30:0] _T_1270 = {_T_1267,_T_1156,_T_1153,_T_1150}; // @[Cat.scala 29:58]
  wire  _T_1306 = io_multiplicand[0] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1309 = io_multiplicand[1] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1312 = io_multiplicand[2] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1315 = io_multiplicand[3] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1318 = io_multiplicand[4] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1321 = io_multiplicand[5] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1324 = io_multiplicand[6] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1327 = io_multiplicand[7] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1330 = io_multiplicand[8] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1333 = io_multiplicand[9] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1336 = io_multiplicand[10] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1339 = io_multiplicand[11] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1342 = io_multiplicand[12] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1345 = io_multiplicand[13] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1348 = io_multiplicand[14] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1351 = io_multiplicand[15] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1354 = io_multiplicand[16] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1357 = io_multiplicand[17] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1360 = io_multiplicand[18] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1363 = io_multiplicand[19] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1366 = io_multiplicand[20] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1369 = io_multiplicand[21] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1372 = io_multiplicand[22] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1375 = io_multiplicand[23] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1378 = io_multiplicand[24] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1381 = io_multiplicand[25] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1384 = io_multiplicand[26] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1387 = io_multiplicand[27] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1390 = io_multiplicand[28] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1393 = io_multiplicand[29] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1396 = io_multiplicand[30] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_1399 = io_multiplicand[31] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1408 = {_T_1399,_T_1396,_T_1393,_T_1390,_T_1387,_T_1384,_T_1381,_T_1378,_T_1375,_T_1372}; // @[Cat.scala 29:58]
  wire [18:0] _T_1417 = {_T_1408,_T_1369,_T_1366,_T_1363,_T_1360,_T_1357,_T_1354,_T_1351,_T_1348,_T_1345}; // @[Cat.scala 29:58]
  wire [27:0] _T_1426 = {_T_1417,_T_1342,_T_1339,_T_1336,_T_1333,_T_1330,_T_1327,_T_1324,_T_1321,_T_1318}; // @[Cat.scala 29:58]
  wire [30:0] _T_1429 = {_T_1426,_T_1315,_T_1312,_T_1309}; // @[Cat.scala 29:58]
  wire  _T_1465 = io_multiplicand[0] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1468 = io_multiplicand[1] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1471 = io_multiplicand[2] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1474 = io_multiplicand[3] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1477 = io_multiplicand[4] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1480 = io_multiplicand[5] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1483 = io_multiplicand[6] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1486 = io_multiplicand[7] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1489 = io_multiplicand[8] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1492 = io_multiplicand[9] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1495 = io_multiplicand[10] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1498 = io_multiplicand[11] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1501 = io_multiplicand[12] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1504 = io_multiplicand[13] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1507 = io_multiplicand[14] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1510 = io_multiplicand[15] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1513 = io_multiplicand[16] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1516 = io_multiplicand[17] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1519 = io_multiplicand[18] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1522 = io_multiplicand[19] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1525 = io_multiplicand[20] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1528 = io_multiplicand[21] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1531 = io_multiplicand[22] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1534 = io_multiplicand[23] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1537 = io_multiplicand[24] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1540 = io_multiplicand[25] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1543 = io_multiplicand[26] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1546 = io_multiplicand[27] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1549 = io_multiplicand[28] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1552 = io_multiplicand[29] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1555 = io_multiplicand[30] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_1558 = io_multiplicand[31] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1567 = {_T_1558,_T_1555,_T_1552,_T_1549,_T_1546,_T_1543,_T_1540,_T_1537,_T_1534,_T_1531}; // @[Cat.scala 29:58]
  wire [18:0] _T_1576 = {_T_1567,_T_1528,_T_1525,_T_1522,_T_1519,_T_1516,_T_1513,_T_1510,_T_1507,_T_1504}; // @[Cat.scala 29:58]
  wire [27:0] _T_1585 = {_T_1576,_T_1501,_T_1498,_T_1495,_T_1492,_T_1489,_T_1486,_T_1483,_T_1480,_T_1477}; // @[Cat.scala 29:58]
  wire [30:0] _T_1588 = {_T_1585,_T_1474,_T_1471,_T_1468}; // @[Cat.scala 29:58]
  wire  _T_1624 = io_multiplicand[0] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1627 = io_multiplicand[1] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1630 = io_multiplicand[2] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1633 = io_multiplicand[3] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1636 = io_multiplicand[4] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1639 = io_multiplicand[5] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1642 = io_multiplicand[6] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1645 = io_multiplicand[7] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1648 = io_multiplicand[8] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1651 = io_multiplicand[9] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1654 = io_multiplicand[10] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1657 = io_multiplicand[11] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1660 = io_multiplicand[12] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1663 = io_multiplicand[13] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1666 = io_multiplicand[14] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1669 = io_multiplicand[15] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1672 = io_multiplicand[16] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1675 = io_multiplicand[17] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1678 = io_multiplicand[18] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1681 = io_multiplicand[19] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1684 = io_multiplicand[20] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1687 = io_multiplicand[21] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1690 = io_multiplicand[22] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1693 = io_multiplicand[23] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1696 = io_multiplicand[24] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1699 = io_multiplicand[25] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1702 = io_multiplicand[26] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1705 = io_multiplicand[27] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1708 = io_multiplicand[28] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1711 = io_multiplicand[29] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1714 = io_multiplicand[30] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_1717 = io_multiplicand[31] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1726 = {_T_1717,_T_1714,_T_1711,_T_1708,_T_1705,_T_1702,_T_1699,_T_1696,_T_1693,_T_1690}; // @[Cat.scala 29:58]
  wire [18:0] _T_1735 = {_T_1726,_T_1687,_T_1684,_T_1681,_T_1678,_T_1675,_T_1672,_T_1669,_T_1666,_T_1663}; // @[Cat.scala 29:58]
  wire [27:0] _T_1744 = {_T_1735,_T_1660,_T_1657,_T_1654,_T_1651,_T_1648,_T_1645,_T_1642,_T_1639,_T_1636}; // @[Cat.scala 29:58]
  wire [30:0] _T_1747 = {_T_1744,_T_1633,_T_1630,_T_1627}; // @[Cat.scala 29:58]
  wire  _T_1783 = io_multiplicand[0] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1786 = io_multiplicand[1] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1789 = io_multiplicand[2] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1792 = io_multiplicand[3] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1795 = io_multiplicand[4] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1798 = io_multiplicand[5] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1801 = io_multiplicand[6] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1804 = io_multiplicand[7] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1807 = io_multiplicand[8] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1810 = io_multiplicand[9] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1813 = io_multiplicand[10] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1816 = io_multiplicand[11] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1819 = io_multiplicand[12] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1822 = io_multiplicand[13] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1825 = io_multiplicand[14] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1828 = io_multiplicand[15] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1831 = io_multiplicand[16] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1834 = io_multiplicand[17] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1837 = io_multiplicand[18] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1840 = io_multiplicand[19] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1843 = io_multiplicand[20] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1846 = io_multiplicand[21] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1849 = io_multiplicand[22] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1852 = io_multiplicand[23] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1855 = io_multiplicand[24] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1858 = io_multiplicand[25] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1861 = io_multiplicand[26] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1864 = io_multiplicand[27] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1867 = io_multiplicand[28] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1870 = io_multiplicand[29] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1873 = io_multiplicand[30] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_1876 = io_multiplicand[31] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1885 = {_T_1876,_T_1873,_T_1870,_T_1867,_T_1864,_T_1861,_T_1858,_T_1855,_T_1852,_T_1849}; // @[Cat.scala 29:58]
  wire [18:0] _T_1894 = {_T_1885,_T_1846,_T_1843,_T_1840,_T_1837,_T_1834,_T_1831,_T_1828,_T_1825,_T_1822}; // @[Cat.scala 29:58]
  wire [27:0] _T_1903 = {_T_1894,_T_1819,_T_1816,_T_1813,_T_1810,_T_1807,_T_1804,_T_1801,_T_1798,_T_1795}; // @[Cat.scala 29:58]
  wire [30:0] _T_1906 = {_T_1903,_T_1792,_T_1789,_T_1786}; // @[Cat.scala 29:58]
  wire  _T_1942 = io_multiplicand[0] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1945 = io_multiplicand[1] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1948 = io_multiplicand[2] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1951 = io_multiplicand[3] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1954 = io_multiplicand[4] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1957 = io_multiplicand[5] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1960 = io_multiplicand[6] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1963 = io_multiplicand[7] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1966 = io_multiplicand[8] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1969 = io_multiplicand[9] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1972 = io_multiplicand[10] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1975 = io_multiplicand[11] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1978 = io_multiplicand[12] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1981 = io_multiplicand[13] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1984 = io_multiplicand[14] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1987 = io_multiplicand[15] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1990 = io_multiplicand[16] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1993 = io_multiplicand[17] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1996 = io_multiplicand[18] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1999 = io_multiplicand[19] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_2002 = io_multiplicand[20] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_2005 = io_multiplicand[21] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_2008 = io_multiplicand[22] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_2011 = io_multiplicand[23] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_2014 = io_multiplicand[24] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_2017 = io_multiplicand[25] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_2020 = io_multiplicand[26] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_2023 = io_multiplicand[27] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_2026 = io_multiplicand[28] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_2029 = io_multiplicand[29] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_2032 = io_multiplicand[30] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_2035 = io_multiplicand[31] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire [9:0] _T_2044 = {_T_2035,_T_2032,_T_2029,_T_2026,_T_2023,_T_2020,_T_2017,_T_2014,_T_2011,_T_2008}; // @[Cat.scala 29:58]
  wire [18:0] _T_2053 = {_T_2044,_T_2005,_T_2002,_T_1999,_T_1996,_T_1993,_T_1990,_T_1987,_T_1984,_T_1981}; // @[Cat.scala 29:58]
  wire [27:0] _T_2062 = {_T_2053,_T_1978,_T_1975,_T_1972,_T_1969,_T_1966,_T_1963,_T_1960,_T_1957,_T_1954}; // @[Cat.scala 29:58]
  wire [30:0] _T_2065 = {_T_2062,_T_1951,_T_1948,_T_1945}; // @[Cat.scala 29:58]
  wire  _T_2101 = io_multiplicand[0] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2104 = io_multiplicand[1] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2107 = io_multiplicand[2] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2110 = io_multiplicand[3] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2113 = io_multiplicand[4] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2116 = io_multiplicand[5] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2119 = io_multiplicand[6] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2122 = io_multiplicand[7] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2125 = io_multiplicand[8] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2128 = io_multiplicand[9] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2131 = io_multiplicand[10] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2134 = io_multiplicand[11] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2137 = io_multiplicand[12] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2140 = io_multiplicand[13] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2143 = io_multiplicand[14] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2146 = io_multiplicand[15] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2149 = io_multiplicand[16] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2152 = io_multiplicand[17] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2155 = io_multiplicand[18] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2158 = io_multiplicand[19] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2161 = io_multiplicand[20] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2164 = io_multiplicand[21] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2167 = io_multiplicand[22] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2170 = io_multiplicand[23] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2173 = io_multiplicand[24] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2176 = io_multiplicand[25] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2179 = io_multiplicand[26] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2182 = io_multiplicand[27] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2185 = io_multiplicand[28] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2188 = io_multiplicand[29] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2191 = io_multiplicand[30] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_2194 = io_multiplicand[31] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire [9:0] _T_2203 = {_T_2194,_T_2191,_T_2188,_T_2185,_T_2182,_T_2179,_T_2176,_T_2173,_T_2170,_T_2167}; // @[Cat.scala 29:58]
  wire [18:0] _T_2212 = {_T_2203,_T_2164,_T_2161,_T_2158,_T_2155,_T_2152,_T_2149,_T_2146,_T_2143,_T_2140}; // @[Cat.scala 29:58]
  wire [27:0] _T_2221 = {_T_2212,_T_2137,_T_2134,_T_2131,_T_2128,_T_2125,_T_2122,_T_2119,_T_2116,_T_2113}; // @[Cat.scala 29:58]
  wire [30:0] _T_2224 = {_T_2221,_T_2110,_T_2107,_T_2104}; // @[Cat.scala 29:58]
  wire  _T_2260 = io_multiplicand[0] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2263 = io_multiplicand[1] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2266 = io_multiplicand[2] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2269 = io_multiplicand[3] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2272 = io_multiplicand[4] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2275 = io_multiplicand[5] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2278 = io_multiplicand[6] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2281 = io_multiplicand[7] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2284 = io_multiplicand[8] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2287 = io_multiplicand[9] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2290 = io_multiplicand[10] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2293 = io_multiplicand[11] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2296 = io_multiplicand[12] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2299 = io_multiplicand[13] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2302 = io_multiplicand[14] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2305 = io_multiplicand[15] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2308 = io_multiplicand[16] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2311 = io_multiplicand[17] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2314 = io_multiplicand[18] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2317 = io_multiplicand[19] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2320 = io_multiplicand[20] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2323 = io_multiplicand[21] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2326 = io_multiplicand[22] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2329 = io_multiplicand[23] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2332 = io_multiplicand[24] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2335 = io_multiplicand[25] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2338 = io_multiplicand[26] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2341 = io_multiplicand[27] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2344 = io_multiplicand[28] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2347 = io_multiplicand[29] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2350 = io_multiplicand[30] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_2353 = io_multiplicand[31] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire [9:0] _T_2362 = {_T_2353,_T_2350,_T_2347,_T_2344,_T_2341,_T_2338,_T_2335,_T_2332,_T_2329,_T_2326}; // @[Cat.scala 29:58]
  wire [18:0] _T_2371 = {_T_2362,_T_2323,_T_2320,_T_2317,_T_2314,_T_2311,_T_2308,_T_2305,_T_2302,_T_2299}; // @[Cat.scala 29:58]
  wire [27:0] _T_2380 = {_T_2371,_T_2296,_T_2293,_T_2290,_T_2287,_T_2284,_T_2281,_T_2278,_T_2275,_T_2272}; // @[Cat.scala 29:58]
  wire [30:0] _T_2383 = {_T_2380,_T_2269,_T_2266,_T_2263}; // @[Cat.scala 29:58]
  wire  _T_2419 = io_multiplicand[0] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2422 = io_multiplicand[1] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2425 = io_multiplicand[2] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2428 = io_multiplicand[3] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2431 = io_multiplicand[4] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2434 = io_multiplicand[5] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2437 = io_multiplicand[6] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2440 = io_multiplicand[7] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2443 = io_multiplicand[8] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2446 = io_multiplicand[9] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2449 = io_multiplicand[10] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2452 = io_multiplicand[11] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2455 = io_multiplicand[12] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2458 = io_multiplicand[13] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2461 = io_multiplicand[14] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2464 = io_multiplicand[15] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2467 = io_multiplicand[16] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2470 = io_multiplicand[17] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2473 = io_multiplicand[18] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2476 = io_multiplicand[19] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2479 = io_multiplicand[20] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2482 = io_multiplicand[21] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2485 = io_multiplicand[22] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2488 = io_multiplicand[23] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2491 = io_multiplicand[24] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2494 = io_multiplicand[25] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2497 = io_multiplicand[26] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2500 = io_multiplicand[27] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2503 = io_multiplicand[28] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2506 = io_multiplicand[29] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2509 = io_multiplicand[30] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_2512 = io_multiplicand[31] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire [9:0] _T_2521 = {_T_2512,_T_2509,_T_2506,_T_2503,_T_2500,_T_2497,_T_2494,_T_2491,_T_2488,_T_2485}; // @[Cat.scala 29:58]
  wire [18:0] _T_2530 = {_T_2521,_T_2482,_T_2479,_T_2476,_T_2473,_T_2470,_T_2467,_T_2464,_T_2461,_T_2458}; // @[Cat.scala 29:58]
  wire [27:0] _T_2539 = {_T_2530,_T_2455,_T_2452,_T_2449,_T_2446,_T_2443,_T_2440,_T_2437,_T_2434,_T_2431}; // @[Cat.scala 29:58]
  wire [30:0] _T_2542 = {_T_2539,_T_2428,_T_2425,_T_2422}; // @[Cat.scala 29:58]
  wire  _T_2578 = io_multiplicand[0] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2581 = io_multiplicand[1] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2584 = io_multiplicand[2] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2587 = io_multiplicand[3] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2590 = io_multiplicand[4] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2593 = io_multiplicand[5] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2596 = io_multiplicand[6] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2599 = io_multiplicand[7] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2602 = io_multiplicand[8] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2605 = io_multiplicand[9] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2608 = io_multiplicand[10] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2611 = io_multiplicand[11] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2614 = io_multiplicand[12] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2617 = io_multiplicand[13] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2620 = io_multiplicand[14] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2623 = io_multiplicand[15] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2626 = io_multiplicand[16] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2629 = io_multiplicand[17] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2632 = io_multiplicand[18] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2635 = io_multiplicand[19] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2638 = io_multiplicand[20] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2641 = io_multiplicand[21] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2644 = io_multiplicand[22] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2647 = io_multiplicand[23] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2650 = io_multiplicand[24] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2653 = io_multiplicand[25] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2656 = io_multiplicand[26] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2659 = io_multiplicand[27] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2662 = io_multiplicand[28] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2665 = io_multiplicand[29] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2668 = io_multiplicand[30] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_2671 = io_multiplicand[31] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire [9:0] _T_2680 = {_T_2671,_T_2668,_T_2665,_T_2662,_T_2659,_T_2656,_T_2653,_T_2650,_T_2647,_T_2644}; // @[Cat.scala 29:58]
  wire [18:0] _T_2689 = {_T_2680,_T_2641,_T_2638,_T_2635,_T_2632,_T_2629,_T_2626,_T_2623,_T_2620,_T_2617}; // @[Cat.scala 29:58]
  wire [27:0] _T_2698 = {_T_2689,_T_2614,_T_2611,_T_2608,_T_2605,_T_2602,_T_2599,_T_2596,_T_2593,_T_2590}; // @[Cat.scala 29:58]
  wire [30:0] _T_2701 = {_T_2698,_T_2587,_T_2584,_T_2581}; // @[Cat.scala 29:58]
  wire  _T_2737 = io_multiplicand[0] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2740 = io_multiplicand[1] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2743 = io_multiplicand[2] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2746 = io_multiplicand[3] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2749 = io_multiplicand[4] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2752 = io_multiplicand[5] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2755 = io_multiplicand[6] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2758 = io_multiplicand[7] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2761 = io_multiplicand[8] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2764 = io_multiplicand[9] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2767 = io_multiplicand[10] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2770 = io_multiplicand[11] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2773 = io_multiplicand[12] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2776 = io_multiplicand[13] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2779 = io_multiplicand[14] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2782 = io_multiplicand[15] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2785 = io_multiplicand[16] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2788 = io_multiplicand[17] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2791 = io_multiplicand[18] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2794 = io_multiplicand[19] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2797 = io_multiplicand[20] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2800 = io_multiplicand[21] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2803 = io_multiplicand[22] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2806 = io_multiplicand[23] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2809 = io_multiplicand[24] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2812 = io_multiplicand[25] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2815 = io_multiplicand[26] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2818 = io_multiplicand[27] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2821 = io_multiplicand[28] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2824 = io_multiplicand[29] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2827 = io_multiplicand[30] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_2830 = io_multiplicand[31] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire [9:0] _T_2839 = {_T_2830,_T_2827,_T_2824,_T_2821,_T_2818,_T_2815,_T_2812,_T_2809,_T_2806,_T_2803}; // @[Cat.scala 29:58]
  wire [18:0] _T_2848 = {_T_2839,_T_2800,_T_2797,_T_2794,_T_2791,_T_2788,_T_2785,_T_2782,_T_2779,_T_2776}; // @[Cat.scala 29:58]
  wire [27:0] _T_2857 = {_T_2848,_T_2773,_T_2770,_T_2767,_T_2764,_T_2761,_T_2758,_T_2755,_T_2752,_T_2749}; // @[Cat.scala 29:58]
  wire [30:0] _T_2860 = {_T_2857,_T_2746,_T_2743,_T_2740}; // @[Cat.scala 29:58]
  wire  _T_2896 = io_multiplicand[0] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2899 = io_multiplicand[1] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2902 = io_multiplicand[2] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2905 = io_multiplicand[3] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2908 = io_multiplicand[4] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2911 = io_multiplicand[5] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2914 = io_multiplicand[6] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2917 = io_multiplicand[7] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2920 = io_multiplicand[8] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2923 = io_multiplicand[9] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2926 = io_multiplicand[10] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2929 = io_multiplicand[11] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2932 = io_multiplicand[12] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2935 = io_multiplicand[13] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2938 = io_multiplicand[14] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2941 = io_multiplicand[15] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2944 = io_multiplicand[16] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2947 = io_multiplicand[17] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2950 = io_multiplicand[18] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2953 = io_multiplicand[19] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2956 = io_multiplicand[20] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2959 = io_multiplicand[21] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2962 = io_multiplicand[22] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2965 = io_multiplicand[23] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2968 = io_multiplicand[24] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2971 = io_multiplicand[25] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2974 = io_multiplicand[26] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2977 = io_multiplicand[27] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2980 = io_multiplicand[28] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2983 = io_multiplicand[29] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2986 = io_multiplicand[30] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_2989 = io_multiplicand[31] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire [9:0] _T_2998 = {_T_2989,_T_2986,_T_2983,_T_2980,_T_2977,_T_2974,_T_2971,_T_2968,_T_2965,_T_2962}; // @[Cat.scala 29:58]
  wire [18:0] _T_3007 = {_T_2998,_T_2959,_T_2956,_T_2953,_T_2950,_T_2947,_T_2944,_T_2941,_T_2938,_T_2935}; // @[Cat.scala 29:58]
  wire [27:0] _T_3016 = {_T_3007,_T_2932,_T_2929,_T_2926,_T_2923,_T_2920,_T_2917,_T_2914,_T_2911,_T_2908}; // @[Cat.scala 29:58]
  wire [30:0] _T_3019 = {_T_3016,_T_2905,_T_2902,_T_2899}; // @[Cat.scala 29:58]
  wire  _T_3055 = io_multiplicand[0] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3058 = io_multiplicand[1] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3061 = io_multiplicand[2] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3064 = io_multiplicand[3] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3067 = io_multiplicand[4] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3070 = io_multiplicand[5] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3073 = io_multiplicand[6] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3076 = io_multiplicand[7] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3079 = io_multiplicand[8] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3082 = io_multiplicand[9] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3085 = io_multiplicand[10] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3088 = io_multiplicand[11] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3091 = io_multiplicand[12] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3094 = io_multiplicand[13] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3097 = io_multiplicand[14] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3100 = io_multiplicand[15] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3103 = io_multiplicand[16] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3106 = io_multiplicand[17] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3109 = io_multiplicand[18] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3112 = io_multiplicand[19] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3115 = io_multiplicand[20] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3118 = io_multiplicand[21] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3121 = io_multiplicand[22] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3124 = io_multiplicand[23] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3127 = io_multiplicand[24] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3130 = io_multiplicand[25] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3133 = io_multiplicand[26] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3136 = io_multiplicand[27] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3139 = io_multiplicand[28] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3142 = io_multiplicand[29] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3145 = io_multiplicand[30] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_3148 = io_multiplicand[31] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire [9:0] _T_3157 = {_T_3148,_T_3145,_T_3142,_T_3139,_T_3136,_T_3133,_T_3130,_T_3127,_T_3124,_T_3121}; // @[Cat.scala 29:58]
  wire [18:0] _T_3166 = {_T_3157,_T_3118,_T_3115,_T_3112,_T_3109,_T_3106,_T_3103,_T_3100,_T_3097,_T_3094}; // @[Cat.scala 29:58]
  wire [27:0] _T_3175 = {_T_3166,_T_3091,_T_3088,_T_3085,_T_3082,_T_3079,_T_3076,_T_3073,_T_3070,_T_3067}; // @[Cat.scala 29:58]
  wire [30:0] _T_3178 = {_T_3175,_T_3064,_T_3061,_T_3058}; // @[Cat.scala 29:58]
  wire  _T_3214 = io_multiplicand[0] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3217 = io_multiplicand[1] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3220 = io_multiplicand[2] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3223 = io_multiplicand[3] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3226 = io_multiplicand[4] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3229 = io_multiplicand[5] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3232 = io_multiplicand[6] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3235 = io_multiplicand[7] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3238 = io_multiplicand[8] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3241 = io_multiplicand[9] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3244 = io_multiplicand[10] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3247 = io_multiplicand[11] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3250 = io_multiplicand[12] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3253 = io_multiplicand[13] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3256 = io_multiplicand[14] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3259 = io_multiplicand[15] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3262 = io_multiplicand[16] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3265 = io_multiplicand[17] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3268 = io_multiplicand[18] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3271 = io_multiplicand[19] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3274 = io_multiplicand[20] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3277 = io_multiplicand[21] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3280 = io_multiplicand[22] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3283 = io_multiplicand[23] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3286 = io_multiplicand[24] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3289 = io_multiplicand[25] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3292 = io_multiplicand[26] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3295 = io_multiplicand[27] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3298 = io_multiplicand[28] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3301 = io_multiplicand[29] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3304 = io_multiplicand[30] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_3307 = io_multiplicand[31] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire [9:0] _T_3316 = {_T_3307,_T_3304,_T_3301,_T_3298,_T_3295,_T_3292,_T_3289,_T_3286,_T_3283,_T_3280}; // @[Cat.scala 29:58]
  wire [18:0] _T_3325 = {_T_3316,_T_3277,_T_3274,_T_3271,_T_3268,_T_3265,_T_3262,_T_3259,_T_3256,_T_3253}; // @[Cat.scala 29:58]
  wire [27:0] _T_3334 = {_T_3325,_T_3250,_T_3247,_T_3244,_T_3241,_T_3238,_T_3235,_T_3232,_T_3229,_T_3226}; // @[Cat.scala 29:58]
  wire [30:0] _T_3337 = {_T_3334,_T_3223,_T_3220,_T_3217}; // @[Cat.scala 29:58]
  wire  _T_3373 = io_multiplicand[0] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3376 = io_multiplicand[1] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3379 = io_multiplicand[2] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3382 = io_multiplicand[3] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3385 = io_multiplicand[4] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3388 = io_multiplicand[5] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3391 = io_multiplicand[6] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3394 = io_multiplicand[7] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3397 = io_multiplicand[8] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3400 = io_multiplicand[9] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3403 = io_multiplicand[10] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3406 = io_multiplicand[11] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3409 = io_multiplicand[12] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3412 = io_multiplicand[13] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3415 = io_multiplicand[14] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3418 = io_multiplicand[15] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3421 = io_multiplicand[16] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3424 = io_multiplicand[17] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3427 = io_multiplicand[18] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3430 = io_multiplicand[19] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3433 = io_multiplicand[20] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3436 = io_multiplicand[21] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3439 = io_multiplicand[22] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3442 = io_multiplicand[23] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3445 = io_multiplicand[24] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3448 = io_multiplicand[25] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3451 = io_multiplicand[26] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3454 = io_multiplicand[27] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3457 = io_multiplicand[28] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3460 = io_multiplicand[29] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3463 = io_multiplicand[30] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_3466 = io_multiplicand[31] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire [9:0] _T_3475 = {_T_3466,_T_3463,_T_3460,_T_3457,_T_3454,_T_3451,_T_3448,_T_3445,_T_3442,_T_3439}; // @[Cat.scala 29:58]
  wire [18:0] _T_3484 = {_T_3475,_T_3436,_T_3433,_T_3430,_T_3427,_T_3424,_T_3421,_T_3418,_T_3415,_T_3412}; // @[Cat.scala 29:58]
  wire [27:0] _T_3493 = {_T_3484,_T_3409,_T_3406,_T_3403,_T_3400,_T_3397,_T_3394,_T_3391,_T_3388,_T_3385}; // @[Cat.scala 29:58]
  wire [30:0] _T_3496 = {_T_3493,_T_3382,_T_3379,_T_3376}; // @[Cat.scala 29:58]
  wire  _T_3532 = io_multiplicand[0] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3535 = io_multiplicand[1] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3538 = io_multiplicand[2] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3541 = io_multiplicand[3] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3544 = io_multiplicand[4] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3547 = io_multiplicand[5] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3550 = io_multiplicand[6] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3553 = io_multiplicand[7] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3556 = io_multiplicand[8] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3559 = io_multiplicand[9] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3562 = io_multiplicand[10] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3565 = io_multiplicand[11] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3568 = io_multiplicand[12] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3571 = io_multiplicand[13] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3574 = io_multiplicand[14] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3577 = io_multiplicand[15] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3580 = io_multiplicand[16] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3583 = io_multiplicand[17] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3586 = io_multiplicand[18] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3589 = io_multiplicand[19] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3592 = io_multiplicand[20] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3595 = io_multiplicand[21] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3598 = io_multiplicand[22] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3601 = io_multiplicand[23] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3604 = io_multiplicand[24] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3607 = io_multiplicand[25] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3610 = io_multiplicand[26] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3613 = io_multiplicand[27] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3616 = io_multiplicand[28] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3619 = io_multiplicand[29] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3622 = io_multiplicand[30] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_3625 = io_multiplicand[31] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire [9:0] _T_3634 = {_T_3625,_T_3622,_T_3619,_T_3616,_T_3613,_T_3610,_T_3607,_T_3604,_T_3601,_T_3598}; // @[Cat.scala 29:58]
  wire [18:0] _T_3643 = {_T_3634,_T_3595,_T_3592,_T_3589,_T_3586,_T_3583,_T_3580,_T_3577,_T_3574,_T_3571}; // @[Cat.scala 29:58]
  wire [27:0] _T_3652 = {_T_3643,_T_3568,_T_3565,_T_3562,_T_3559,_T_3556,_T_3553,_T_3550,_T_3547,_T_3544}; // @[Cat.scala 29:58]
  wire [30:0] _T_3655 = {_T_3652,_T_3541,_T_3538,_T_3535}; // @[Cat.scala 29:58]
  wire  _T_3691 = io_multiplicand[0] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3694 = io_multiplicand[1] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3697 = io_multiplicand[2] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3700 = io_multiplicand[3] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3703 = io_multiplicand[4] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3706 = io_multiplicand[5] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3709 = io_multiplicand[6] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3712 = io_multiplicand[7] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3715 = io_multiplicand[8] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3718 = io_multiplicand[9] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3721 = io_multiplicand[10] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3724 = io_multiplicand[11] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3727 = io_multiplicand[12] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3730 = io_multiplicand[13] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3733 = io_multiplicand[14] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3736 = io_multiplicand[15] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3739 = io_multiplicand[16] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3742 = io_multiplicand[17] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3745 = io_multiplicand[18] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3748 = io_multiplicand[19] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3751 = io_multiplicand[20] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3754 = io_multiplicand[21] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3757 = io_multiplicand[22] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3760 = io_multiplicand[23] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3763 = io_multiplicand[24] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3766 = io_multiplicand[25] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3769 = io_multiplicand[26] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3772 = io_multiplicand[27] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3775 = io_multiplicand[28] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3778 = io_multiplicand[29] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3781 = io_multiplicand[30] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_3784 = io_multiplicand[31] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire [9:0] _T_3793 = {_T_3784,_T_3781,_T_3778,_T_3775,_T_3772,_T_3769,_T_3766,_T_3763,_T_3760,_T_3757}; // @[Cat.scala 29:58]
  wire [18:0] _T_3802 = {_T_3793,_T_3754,_T_3751,_T_3748,_T_3745,_T_3742,_T_3739,_T_3736,_T_3733,_T_3730}; // @[Cat.scala 29:58]
  wire [27:0] _T_3811 = {_T_3802,_T_3727,_T_3724,_T_3721,_T_3718,_T_3715,_T_3712,_T_3709,_T_3706,_T_3703}; // @[Cat.scala 29:58]
  wire [30:0] _T_3814 = {_T_3811,_T_3700,_T_3697,_T_3694}; // @[Cat.scala 29:58]
  wire  _T_3850 = io_multiplicand[0] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3853 = io_multiplicand[1] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3856 = io_multiplicand[2] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3859 = io_multiplicand[3] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3862 = io_multiplicand[4] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3865 = io_multiplicand[5] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3868 = io_multiplicand[6] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3871 = io_multiplicand[7] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3874 = io_multiplicand[8] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3877 = io_multiplicand[9] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3880 = io_multiplicand[10] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3883 = io_multiplicand[11] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3886 = io_multiplicand[12] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3889 = io_multiplicand[13] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3892 = io_multiplicand[14] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3895 = io_multiplicand[15] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3898 = io_multiplicand[16] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3901 = io_multiplicand[17] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3904 = io_multiplicand[18] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3907 = io_multiplicand[19] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3910 = io_multiplicand[20] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3913 = io_multiplicand[21] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3916 = io_multiplicand[22] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3919 = io_multiplicand[23] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3922 = io_multiplicand[24] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3925 = io_multiplicand[25] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3928 = io_multiplicand[26] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3931 = io_multiplicand[27] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3934 = io_multiplicand[28] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3937 = io_multiplicand[29] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3940 = io_multiplicand[30] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_3943 = io_multiplicand[31] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire [9:0] _T_3952 = {_T_3943,_T_3940,_T_3937,_T_3934,_T_3931,_T_3928,_T_3925,_T_3922,_T_3919,_T_3916}; // @[Cat.scala 29:58]
  wire [18:0] _T_3961 = {_T_3952,_T_3913,_T_3910,_T_3907,_T_3904,_T_3901,_T_3898,_T_3895,_T_3892,_T_3889}; // @[Cat.scala 29:58]
  wire [27:0] _T_3970 = {_T_3961,_T_3886,_T_3883,_T_3880,_T_3877,_T_3874,_T_3871,_T_3868,_T_3865,_T_3862}; // @[Cat.scala 29:58]
  wire [30:0] _T_3973 = {_T_3970,_T_3859,_T_3856,_T_3853}; // @[Cat.scala 29:58]
  wire  _T_4009 = io_multiplicand[0] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4012 = io_multiplicand[1] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4015 = io_multiplicand[2] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4018 = io_multiplicand[3] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4021 = io_multiplicand[4] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4024 = io_multiplicand[5] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4027 = io_multiplicand[6] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4030 = io_multiplicand[7] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4033 = io_multiplicand[8] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4036 = io_multiplicand[9] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4039 = io_multiplicand[10] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4042 = io_multiplicand[11] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4045 = io_multiplicand[12] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4048 = io_multiplicand[13] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4051 = io_multiplicand[14] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4054 = io_multiplicand[15] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4057 = io_multiplicand[16] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4060 = io_multiplicand[17] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4063 = io_multiplicand[18] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4066 = io_multiplicand[19] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4069 = io_multiplicand[20] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4072 = io_multiplicand[21] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4075 = io_multiplicand[22] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4078 = io_multiplicand[23] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4081 = io_multiplicand[24] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4084 = io_multiplicand[25] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4087 = io_multiplicand[26] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4090 = io_multiplicand[27] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4093 = io_multiplicand[28] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4096 = io_multiplicand[29] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4099 = io_multiplicand[30] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_4102 = io_multiplicand[31] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire [9:0] _T_4111 = {_T_4102,_T_4099,_T_4096,_T_4093,_T_4090,_T_4087,_T_4084,_T_4081,_T_4078,_T_4075}; // @[Cat.scala 29:58]
  wire [18:0] _T_4120 = {_T_4111,_T_4072,_T_4069,_T_4066,_T_4063,_T_4060,_T_4057,_T_4054,_T_4051,_T_4048}; // @[Cat.scala 29:58]
  wire [27:0] _T_4129 = {_T_4120,_T_4045,_T_4042,_T_4039,_T_4036,_T_4033,_T_4030,_T_4027,_T_4024,_T_4021}; // @[Cat.scala 29:58]
  wire [30:0] _T_4132 = {_T_4129,_T_4018,_T_4015,_T_4012}; // @[Cat.scala 29:58]
  wire  _T_4168 = io_multiplicand[0] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4171 = io_multiplicand[1] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4174 = io_multiplicand[2] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4177 = io_multiplicand[3] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4180 = io_multiplicand[4] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4183 = io_multiplicand[5] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4186 = io_multiplicand[6] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4189 = io_multiplicand[7] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4192 = io_multiplicand[8] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4195 = io_multiplicand[9] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4198 = io_multiplicand[10] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4201 = io_multiplicand[11] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4204 = io_multiplicand[12] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4207 = io_multiplicand[13] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4210 = io_multiplicand[14] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4213 = io_multiplicand[15] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4216 = io_multiplicand[16] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4219 = io_multiplicand[17] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4222 = io_multiplicand[18] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4225 = io_multiplicand[19] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4228 = io_multiplicand[20] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4231 = io_multiplicand[21] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4234 = io_multiplicand[22] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4237 = io_multiplicand[23] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4240 = io_multiplicand[24] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4243 = io_multiplicand[25] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4246 = io_multiplicand[26] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4249 = io_multiplicand[27] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4252 = io_multiplicand[28] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4255 = io_multiplicand[29] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4258 = io_multiplicand[30] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_4261 = io_multiplicand[31] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire [9:0] _T_4270 = {_T_4261,_T_4258,_T_4255,_T_4252,_T_4249,_T_4246,_T_4243,_T_4240,_T_4237,_T_4234}; // @[Cat.scala 29:58]
  wire [18:0] _T_4279 = {_T_4270,_T_4231,_T_4228,_T_4225,_T_4222,_T_4219,_T_4216,_T_4213,_T_4210,_T_4207}; // @[Cat.scala 29:58]
  wire [27:0] _T_4288 = {_T_4279,_T_4204,_T_4201,_T_4198,_T_4195,_T_4192,_T_4189,_T_4186,_T_4183,_T_4180}; // @[Cat.scala 29:58]
  wire [30:0] _T_4291 = {_T_4288,_T_4177,_T_4174,_T_4171}; // @[Cat.scala 29:58]
  wire  _T_4327 = io_multiplicand[0] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4330 = io_multiplicand[1] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4333 = io_multiplicand[2] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4336 = io_multiplicand[3] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4339 = io_multiplicand[4] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4342 = io_multiplicand[5] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4345 = io_multiplicand[6] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4348 = io_multiplicand[7] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4351 = io_multiplicand[8] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4354 = io_multiplicand[9] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4357 = io_multiplicand[10] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4360 = io_multiplicand[11] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4363 = io_multiplicand[12] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4366 = io_multiplicand[13] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4369 = io_multiplicand[14] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4372 = io_multiplicand[15] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4375 = io_multiplicand[16] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4378 = io_multiplicand[17] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4381 = io_multiplicand[18] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4384 = io_multiplicand[19] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4387 = io_multiplicand[20] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4390 = io_multiplicand[21] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4393 = io_multiplicand[22] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4396 = io_multiplicand[23] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4399 = io_multiplicand[24] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4402 = io_multiplicand[25] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4405 = io_multiplicand[26] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4408 = io_multiplicand[27] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4411 = io_multiplicand[28] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4414 = io_multiplicand[29] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4417 = io_multiplicand[30] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_4420 = io_multiplicand[31] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire [9:0] _T_4429 = {_T_4420,_T_4417,_T_4414,_T_4411,_T_4408,_T_4405,_T_4402,_T_4399,_T_4396,_T_4393}; // @[Cat.scala 29:58]
  wire [18:0] _T_4438 = {_T_4429,_T_4390,_T_4387,_T_4384,_T_4381,_T_4378,_T_4375,_T_4372,_T_4369,_T_4366}; // @[Cat.scala 29:58]
  wire [27:0] _T_4447 = {_T_4438,_T_4363,_T_4360,_T_4357,_T_4354,_T_4351,_T_4348,_T_4345,_T_4342,_T_4339}; // @[Cat.scala 29:58]
  wire [30:0] _T_4450 = {_T_4447,_T_4336,_T_4333,_T_4330}; // @[Cat.scala 29:58]
  wire  _T_4486 = io_multiplicand[0] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4489 = io_multiplicand[1] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4492 = io_multiplicand[2] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4495 = io_multiplicand[3] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4498 = io_multiplicand[4] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4501 = io_multiplicand[5] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4504 = io_multiplicand[6] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4507 = io_multiplicand[7] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4510 = io_multiplicand[8] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4513 = io_multiplicand[9] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4516 = io_multiplicand[10] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4519 = io_multiplicand[11] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4522 = io_multiplicand[12] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4525 = io_multiplicand[13] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4528 = io_multiplicand[14] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4531 = io_multiplicand[15] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4534 = io_multiplicand[16] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4537 = io_multiplicand[17] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4540 = io_multiplicand[18] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4543 = io_multiplicand[19] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4546 = io_multiplicand[20] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4549 = io_multiplicand[21] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4552 = io_multiplicand[22] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4555 = io_multiplicand[23] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4558 = io_multiplicand[24] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4561 = io_multiplicand[25] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4564 = io_multiplicand[26] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4567 = io_multiplicand[27] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4570 = io_multiplicand[28] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4573 = io_multiplicand[29] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4576 = io_multiplicand[30] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_4579 = io_multiplicand[31] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire [9:0] _T_4588 = {_T_4579,_T_4576,_T_4573,_T_4570,_T_4567,_T_4564,_T_4561,_T_4558,_T_4555,_T_4552}; // @[Cat.scala 29:58]
  wire [18:0] _T_4597 = {_T_4588,_T_4549,_T_4546,_T_4543,_T_4540,_T_4537,_T_4534,_T_4531,_T_4528,_T_4525}; // @[Cat.scala 29:58]
  wire [27:0] _T_4606 = {_T_4597,_T_4522,_T_4519,_T_4516,_T_4513,_T_4510,_T_4507,_T_4504,_T_4501,_T_4498}; // @[Cat.scala 29:58]
  wire [30:0] _T_4609 = {_T_4606,_T_4495,_T_4492,_T_4489}; // @[Cat.scala 29:58]
  wire  _T_4645 = io_multiplicand[0] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4648 = io_multiplicand[1] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4651 = io_multiplicand[2] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4654 = io_multiplicand[3] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4657 = io_multiplicand[4] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4660 = io_multiplicand[5] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4663 = io_multiplicand[6] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4666 = io_multiplicand[7] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4669 = io_multiplicand[8] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4672 = io_multiplicand[9] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4675 = io_multiplicand[10] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4678 = io_multiplicand[11] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4681 = io_multiplicand[12] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4684 = io_multiplicand[13] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4687 = io_multiplicand[14] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4690 = io_multiplicand[15] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4693 = io_multiplicand[16] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4696 = io_multiplicand[17] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4699 = io_multiplicand[18] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4702 = io_multiplicand[19] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4705 = io_multiplicand[20] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4708 = io_multiplicand[21] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4711 = io_multiplicand[22] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4714 = io_multiplicand[23] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4717 = io_multiplicand[24] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4720 = io_multiplicand[25] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4723 = io_multiplicand[26] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4726 = io_multiplicand[27] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4729 = io_multiplicand[28] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4732 = io_multiplicand[29] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4735 = io_multiplicand[30] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_4738 = io_multiplicand[31] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire [9:0] _T_4747 = {_T_4738,_T_4735,_T_4732,_T_4729,_T_4726,_T_4723,_T_4720,_T_4717,_T_4714,_T_4711}; // @[Cat.scala 29:58]
  wire [18:0] _T_4756 = {_T_4747,_T_4708,_T_4705,_T_4702,_T_4699,_T_4696,_T_4693,_T_4690,_T_4687,_T_4684}; // @[Cat.scala 29:58]
  wire [27:0] _T_4765 = {_T_4756,_T_4681,_T_4678,_T_4675,_T_4672,_T_4669,_T_4666,_T_4663,_T_4660,_T_4657}; // @[Cat.scala 29:58]
  wire [30:0] _T_4768 = {_T_4765,_T_4654,_T_4651,_T_4648}; // @[Cat.scala 29:58]
  wire  _T_4804 = io_multiplicand[0] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4807 = io_multiplicand[1] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4810 = io_multiplicand[2] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4813 = io_multiplicand[3] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4816 = io_multiplicand[4] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4819 = io_multiplicand[5] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4822 = io_multiplicand[6] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4825 = io_multiplicand[7] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4828 = io_multiplicand[8] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4831 = io_multiplicand[9] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4834 = io_multiplicand[10] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4837 = io_multiplicand[11] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4840 = io_multiplicand[12] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4843 = io_multiplicand[13] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4846 = io_multiplicand[14] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4849 = io_multiplicand[15] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4852 = io_multiplicand[16] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4855 = io_multiplicand[17] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4858 = io_multiplicand[18] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4861 = io_multiplicand[19] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4864 = io_multiplicand[20] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4867 = io_multiplicand[21] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4870 = io_multiplicand[22] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4873 = io_multiplicand[23] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4876 = io_multiplicand[24] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4879 = io_multiplicand[25] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4882 = io_multiplicand[26] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4885 = io_multiplicand[27] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4888 = io_multiplicand[28] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4891 = io_multiplicand[29] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4894 = io_multiplicand[30] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_4897 = io_multiplicand[31] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire [9:0] _T_4906 = {_T_4897,_T_4894,_T_4891,_T_4888,_T_4885,_T_4882,_T_4879,_T_4876,_T_4873,_T_4870}; // @[Cat.scala 29:58]
  wire [18:0] _T_4915 = {_T_4906,_T_4867,_T_4864,_T_4861,_T_4858,_T_4855,_T_4852,_T_4849,_T_4846,_T_4843}; // @[Cat.scala 29:58]
  wire [27:0] _T_4924 = {_T_4915,_T_4840,_T_4837,_T_4834,_T_4831,_T_4828,_T_4825,_T_4822,_T_4819,_T_4816}; // @[Cat.scala 29:58]
  wire [30:0] _T_4927 = {_T_4924,_T_4813,_T_4810,_T_4807}; // @[Cat.scala 29:58]
  wire  _T_4963 = io_multiplicand[0] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_4966 = io_multiplicand[1] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_4969 = io_multiplicand[2] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_4972 = io_multiplicand[3] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_4975 = io_multiplicand[4] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_4978 = io_multiplicand[5] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_4981 = io_multiplicand[6] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_4984 = io_multiplicand[7] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_4987 = io_multiplicand[8] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_4990 = io_multiplicand[9] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_4993 = io_multiplicand[10] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_4996 = io_multiplicand[11] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_4999 = io_multiplicand[12] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5002 = io_multiplicand[13] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5005 = io_multiplicand[14] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5008 = io_multiplicand[15] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5011 = io_multiplicand[16] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5014 = io_multiplicand[17] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5017 = io_multiplicand[18] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5020 = io_multiplicand[19] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5023 = io_multiplicand[20] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5026 = io_multiplicand[21] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5029 = io_multiplicand[22] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5032 = io_multiplicand[23] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5035 = io_multiplicand[24] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5038 = io_multiplicand[25] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5041 = io_multiplicand[26] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5044 = io_multiplicand[27] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5047 = io_multiplicand[28] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5050 = io_multiplicand[29] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5053 = io_multiplicand[30] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_5056 = io_multiplicand[31] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire [9:0] _T_5065 = {_T_5056,_T_5053,_T_5050,_T_5047,_T_5044,_T_5041,_T_5038,_T_5035,_T_5032,_T_5029}; // @[Cat.scala 29:58]
  wire [18:0] _T_5074 = {_T_5065,_T_5026,_T_5023,_T_5020,_T_5017,_T_5014,_T_5011,_T_5008,_T_5005,_T_5002}; // @[Cat.scala 29:58]
  wire [27:0] _T_5083 = {_T_5074,_T_4999,_T_4996,_T_4993,_T_4990,_T_4987,_T_4984,_T_4981,_T_4978,_T_4975}; // @[Cat.scala 29:58]
  wire [30:0] _T_5086 = {_T_5083,_T_4972,_T_4969,_T_4966}; // @[Cat.scala 29:58]
  assign io_outs_0 = {_T_157,_T_34}; // @[partialprod.scala 18:16]
  assign io_outs_1 = {_T_316,_T_193}; // @[partialprod.scala 18:16]
  assign io_outs_2 = {_T_475,_T_352}; // @[partialprod.scala 18:16]
  assign io_outs_3 = {_T_634,_T_511}; // @[partialprod.scala 18:16]
  assign io_outs_4 = {_T_793,_T_670}; // @[partialprod.scala 18:16]
  assign io_outs_5 = {_T_952,_T_829}; // @[partialprod.scala 18:16]
  assign io_outs_6 = {_T_1111,_T_988}; // @[partialprod.scala 18:16]
  assign io_outs_7 = {_T_1270,_T_1147}; // @[partialprod.scala 18:16]
  assign io_outs_8 = {_T_1429,_T_1306}; // @[partialprod.scala 18:16]
  assign io_outs_9 = {_T_1588,_T_1465}; // @[partialprod.scala 18:16]
  assign io_outs_10 = {_T_1747,_T_1624}; // @[partialprod.scala 18:16]
  assign io_outs_11 = {_T_1906,_T_1783}; // @[partialprod.scala 18:16]
  assign io_outs_12 = {_T_2065,_T_1942}; // @[partialprod.scala 18:16]
  assign io_outs_13 = {_T_2224,_T_2101}; // @[partialprod.scala 18:16]
  assign io_outs_14 = {_T_2383,_T_2260}; // @[partialprod.scala 18:16]
  assign io_outs_15 = {_T_2542,_T_2419}; // @[partialprod.scala 18:16]
  assign io_outs_16 = {_T_2701,_T_2578}; // @[partialprod.scala 18:16]
  assign io_outs_17 = {_T_2860,_T_2737}; // @[partialprod.scala 18:16]
  assign io_outs_18 = {_T_3019,_T_2896}; // @[partialprod.scala 18:16]
  assign io_outs_19 = {_T_3178,_T_3055}; // @[partialprod.scala 18:16]
  assign io_outs_20 = {_T_3337,_T_3214}; // @[partialprod.scala 18:16]
  assign io_outs_21 = {_T_3496,_T_3373}; // @[partialprod.scala 18:16]
  assign io_outs_22 = {_T_3655,_T_3532}; // @[partialprod.scala 18:16]
  assign io_outs_23 = {_T_3814,_T_3691}; // @[partialprod.scala 18:16]
  assign io_outs_24 = {_T_3973,_T_3850}; // @[partialprod.scala 18:16]
  assign io_outs_25 = {_T_4132,_T_4009}; // @[partialprod.scala 18:16]
  assign io_outs_26 = {_T_4291,_T_4168}; // @[partialprod.scala 18:16]
  assign io_outs_27 = {_T_4450,_T_4327}; // @[partialprod.scala 18:16]
  assign io_outs_28 = {_T_4609,_T_4486}; // @[partialprod.scala 18:16]
  assign io_outs_29 = {_T_4768,_T_4645}; // @[partialprod.scala 18:16]
  assign io_outs_30 = {_T_4927,_T_4804}; // @[partialprod.scala 18:16]
  assign io_outs_31 = {_T_5086,_T_4963}; // @[partialprod.scala 18:16]
endmodule
module HalfAdder(
  input   io_a,
  input   io_b,
  output  io_s,
  output  io_co
);
  assign io_s = io_a ^ io_b; // @[comp.scala 15:8]
  assign io_co = io_a & io_b; // @[comp.scala 16:9]
endmodule
module FullAdder(
  input   io_a,
  input   io_b,
  input   io_ci,
  output  io_s,
  output  io_co
);
  wire  a_xor_b = io_a ^ io_b; // @[comp.scala 28:22]
  wire  a_and_b = io_a & io_b; // @[comp.scala 31:22]
  wire  a_and_cin = io_a & io_ci; // @[comp.scala 32:24]
  wire  b_and_cin = io_b & io_ci; // @[comp.scala 33:24]
  wire  _T_1 = a_and_b | b_and_cin; // @[comp.scala 34:20]
  assign io_s = a_xor_b ^ io_ci; // @[comp.scala 29:8]
  assign io_co = _T_1 | a_and_cin; // @[comp.scala 34:9]
endmodule
module Wallace(
  input  [31:0] io_pp_0,
  input  [31:0] io_pp_1,
  input  [31:0] io_pp_2,
  input  [31:0] io_pp_3,
  input  [31:0] io_pp_4,
  input  [31:0] io_pp_5,
  input  [31:0] io_pp_6,
  input  [31:0] io_pp_7,
  input  [31:0] io_pp_8,
  input  [31:0] io_pp_9,
  input  [31:0] io_pp_10,
  input  [31:0] io_pp_11,
  input  [31:0] io_pp_12,
  input  [31:0] io_pp_13,
  input  [31:0] io_pp_14,
  input  [31:0] io_pp_15,
  input  [31:0] io_pp_16,
  input  [31:0] io_pp_17,
  input  [31:0] io_pp_18,
  input  [31:0] io_pp_19,
  input  [31:0] io_pp_20,
  input  [31:0] io_pp_21,
  input  [31:0] io_pp_22,
  input  [31:0] io_pp_23,
  input  [31:0] io_pp_24,
  input  [31:0] io_pp_25,
  input  [31:0] io_pp_26,
  input  [31:0] io_pp_27,
  input  [31:0] io_pp_28,
  input  [31:0] io_pp_29,
  input  [31:0] io_pp_30,
  input  [31:0] io_pp_31,
  output [63:0] io_augend,
  output [63:0] io_addend
);
  wire  HalfAdder_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_1_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_1_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_1_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_1_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_2_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_2_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_2_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_2_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_4_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_4_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_4_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_4_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_4_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_5_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_5_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_5_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_5_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_5_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_6_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_6_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_6_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_6_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_6_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_7_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_7_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_7_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_7_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_7_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_8_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_8_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_8_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_8_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_8_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_9_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_9_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_9_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_9_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_9_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_10_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_10_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_10_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_10_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_10_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_11_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_11_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_11_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_11_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_11_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_12_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_12_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_12_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_12_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_12_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_13_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_13_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_13_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_13_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_13_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_14_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_14_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_14_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_14_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_14_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_15_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_15_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_15_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_15_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_15_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_16_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_16_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_16_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_16_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_16_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_3_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_3_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_3_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_3_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_17_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_17_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_17_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_17_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_17_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_18_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_18_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_18_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_18_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_18_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_19_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_19_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_19_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_19_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_19_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_20_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_20_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_20_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_20_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_20_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_21_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_21_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_21_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_21_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_21_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_22_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_22_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_22_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_22_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_22_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_23_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_23_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_23_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_23_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_23_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_24_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_24_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_24_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_24_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_24_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_25_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_25_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_25_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_25_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_25_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_26_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_26_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_26_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_26_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_26_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_27_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_27_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_27_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_27_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_27_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_28_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_28_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_28_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_28_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_28_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_4_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_4_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_4_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_4_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_29_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_29_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_29_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_29_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_29_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_30_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_30_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_30_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_30_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_30_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_31_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_31_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_31_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_31_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_31_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_32_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_32_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_32_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_32_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_32_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_33_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_33_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_33_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_33_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_33_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_34_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_34_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_34_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_34_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_34_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_35_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_35_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_35_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_35_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_35_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_36_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_36_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_36_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_36_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_36_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_37_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_37_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_37_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_37_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_37_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_38_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_38_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_38_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_38_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_38_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_39_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_39_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_39_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_39_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_39_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_40_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_40_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_40_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_40_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_40_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_41_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_41_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_41_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_41_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_41_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_42_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_42_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_42_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_42_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_42_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_43_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_43_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_43_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_43_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_43_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_5_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_5_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_5_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_5_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_44_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_44_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_44_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_44_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_44_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_45_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_45_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_45_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_45_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_45_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_46_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_46_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_46_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_46_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_46_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_47_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_47_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_47_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_47_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_47_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_48_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_48_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_48_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_48_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_48_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_49_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_49_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_49_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_49_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_49_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_50_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_50_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_50_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_50_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_50_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_51_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_51_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_51_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_51_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_51_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_52_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_52_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_52_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_52_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_52_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_53_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_53_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_53_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_53_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_53_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_54_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_54_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_54_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_54_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_54_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_55_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_55_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_55_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_55_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_55_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_56_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_56_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_56_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_56_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_56_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_57_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_57_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_57_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_57_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_57_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_58_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_58_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_58_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_58_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_58_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_59_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_59_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_59_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_59_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_59_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_60_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_60_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_60_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_60_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_60_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_61_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_61_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_61_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_61_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_61_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_62_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_62_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_62_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_62_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_62_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_63_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_63_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_63_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_63_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_63_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_64_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_64_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_64_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_64_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_64_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_65_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_65_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_65_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_65_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_65_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_66_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_66_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_66_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_66_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_66_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_67_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_67_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_67_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_67_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_67_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_68_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_68_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_68_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_68_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_68_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_69_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_69_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_69_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_69_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_69_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_70_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_70_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_70_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_70_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_70_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_71_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_71_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_71_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_71_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_71_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_72_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_72_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_72_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_72_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_72_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_73_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_73_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_73_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_73_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_73_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_74_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_74_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_74_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_74_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_74_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_75_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_75_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_75_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_75_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_75_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_76_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_76_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_76_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_76_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_76_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_77_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_77_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_77_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_77_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_77_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_78_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_78_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_78_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_78_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_78_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_79_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_79_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_79_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_79_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_79_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_80_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_80_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_80_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_80_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_80_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_81_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_81_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_81_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_81_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_81_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_82_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_82_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_82_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_82_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_82_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_6_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_6_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_6_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_6_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_83_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_83_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_83_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_83_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_83_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_84_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_84_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_84_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_84_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_84_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_85_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_85_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_85_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_85_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_85_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_86_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_86_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_86_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_86_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_86_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_87_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_87_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_87_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_87_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_87_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_88_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_88_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_88_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_88_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_88_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_89_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_89_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_89_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_89_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_89_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_90_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_90_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_90_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_90_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_90_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_91_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_91_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_91_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_91_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_91_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_92_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_92_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_92_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_92_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_92_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_93_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_93_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_93_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_93_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_93_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_94_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_94_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_94_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_94_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_94_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_95_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_95_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_95_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_95_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_95_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_96_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_96_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_96_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_96_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_96_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_97_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_97_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_97_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_97_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_97_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_98_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_98_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_98_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_98_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_98_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_99_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_99_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_99_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_99_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_99_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_100_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_100_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_100_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_100_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_100_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_101_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_101_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_101_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_101_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_101_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_102_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_102_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_102_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_102_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_102_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_103_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_103_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_103_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_103_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_103_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_104_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_104_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_104_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_104_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_104_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_105_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_105_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_105_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_105_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_105_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_106_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_106_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_106_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_106_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_106_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_107_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_107_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_107_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_107_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_107_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_108_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_108_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_108_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_108_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_108_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_109_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_109_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_109_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_109_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_109_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_110_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_110_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_110_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_110_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_110_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_111_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_111_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_111_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_111_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_111_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_112_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_112_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_112_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_112_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_112_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_113_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_113_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_113_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_113_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_113_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_114_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_114_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_114_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_114_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_114_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_115_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_115_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_115_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_115_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_115_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_116_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_116_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_116_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_116_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_116_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_117_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_117_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_117_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_117_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_117_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_118_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_118_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_118_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_118_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_118_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_119_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_119_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_119_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_119_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_119_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_120_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_120_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_120_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_120_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_120_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_121_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_121_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_121_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_121_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_121_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_122_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_122_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_122_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_122_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_122_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_123_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_123_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_123_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_123_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_123_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_124_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_124_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_124_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_124_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_124_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_125_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_125_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_125_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_125_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_125_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_126_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_126_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_126_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_126_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_126_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_127_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_127_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_127_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_127_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_127_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_128_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_128_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_128_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_128_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_128_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_129_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_129_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_129_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_129_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_129_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_130_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_130_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_130_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_130_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_130_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_131_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_131_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_131_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_131_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_131_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_132_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_132_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_132_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_132_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_132_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_133_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_133_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_133_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_133_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_133_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_7_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_7_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_7_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_7_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_134_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_134_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_134_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_134_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_134_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_135_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_135_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_135_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_135_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_135_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_136_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_136_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_136_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_136_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_136_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_137_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_137_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_137_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_137_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_137_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_138_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_138_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_138_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_138_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_138_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_139_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_139_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_139_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_139_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_139_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_140_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_140_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_140_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_140_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_140_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_141_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_141_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_141_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_141_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_141_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_142_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_142_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_142_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_142_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_142_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_143_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_143_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_143_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_143_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_143_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_144_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_144_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_144_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_144_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_144_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_145_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_145_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_145_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_145_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_145_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_146_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_146_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_146_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_146_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_146_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_147_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_147_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_147_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_147_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_147_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_148_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_148_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_148_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_148_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_148_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_149_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_149_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_149_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_149_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_149_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_150_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_150_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_150_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_150_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_150_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_151_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_151_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_151_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_151_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_151_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_152_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_152_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_152_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_152_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_152_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_153_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_153_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_153_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_153_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_153_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_154_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_154_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_154_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_154_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_154_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_155_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_155_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_155_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_155_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_155_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_156_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_156_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_156_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_156_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_156_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_157_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_157_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_157_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_157_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_157_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_158_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_158_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_158_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_158_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_158_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_159_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_159_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_159_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_159_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_159_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_160_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_160_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_160_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_160_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_160_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_161_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_161_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_161_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_161_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_161_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_162_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_162_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_162_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_162_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_162_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_163_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_163_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_163_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_163_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_163_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_164_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_164_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_164_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_164_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_164_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_165_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_165_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_165_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_165_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_165_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_166_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_166_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_166_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_166_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_166_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_167_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_167_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_167_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_167_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_167_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_168_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_168_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_168_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_168_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_168_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_169_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_169_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_169_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_169_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_169_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_170_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_170_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_170_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_170_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_170_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_171_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_171_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_171_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_171_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_171_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_172_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_172_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_172_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_172_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_172_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_173_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_173_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_173_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_173_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_173_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_174_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_174_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_174_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_174_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_174_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_175_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_175_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_175_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_175_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_175_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_176_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_176_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_176_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_176_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_176_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_177_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_177_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_177_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_177_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_177_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_178_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_178_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_178_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_178_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_178_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_179_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_179_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_179_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_179_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_179_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_180_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_180_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_180_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_180_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_180_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_181_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_181_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_181_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_181_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_181_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_182_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_182_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_182_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_182_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_182_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_183_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_183_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_183_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_183_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_183_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_184_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_184_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_184_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_184_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_184_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_185_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_185_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_185_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_185_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_185_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_186_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_186_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_186_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_186_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_186_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_187_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_187_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_187_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_187_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_187_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_188_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_188_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_188_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_188_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_188_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_189_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_189_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_189_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_189_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_189_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_190_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_190_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_190_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_190_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_190_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_191_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_191_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_191_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_191_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_191_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_192_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_192_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_192_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_192_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_192_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_8_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_8_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_8_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_8_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_193_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_193_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_193_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_193_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_193_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_194_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_194_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_194_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_194_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_194_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_195_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_195_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_195_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_195_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_195_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_196_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_196_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_196_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_196_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_196_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_197_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_197_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_197_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_197_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_197_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_198_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_198_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_198_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_198_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_198_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_199_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_199_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_199_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_199_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_199_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_200_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_200_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_200_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_200_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_200_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_201_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_201_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_201_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_201_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_201_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_202_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_202_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_202_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_202_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_202_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_203_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_203_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_203_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_203_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_203_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_204_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_204_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_204_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_204_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_204_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_205_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_205_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_205_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_205_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_205_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_206_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_206_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_206_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_206_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_206_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_207_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_207_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_207_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_207_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_207_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_208_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_208_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_208_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_208_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_208_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_209_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_209_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_209_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_209_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_209_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_210_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_210_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_210_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_210_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_210_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_211_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_211_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_211_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_211_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_211_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_212_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_212_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_212_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_212_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_212_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_213_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_213_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_213_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_213_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_213_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_214_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_214_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_214_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_214_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_214_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_215_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_215_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_215_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_215_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_215_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_216_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_216_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_216_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_216_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_216_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_217_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_217_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_217_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_217_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_217_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_218_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_218_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_218_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_218_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_218_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_9_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_9_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_9_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_9_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_219_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_219_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_219_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_219_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_219_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_220_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_220_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_220_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_220_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_220_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_221_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_221_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_221_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_221_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_221_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_222_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_222_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_222_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_222_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_222_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_223_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_223_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_223_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_223_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_223_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_224_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_224_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_224_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_224_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_224_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_225_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_225_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_225_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_225_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_225_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_226_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_226_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_226_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_226_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_226_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_227_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_227_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_227_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_227_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_227_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_228_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_228_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_228_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_228_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_228_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_229_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_229_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_229_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_229_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_229_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_230_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_230_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_230_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_230_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_230_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_231_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_231_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_231_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_231_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_231_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_232_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_232_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_232_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_232_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_232_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_233_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_233_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_233_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_233_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_233_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_234_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_234_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_234_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_234_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_234_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_235_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_235_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_235_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_235_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_235_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_236_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_236_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_236_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_236_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_236_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_237_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_237_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_237_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_237_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_237_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_238_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_238_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_238_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_238_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_238_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_239_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_239_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_239_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_239_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_239_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_240_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_240_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_240_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_240_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_240_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_241_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_241_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_241_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_241_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_241_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_242_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_242_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_242_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_242_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_242_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_243_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_243_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_243_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_243_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_243_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_244_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_244_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_244_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_244_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_244_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_245_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_245_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_245_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_245_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_245_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_246_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_246_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_246_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_246_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_246_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_247_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_247_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_247_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_247_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_247_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_248_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_248_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_248_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_248_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_248_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_249_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_249_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_249_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_249_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_249_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_250_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_250_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_250_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_250_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_250_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_251_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_251_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_251_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_251_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_251_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_252_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_252_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_252_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_252_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_252_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_253_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_253_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_253_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_253_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_253_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_254_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_254_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_254_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_254_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_254_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_255_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_255_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_255_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_255_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_255_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_256_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_256_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_256_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_256_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_256_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_257_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_257_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_257_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_257_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_257_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_258_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_258_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_258_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_258_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_258_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_259_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_259_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_259_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_259_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_259_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_260_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_260_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_260_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_260_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_260_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_261_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_261_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_261_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_261_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_261_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_262_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_262_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_262_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_262_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_262_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_263_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_263_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_263_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_263_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_263_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_264_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_264_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_264_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_264_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_264_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_265_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_265_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_265_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_265_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_265_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_266_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_266_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_266_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_266_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_266_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_267_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_267_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_267_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_267_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_267_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_268_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_268_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_268_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_268_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_268_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_269_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_269_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_269_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_269_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_269_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_270_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_270_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_270_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_270_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_270_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_271_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_271_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_271_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_271_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_271_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_272_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_272_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_272_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_272_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_272_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_273_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_273_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_273_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_273_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_273_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_274_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_274_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_274_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_274_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_274_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_275_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_275_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_275_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_275_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_275_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_276_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_276_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_276_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_276_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_276_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_277_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_277_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_277_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_277_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_277_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_278_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_278_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_278_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_278_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_278_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_10_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_10_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_10_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_10_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_279_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_279_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_279_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_279_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_279_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_280_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_280_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_280_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_280_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_280_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_281_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_281_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_281_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_281_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_281_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_282_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_282_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_282_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_282_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_282_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_283_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_283_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_283_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_283_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_283_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_284_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_284_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_284_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_284_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_284_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_285_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_285_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_285_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_285_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_285_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_286_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_286_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_286_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_286_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_286_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_287_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_287_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_287_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_287_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_287_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_288_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_288_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_288_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_288_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_288_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_289_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_289_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_289_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_289_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_289_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_290_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_290_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_290_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_290_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_290_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_291_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_291_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_291_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_291_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_291_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_292_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_292_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_292_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_292_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_292_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_293_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_293_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_293_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_293_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_293_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_294_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_294_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_294_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_294_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_294_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_295_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_295_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_295_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_295_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_295_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_296_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_296_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_296_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_296_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_296_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_297_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_297_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_297_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_297_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_297_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_298_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_298_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_298_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_298_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_298_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_299_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_299_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_299_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_299_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_299_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_300_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_300_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_300_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_300_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_300_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_301_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_301_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_301_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_301_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_301_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_302_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_302_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_302_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_302_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_302_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_303_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_303_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_303_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_303_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_303_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_11_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_11_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_11_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_11_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_304_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_304_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_304_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_304_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_304_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_305_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_305_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_305_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_305_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_305_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_306_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_306_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_306_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_306_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_306_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_307_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_307_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_307_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_307_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_307_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_308_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_308_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_308_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_308_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_308_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_309_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_309_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_309_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_309_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_309_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_310_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_310_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_310_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_310_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_310_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_311_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_311_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_311_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_311_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_311_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_12_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_12_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_12_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_12_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_312_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_312_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_312_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_312_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_312_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_313_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_313_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_313_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_313_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_313_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_314_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_314_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_314_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_314_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_314_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_315_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_315_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_315_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_315_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_315_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_316_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_316_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_316_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_316_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_316_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_13_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_13_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_13_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_13_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_317_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_317_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_317_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_317_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_317_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_318_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_318_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_318_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_318_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_318_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_14_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_14_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_14_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_14_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_15_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_15_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_15_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_15_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_16_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_16_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_16_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_16_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_319_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_319_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_319_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_319_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_319_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_320_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_320_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_320_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_320_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_320_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_321_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_321_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_321_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_321_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_321_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_322_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_322_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_322_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_322_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_322_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_17_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_17_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_17_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_17_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_323_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_323_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_323_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_323_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_323_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_324_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_324_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_324_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_324_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_324_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_325_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_325_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_325_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_325_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_325_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_326_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_326_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_326_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_326_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_326_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_327_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_327_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_327_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_327_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_327_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_328_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_328_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_328_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_328_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_328_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_18_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_18_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_18_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_18_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_329_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_329_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_329_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_329_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_329_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_330_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_330_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_330_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_330_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_330_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_19_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_19_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_19_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_19_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_331_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_331_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_331_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_331_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_331_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_332_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_332_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_332_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_332_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_332_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_20_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_20_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_20_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_20_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_333_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_333_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_333_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_333_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_333_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_334_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_334_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_334_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_334_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_334_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_335_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_335_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_335_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_335_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_335_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_336_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_336_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_336_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_336_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_336_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_337_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_337_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_337_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_337_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_337_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_338_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_338_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_338_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_338_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_338_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_339_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_339_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_339_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_339_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_339_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_340_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_340_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_340_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_340_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_340_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_341_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_341_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_341_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_341_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_341_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_342_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_342_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_342_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_342_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_342_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_343_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_343_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_343_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_343_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_343_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_344_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_344_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_344_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_344_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_344_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_345_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_345_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_345_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_345_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_345_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_346_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_346_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_346_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_346_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_346_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_347_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_347_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_347_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_347_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_347_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_348_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_348_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_348_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_348_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_348_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_349_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_349_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_349_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_349_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_349_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_350_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_350_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_350_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_350_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_350_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_351_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_351_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_351_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_351_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_351_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_352_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_352_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_352_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_352_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_352_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_353_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_353_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_353_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_353_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_353_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_354_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_354_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_354_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_354_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_354_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_355_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_355_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_355_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_355_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_355_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_356_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_356_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_356_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_356_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_356_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_357_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_357_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_357_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_357_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_357_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_358_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_358_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_358_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_358_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_358_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_359_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_359_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_359_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_359_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_359_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_360_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_360_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_360_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_360_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_360_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_361_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_361_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_361_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_361_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_361_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_362_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_362_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_362_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_362_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_362_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_363_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_363_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_363_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_363_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_363_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_364_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_364_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_364_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_364_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_364_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_365_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_365_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_365_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_365_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_365_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_366_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_366_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_366_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_366_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_366_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_21_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_21_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_21_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_21_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_367_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_367_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_367_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_367_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_367_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_368_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_368_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_368_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_368_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_368_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_369_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_369_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_369_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_369_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_369_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_370_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_370_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_370_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_370_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_370_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_371_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_371_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_371_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_371_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_371_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_372_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_372_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_372_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_372_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_372_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_373_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_373_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_373_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_373_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_373_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_374_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_374_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_374_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_374_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_374_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_375_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_375_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_375_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_375_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_375_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_376_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_376_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_376_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_376_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_376_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_377_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_377_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_377_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_377_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_377_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_378_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_378_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_378_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_378_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_378_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_379_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_379_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_379_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_379_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_379_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_380_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_380_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_380_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_380_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_380_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_381_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_381_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_381_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_381_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_381_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_382_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_382_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_382_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_382_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_382_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_383_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_383_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_383_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_383_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_383_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_384_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_384_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_384_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_384_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_384_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_385_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_385_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_385_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_385_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_385_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_386_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_386_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_386_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_386_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_386_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_22_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_22_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_22_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_22_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_387_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_387_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_387_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_387_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_387_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_388_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_388_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_388_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_388_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_388_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_389_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_389_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_389_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_389_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_389_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_390_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_390_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_390_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_390_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_390_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_391_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_391_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_391_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_391_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_391_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_392_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_392_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_392_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_392_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_392_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_393_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_393_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_393_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_393_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_393_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_394_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_394_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_394_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_394_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_394_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_395_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_395_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_395_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_395_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_395_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_396_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_396_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_396_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_396_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_396_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_397_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_397_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_397_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_397_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_397_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_398_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_398_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_398_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_398_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_398_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_399_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_399_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_399_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_399_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_399_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_400_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_400_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_400_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_400_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_400_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_401_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_401_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_401_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_401_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_401_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_402_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_402_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_402_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_402_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_402_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_403_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_403_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_403_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_403_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_403_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_404_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_404_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_404_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_404_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_404_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_23_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_23_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_23_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_23_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_405_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_405_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_405_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_405_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_405_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_406_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_406_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_406_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_406_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_406_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_407_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_407_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_407_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_407_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_407_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_408_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_408_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_408_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_408_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_408_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_409_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_409_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_409_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_409_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_409_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_410_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_410_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_410_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_410_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_410_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_24_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_24_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_24_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_24_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_411_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_411_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_411_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_411_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_411_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_412_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_412_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_412_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_412_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_412_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_413_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_413_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_413_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_413_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_413_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_414_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_414_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_414_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_414_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_414_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_415_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_415_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_415_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_415_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_415_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_416_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_416_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_416_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_416_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_416_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_417_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_417_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_417_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_417_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_417_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_418_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_418_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_418_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_418_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_418_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_419_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_419_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_419_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_419_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_419_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_420_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_420_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_420_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_420_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_420_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_421_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_421_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_421_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_421_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_421_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_422_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_422_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_422_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_422_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_422_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_423_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_423_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_423_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_423_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_423_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_424_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_424_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_424_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_424_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_424_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_425_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_425_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_425_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_425_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_425_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_426_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_426_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_426_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_426_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_426_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_427_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_427_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_427_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_427_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_427_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_428_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_428_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_428_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_428_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_428_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_429_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_429_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_429_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_429_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_429_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_430_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_430_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_430_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_430_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_430_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_431_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_431_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_431_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_431_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_431_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_432_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_432_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_432_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_432_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_432_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_433_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_433_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_433_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_433_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_433_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_434_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_434_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_434_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_434_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_434_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_435_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_435_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_435_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_435_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_435_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_436_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_436_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_436_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_436_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_436_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_437_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_437_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_437_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_437_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_437_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_438_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_438_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_438_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_438_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_438_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_439_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_439_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_439_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_439_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_439_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_440_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_440_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_440_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_440_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_440_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_441_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_441_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_441_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_441_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_441_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_442_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_442_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_442_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_442_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_442_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_443_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_443_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_443_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_443_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_443_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_444_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_444_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_444_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_444_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_444_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_445_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_445_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_445_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_445_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_445_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_446_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_446_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_446_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_446_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_446_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_447_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_447_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_447_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_447_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_447_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_448_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_448_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_448_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_448_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_448_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_449_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_449_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_449_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_449_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_449_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_450_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_450_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_450_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_450_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_450_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_451_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_451_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_451_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_451_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_451_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_452_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_452_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_452_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_452_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_452_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_453_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_453_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_453_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_453_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_453_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_454_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_454_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_454_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_454_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_454_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_455_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_455_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_455_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_455_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_455_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_456_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_456_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_456_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_456_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_456_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_457_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_457_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_457_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_457_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_457_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_458_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_458_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_458_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_458_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_458_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_459_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_459_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_459_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_459_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_459_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_460_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_460_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_460_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_460_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_460_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_461_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_461_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_461_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_461_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_461_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_462_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_462_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_462_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_462_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_462_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_463_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_463_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_463_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_463_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_463_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_464_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_464_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_464_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_464_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_464_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_465_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_465_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_465_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_465_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_465_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_466_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_466_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_466_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_466_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_466_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_25_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_25_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_25_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_25_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_467_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_467_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_467_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_467_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_467_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_468_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_468_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_468_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_468_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_468_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_469_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_469_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_469_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_469_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_469_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_470_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_470_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_470_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_470_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_470_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_471_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_471_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_471_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_471_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_471_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_26_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_26_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_26_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_26_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_472_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_472_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_472_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_472_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_472_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_473_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_473_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_473_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_473_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_473_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_474_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_474_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_474_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_474_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_474_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_475_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_475_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_475_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_475_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_475_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_476_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_476_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_476_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_476_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_476_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_477_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_477_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_477_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_477_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_477_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_478_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_478_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_478_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_478_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_478_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_479_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_479_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_479_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_479_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_479_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_480_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_480_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_480_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_480_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_480_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_481_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_481_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_481_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_481_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_481_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_482_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_482_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_482_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_482_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_482_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_483_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_483_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_483_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_483_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_483_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_484_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_484_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_484_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_484_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_484_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_485_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_485_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_485_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_485_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_485_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_486_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_486_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_486_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_486_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_486_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_487_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_487_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_487_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_487_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_487_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_488_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_488_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_488_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_488_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_488_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_489_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_489_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_489_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_489_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_489_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_490_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_490_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_490_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_490_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_490_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_491_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_491_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_491_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_491_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_491_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_492_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_492_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_492_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_492_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_492_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_493_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_493_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_493_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_493_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_493_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_494_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_494_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_494_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_494_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_494_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_495_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_495_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_495_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_495_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_495_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_496_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_496_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_496_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_496_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_496_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_497_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_497_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_497_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_497_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_497_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_498_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_498_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_498_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_498_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_498_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_499_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_499_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_499_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_499_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_499_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_500_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_500_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_500_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_500_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_500_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_501_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_501_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_501_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_501_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_501_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_502_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_502_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_502_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_502_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_502_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_503_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_503_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_503_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_503_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_503_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_504_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_504_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_504_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_504_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_504_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_505_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_505_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_505_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_505_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_505_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_27_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_27_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_27_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_27_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_506_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_506_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_506_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_506_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_506_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_507_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_507_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_507_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_507_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_507_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_508_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_508_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_508_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_508_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_508_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_509_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_509_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_509_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_509_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_509_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_510_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_510_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_510_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_510_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_510_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_511_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_511_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_511_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_511_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_511_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_512_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_512_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_512_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_512_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_512_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_513_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_513_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_513_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_513_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_513_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_514_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_514_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_514_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_514_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_514_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_515_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_515_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_515_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_515_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_515_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_516_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_516_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_516_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_516_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_516_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_517_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_517_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_517_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_517_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_517_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_518_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_518_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_518_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_518_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_518_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_519_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_519_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_519_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_519_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_519_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_28_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_28_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_28_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_28_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_520_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_520_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_520_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_520_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_520_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_521_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_521_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_521_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_521_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_521_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_522_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_522_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_522_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_522_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_522_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_523_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_523_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_523_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_523_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_523_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_524_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_524_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_524_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_524_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_524_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_525_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_525_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_525_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_525_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_525_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_526_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_526_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_526_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_526_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_526_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_29_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_29_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_29_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_29_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_527_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_527_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_527_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_527_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_527_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_30_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_30_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_30_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_30_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_31_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_31_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_31_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_31_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_32_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_32_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_32_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_32_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_33_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_33_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_33_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_33_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_528_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_528_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_528_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_528_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_528_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_34_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_34_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_34_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_34_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_35_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_35_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_35_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_35_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_36_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_36_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_36_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_36_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_529_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_529_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_529_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_529_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_529_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_530_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_530_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_530_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_530_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_530_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_531_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_531_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_531_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_531_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_531_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_532_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_532_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_532_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_532_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_532_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_533_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_533_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_533_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_533_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_533_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_534_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_534_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_534_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_534_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_534_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_37_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_37_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_37_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_37_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_535_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_535_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_535_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_535_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_535_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_536_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_536_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_536_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_536_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_536_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_537_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_537_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_537_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_537_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_537_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_538_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_538_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_538_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_538_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_538_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_539_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_539_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_539_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_539_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_539_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_540_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_540_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_540_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_540_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_540_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_541_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_541_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_541_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_541_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_541_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_542_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_542_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_542_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_542_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_542_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_543_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_543_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_543_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_543_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_543_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_544_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_544_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_544_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_544_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_544_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_545_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_545_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_545_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_545_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_545_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_546_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_546_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_546_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_546_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_546_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_38_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_38_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_38_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_38_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_547_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_547_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_547_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_547_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_547_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_548_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_548_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_548_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_548_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_548_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_39_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_39_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_39_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_39_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_549_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_549_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_549_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_549_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_549_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_550_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_550_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_550_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_550_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_550_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_40_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_40_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_40_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_40_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_551_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_551_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_551_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_551_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_551_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_552_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_552_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_552_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_552_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_552_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_41_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_41_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_41_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_41_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_553_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_553_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_553_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_553_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_553_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_554_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_554_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_554_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_554_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_554_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_555_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_555_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_555_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_555_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_555_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_556_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_556_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_556_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_556_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_556_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_557_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_557_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_557_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_557_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_557_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_558_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_558_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_558_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_558_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_558_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_559_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_559_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_559_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_559_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_559_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_560_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_560_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_560_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_560_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_560_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_561_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_561_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_561_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_561_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_561_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_562_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_562_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_562_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_562_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_562_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_563_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_563_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_563_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_563_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_563_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_564_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_564_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_564_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_564_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_564_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_42_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_42_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_42_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_42_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_565_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_565_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_565_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_565_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_565_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_566_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_566_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_566_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_566_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_566_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_567_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_567_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_567_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_567_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_567_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_43_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_43_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_43_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_43_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_568_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_568_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_568_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_568_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_568_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_569_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_569_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_569_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_569_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_569_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_570_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_570_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_570_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_570_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_570_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_571_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_571_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_571_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_571_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_571_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_572_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_572_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_572_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_572_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_572_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_573_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_573_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_573_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_573_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_573_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_574_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_574_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_574_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_574_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_574_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_575_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_575_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_575_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_575_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_575_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_576_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_576_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_576_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_576_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_576_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_577_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_577_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_577_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_577_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_577_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_578_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_578_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_578_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_578_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_578_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_579_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_579_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_579_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_579_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_579_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_580_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_580_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_580_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_580_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_580_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_581_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_581_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_581_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_581_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_581_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_582_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_582_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_582_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_582_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_582_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_583_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_583_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_583_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_583_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_583_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_584_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_584_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_584_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_584_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_584_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_585_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_585_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_585_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_585_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_585_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_586_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_586_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_586_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_586_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_586_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_587_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_587_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_587_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_587_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_587_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_44_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_44_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_44_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_44_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_588_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_588_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_588_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_588_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_588_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_589_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_589_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_589_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_589_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_589_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_590_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_590_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_590_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_590_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_590_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_591_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_591_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_591_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_591_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_591_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_592_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_592_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_592_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_592_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_592_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_593_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_593_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_593_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_593_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_593_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_594_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_594_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_594_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_594_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_594_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_595_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_595_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_595_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_595_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_595_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_596_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_596_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_596_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_596_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_596_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_597_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_597_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_597_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_597_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_597_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_598_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_598_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_598_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_598_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_598_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_599_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_599_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_599_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_599_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_599_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_600_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_600_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_600_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_600_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_600_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_45_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_45_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_45_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_45_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_601_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_601_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_601_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_601_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_601_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_602_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_602_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_602_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_602_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_602_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_603_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_603_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_603_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_603_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_603_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_604_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_604_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_604_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_604_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_604_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_605_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_605_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_605_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_605_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_605_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_606_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_606_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_606_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_606_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_606_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_607_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_607_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_607_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_607_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_607_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_608_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_608_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_608_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_608_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_608_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_609_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_609_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_609_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_609_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_609_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_610_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_610_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_610_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_610_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_610_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_611_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_611_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_611_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_611_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_611_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_612_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_612_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_612_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_612_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_612_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_613_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_613_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_613_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_613_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_613_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_614_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_614_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_614_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_614_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_614_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_615_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_615_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_615_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_615_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_615_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_616_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_616_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_616_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_616_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_616_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_617_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_617_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_617_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_617_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_617_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_618_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_618_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_618_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_618_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_618_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_619_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_619_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_619_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_619_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_619_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_620_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_620_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_620_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_620_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_620_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_621_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_621_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_621_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_621_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_621_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_622_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_622_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_622_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_622_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_622_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_623_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_623_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_623_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_623_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_623_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_624_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_624_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_624_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_624_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_624_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_625_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_625_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_625_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_625_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_625_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_626_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_626_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_626_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_626_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_626_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_627_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_627_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_627_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_627_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_627_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_628_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_628_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_628_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_628_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_628_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_629_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_629_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_629_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_629_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_629_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_630_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_630_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_630_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_630_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_630_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_631_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_631_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_631_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_631_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_631_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_632_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_632_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_632_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_632_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_632_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_46_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_46_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_46_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_46_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_633_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_633_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_633_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_633_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_633_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_634_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_634_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_634_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_634_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_634_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_635_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_635_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_635_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_635_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_635_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_636_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_636_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_636_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_636_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_636_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_637_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_637_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_637_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_637_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_637_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_638_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_638_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_638_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_638_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_638_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_639_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_639_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_639_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_639_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_639_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_640_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_640_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_640_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_640_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_640_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_641_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_641_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_641_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_641_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_641_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_642_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_642_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_642_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_642_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_642_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_643_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_643_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_643_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_643_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_643_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_644_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_644_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_644_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_644_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_644_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_645_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_645_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_645_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_645_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_645_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_646_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_646_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_646_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_646_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_646_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_647_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_647_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_647_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_647_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_647_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_648_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_648_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_648_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_648_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_648_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_649_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_649_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_649_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_649_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_649_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_650_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_650_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_650_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_650_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_650_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_651_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_651_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_651_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_651_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_651_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_652_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_652_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_652_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_652_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_652_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_47_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_47_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_47_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_47_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_653_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_653_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_653_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_653_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_653_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_654_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_654_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_654_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_654_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_654_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_655_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_655_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_655_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_655_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_655_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_656_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_656_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_656_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_656_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_656_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_657_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_657_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_657_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_657_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_657_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_658_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_658_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_658_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_658_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_658_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_659_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_659_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_659_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_659_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_659_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_660_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_660_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_660_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_660_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_660_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_661_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_661_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_661_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_661_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_661_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_662_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_662_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_662_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_662_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_662_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_663_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_663_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_663_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_663_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_663_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_48_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_48_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_48_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_48_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_664_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_664_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_664_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_664_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_664_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_49_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_49_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_49_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_49_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_665_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_665_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_665_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_665_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_665_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_50_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_50_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_50_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_50_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_666_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_666_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_666_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_666_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_666_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_667_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_667_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_667_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_667_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_667_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_668_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_668_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_668_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_668_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_668_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_51_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_51_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_51_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_51_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_52_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_52_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_52_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_52_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_53_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_53_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_53_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_53_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_54_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_54_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_54_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_54_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_55_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_55_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_55_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_55_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_56_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_56_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_56_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_56_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_669_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_669_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_669_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_669_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_669_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_670_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_670_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_670_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_670_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_670_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_671_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_671_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_671_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_671_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_671_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_672_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_672_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_672_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_672_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_672_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_673_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_673_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_673_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_673_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_673_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_674_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_674_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_674_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_674_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_674_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_675_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_675_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_675_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_675_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_675_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_676_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_676_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_676_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_676_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_676_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_57_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_57_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_57_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_57_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_58_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_58_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_58_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_58_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_59_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_59_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_59_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_59_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_60_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_60_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_60_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_60_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_677_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_677_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_677_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_677_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_677_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_678_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_678_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_678_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_678_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_678_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_679_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_679_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_679_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_679_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_679_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_680_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_680_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_680_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_680_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_680_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_681_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_681_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_681_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_681_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_681_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_682_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_682_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_682_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_682_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_682_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_683_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_683_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_683_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_683_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_683_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_684_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_684_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_684_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_684_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_684_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_685_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_685_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_685_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_685_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_685_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_686_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_686_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_686_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_686_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_686_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_687_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_687_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_687_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_687_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_687_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_688_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_688_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_688_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_688_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_688_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_689_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_689_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_689_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_689_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_689_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_690_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_690_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_690_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_690_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_690_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_691_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_691_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_691_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_691_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_691_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_61_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_61_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_61_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_61_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_62_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_62_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_62_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_62_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_692_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_692_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_692_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_692_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_692_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_693_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_693_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_693_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_693_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_693_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_694_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_694_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_694_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_694_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_694_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_695_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_695_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_695_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_695_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_695_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_63_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_63_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_63_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_63_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_696_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_696_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_696_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_696_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_696_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_697_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_697_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_697_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_697_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_697_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_698_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_698_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_698_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_698_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_698_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_699_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_699_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_699_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_699_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_699_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_700_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_700_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_700_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_700_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_700_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_701_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_701_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_701_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_701_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_701_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_702_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_702_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_702_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_702_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_702_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_703_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_703_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_703_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_703_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_703_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_704_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_704_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_704_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_704_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_704_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_705_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_705_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_705_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_705_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_705_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_706_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_706_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_706_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_706_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_706_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_707_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_707_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_707_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_707_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_707_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_708_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_708_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_708_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_708_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_708_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_709_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_709_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_709_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_709_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_709_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_710_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_710_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_710_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_710_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_710_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_711_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_711_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_711_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_711_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_711_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_712_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_712_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_712_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_712_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_712_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_713_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_713_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_713_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_713_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_713_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_714_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_714_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_714_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_714_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_714_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_715_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_715_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_715_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_715_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_715_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_716_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_716_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_716_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_716_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_716_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_717_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_717_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_717_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_717_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_717_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_718_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_718_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_718_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_718_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_718_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_719_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_719_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_719_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_719_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_719_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_720_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_720_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_720_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_720_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_720_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_721_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_721_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_721_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_721_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_721_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_722_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_722_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_722_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_722_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_722_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_723_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_723_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_723_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_723_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_723_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_724_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_724_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_724_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_724_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_724_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_725_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_725_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_725_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_725_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_725_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_726_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_726_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_726_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_726_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_726_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_727_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_727_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_727_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_727_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_727_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_728_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_728_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_728_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_728_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_728_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_729_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_729_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_729_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_729_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_729_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_730_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_730_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_730_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_730_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_730_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_731_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_731_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_731_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_731_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_731_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_732_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_732_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_732_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_732_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_732_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_64_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_64_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_64_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_64_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_733_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_733_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_733_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_733_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_733_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_734_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_734_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_734_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_734_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_734_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_65_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_65_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_65_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_65_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_735_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_735_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_735_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_735_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_735_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_736_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_736_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_736_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_736_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_736_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_737_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_737_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_737_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_737_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_737_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_738_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_738_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_738_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_738_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_738_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_739_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_739_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_739_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_739_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_739_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_740_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_740_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_740_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_740_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_740_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_741_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_741_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_741_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_741_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_741_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_742_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_742_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_742_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_742_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_742_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_743_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_743_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_743_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_743_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_743_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_744_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_744_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_744_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_744_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_744_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_745_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_745_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_745_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_745_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_745_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_746_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_746_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_746_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_746_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_746_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_747_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_747_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_747_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_747_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_747_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_748_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_748_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_748_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_748_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_748_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_749_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_749_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_749_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_749_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_749_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_66_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_66_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_66_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_66_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_750_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_750_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_750_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_750_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_750_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_67_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_67_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_67_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_67_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_751_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_751_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_751_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_751_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_751_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_752_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_752_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_752_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_752_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_752_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_753_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_753_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_753_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_753_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_753_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_754_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_754_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_754_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_754_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_754_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_68_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_68_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_68_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_68_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_69_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_69_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_69_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_69_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_755_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_755_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_755_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_755_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_755_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_756_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_756_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_756_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_756_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_756_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_70_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_70_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_70_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_70_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_757_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_757_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_757_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_757_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_757_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_758_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_758_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_758_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_758_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_758_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_71_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_71_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_71_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_71_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_72_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_72_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_72_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_72_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_73_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_73_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_73_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_73_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_74_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_74_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_74_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_74_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_75_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_75_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_75_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_75_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_759_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_759_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_759_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_759_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_759_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_76_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_76_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_76_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_76_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_77_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_77_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_77_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_77_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_760_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_760_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_760_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_760_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_760_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_761_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_761_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_761_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_761_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_761_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_762_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_762_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_762_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_762_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_762_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_763_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_763_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_763_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_763_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_763_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_764_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_764_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_764_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_764_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_764_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_765_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_765_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_765_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_765_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_765_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_78_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_78_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_78_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_78_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_79_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_79_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_79_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_79_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_80_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_80_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_80_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_80_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_766_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_766_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_766_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_766_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_766_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_767_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_767_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_767_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_767_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_767_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_768_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_768_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_768_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_768_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_768_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_769_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_769_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_769_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_769_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_769_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_770_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_770_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_770_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_770_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_770_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_81_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_81_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_81_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_81_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_771_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_771_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_771_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_771_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_771_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_772_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_772_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_772_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_772_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_772_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_773_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_773_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_773_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_773_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_773_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_82_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_82_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_82_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_82_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_83_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_83_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_83_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_83_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_84_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_84_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_84_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_84_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_774_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_774_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_774_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_774_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_774_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_775_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_775_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_775_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_775_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_775_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_776_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_776_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_776_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_776_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_776_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_85_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_85_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_85_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_85_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_777_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_777_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_777_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_777_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_777_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_778_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_778_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_778_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_778_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_778_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_779_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_779_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_779_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_779_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_779_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_780_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_780_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_780_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_780_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_780_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_781_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_781_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_781_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_781_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_781_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_782_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_782_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_782_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_782_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_782_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_783_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_783_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_783_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_783_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_783_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_784_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_784_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_784_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_784_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_784_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_785_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_785_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_785_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_785_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_785_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_786_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_786_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_786_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_786_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_786_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_787_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_787_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_787_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_787_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_787_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_788_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_788_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_788_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_788_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_788_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_789_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_789_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_789_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_789_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_789_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_790_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_790_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_790_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_790_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_790_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_791_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_791_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_791_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_791_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_791_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_792_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_792_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_792_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_792_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_792_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_793_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_793_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_793_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_793_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_793_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_794_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_794_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_794_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_794_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_794_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_795_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_795_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_795_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_795_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_795_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_796_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_796_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_796_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_796_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_796_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_797_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_797_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_797_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_797_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_797_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_798_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_798_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_798_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_798_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_798_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_799_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_799_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_799_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_799_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_799_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_800_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_800_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_800_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_800_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_800_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_801_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_801_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_801_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_801_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_801_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_802_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_802_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_802_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_802_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_802_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_803_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_803_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_803_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_803_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_803_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_86_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_86_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_86_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_86_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_87_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_87_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_87_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_87_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_88_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_88_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_88_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_88_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_804_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_804_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_804_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_804_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_804_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_89_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_89_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_89_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_89_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_805_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_805_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_805_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_805_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_805_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_806_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_806_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_806_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_806_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_806_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_807_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_807_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_807_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_807_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_807_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_808_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_808_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_808_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_808_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_808_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_809_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_809_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_809_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_809_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_809_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_810_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_810_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_810_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_810_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_810_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_811_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_811_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_811_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_811_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_811_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_90_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_90_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_90_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_90_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_91_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_91_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_91_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_91_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_812_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_812_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_812_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_812_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_812_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_813_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_813_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_813_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_813_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_813_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_814_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_814_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_814_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_814_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_814_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_92_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_92_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_92_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_92_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_815_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_815_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_815_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_815_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_815_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_816_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_816_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_816_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_816_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_816_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_93_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_93_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_93_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_93_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_94_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_94_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_94_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_94_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_95_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_95_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_95_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_95_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_96_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_96_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_96_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_96_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_97_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_97_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_97_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_97_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_98_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_98_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_98_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_98_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_99_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_99_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_99_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_99_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_100_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_100_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_100_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_100_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_101_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_101_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_101_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_101_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_817_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_817_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_817_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_817_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_817_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_102_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_102_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_102_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_102_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_103_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_103_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_103_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_103_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_818_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_818_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_818_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_818_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_818_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_819_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_819_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_819_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_819_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_819_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_104_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_104_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_104_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_104_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_105_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_105_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_105_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_105_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_820_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_820_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_820_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_820_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_820_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_821_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_821_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_821_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_821_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_821_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_822_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_822_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_822_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_822_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_822_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_823_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_823_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_823_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_823_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_823_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_824_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_824_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_824_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_824_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_824_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_825_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_825_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_825_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_825_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_825_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_826_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_826_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_826_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_826_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_826_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_827_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_827_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_827_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_827_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_827_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_106_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_106_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_106_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_106_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_107_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_107_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_107_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_107_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_828_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_828_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_828_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_828_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_828_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_108_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_108_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_108_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_108_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_109_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_109_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_109_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_109_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_829_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_829_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_829_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_829_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_829_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_830_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_830_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_830_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_830_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_830_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_831_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_831_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_831_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_831_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_831_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_110_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_110_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_110_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_110_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_832_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_832_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_832_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_832_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_832_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_833_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_833_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_833_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_833_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_833_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_111_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_111_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_111_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_111_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_834_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_834_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_834_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_834_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_834_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_835_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_835_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_835_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_835_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_835_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_836_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_836_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_836_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_836_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_836_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_837_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_837_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_837_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_837_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_837_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_838_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_838_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_838_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_838_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_838_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_839_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_839_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_839_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_839_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_839_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_840_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_840_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_840_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_840_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_840_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_841_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_841_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_841_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_841_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_841_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_842_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_842_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_842_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_842_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_842_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_112_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_112_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_112_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_112_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_113_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_113_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_113_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_113_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_843_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_843_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_843_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_843_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_843_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_844_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_844_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_844_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_844_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_844_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_845_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_845_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_845_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_845_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_845_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_846_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_846_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_846_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_846_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_846_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_847_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_847_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_847_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_847_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_847_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_848_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_848_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_848_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_848_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_848_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_849_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_849_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_849_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_849_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_849_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_114_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_114_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_114_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_114_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_850_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_850_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_850_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_850_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_850_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_115_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_115_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_115_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_115_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_116_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_116_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_116_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_116_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_117_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_117_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_117_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_117_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_851_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_851_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_851_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_851_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_851_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_118_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_118_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_118_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_118_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_852_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_852_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_852_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_852_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_852_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_119_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_119_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_119_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_119_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_853_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_853_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_853_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_853_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_853_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_120_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_120_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_120_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_120_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_121_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_121_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_121_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_121_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_122_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_122_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_122_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_122_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_854_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_854_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_854_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_854_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_854_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_855_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_855_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_855_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_855_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_855_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_856_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_856_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_856_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_856_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_856_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_123_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_123_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_123_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_123_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_124_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_124_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_124_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_124_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_125_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_125_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_125_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_125_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_126_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_126_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_126_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_126_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_857_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_857_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_857_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_857_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_857_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_858_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_858_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_858_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_858_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_858_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_127_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_127_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_127_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_127_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_128_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_128_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_128_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_128_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_859_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_859_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_859_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_859_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_859_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_129_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_129_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_129_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_129_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_860_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_860_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_860_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_860_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_860_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_861_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_861_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_861_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_861_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_861_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_862_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_862_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_862_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_862_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_862_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_863_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_863_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_863_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_863_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_863_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_864_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_864_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_864_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_864_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_864_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_865_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_865_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_865_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_865_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_865_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_866_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_866_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_866_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_866_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_866_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_867_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_867_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_867_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_867_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_867_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_868_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_868_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_868_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_868_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_868_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_869_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_869_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_869_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_869_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_869_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_870_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_870_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_870_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_870_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_870_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_130_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_130_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_130_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_130_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_871_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_871_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_871_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_871_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_871_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_872_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_872_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_872_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_872_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_872_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_131_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_131_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_131_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_131_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_132_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_132_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_132_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_132_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_873_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_873_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_873_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_873_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_873_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_874_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_874_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_874_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_874_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_874_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_875_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_875_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_875_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_875_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_875_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_133_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_133_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_133_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_133_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_876_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_876_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_876_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_876_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_876_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_877_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_877_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_877_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_877_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_877_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_134_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_134_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_134_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_134_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_878_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_878_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_878_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_878_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_878_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_135_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_135_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_135_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_135_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_136_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_136_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_136_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_136_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_137_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_137_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_137_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_137_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_138_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_138_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_138_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_138_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_139_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_139_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_139_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_139_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_140_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_140_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_140_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_140_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_879_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_879_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_879_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_879_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_879_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_141_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_141_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_141_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_141_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_142_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_142_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_142_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_142_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_880_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_880_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_880_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_880_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_880_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_143_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_143_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_143_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_143_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_881_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_881_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_881_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_881_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_881_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_144_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_144_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_144_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_144_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_145_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_145_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_145_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_145_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_882_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_882_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_882_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_882_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_882_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_883_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_883_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_883_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_883_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_883_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_146_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_146_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_146_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_146_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_884_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_884_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_884_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_884_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_884_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_147_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_147_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_147_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_147_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_885_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_885_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_885_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_885_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_885_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_886_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_886_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_886_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_886_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_886_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_148_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_148_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_148_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_148_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_149_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_149_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_149_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_149_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_887_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_887_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_887_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_887_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_887_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_888_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_888_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_888_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_888_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_888_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_889_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_889_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_889_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_889_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_889_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_150_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_150_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_150_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_150_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_151_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_151_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_151_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_151_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_152_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_152_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_152_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_152_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_890_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_890_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_890_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_890_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_890_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_153_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_153_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_153_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_153_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_891_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_891_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_891_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_891_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_891_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_892_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_892_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_892_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_892_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_892_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_154_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_154_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_154_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_154_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_893_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_893_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_893_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_893_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_893_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_155_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_155_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_155_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_155_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_156_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_156_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_156_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_156_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_157_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_157_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_157_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_157_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_894_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_894_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_894_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_894_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_894_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_158_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_158_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_158_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_158_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_159_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_159_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_159_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_159_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_160_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_160_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_160_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_160_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_895_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_895_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_895_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_895_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_895_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_161_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_161_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_161_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_161_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_162_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_162_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_162_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_162_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_896_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_896_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_896_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_896_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_896_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_163_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_163_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_163_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_163_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_164_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_164_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_164_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_164_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_897_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_897_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_897_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_897_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_897_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_898_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_898_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_898_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_898_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_898_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_165_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_165_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_165_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_165_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_899_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_899_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_899_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_899_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_899_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_166_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_166_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_166_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_166_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_167_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_167_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_167_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_167_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_900_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_900_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_900_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_900_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_900_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_901_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_901_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_901_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_901_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_901_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_168_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_168_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_168_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_168_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_169_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_169_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_169_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_169_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_902_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_902_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_902_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_902_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_902_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_170_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_170_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_170_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_170_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_903_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_903_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_903_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_903_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_903_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_904_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_904_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_904_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_904_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_904_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_905_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_905_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_905_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_905_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_905_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_171_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_171_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_171_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_171_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_906_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_906_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_906_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_906_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_906_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_907_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_907_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_907_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_907_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_907_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_908_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_908_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_908_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_908_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_908_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_172_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_172_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_172_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_172_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_173_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_173_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_173_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_173_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_909_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_909_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_909_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_909_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_909_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_174_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_174_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_174_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_174_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_175_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_175_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_175_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_175_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_176_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_176_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_176_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_176_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_910_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_910_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_910_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_910_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_910_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_177_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_177_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_177_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_177_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_911_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_911_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_911_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_911_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_911_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_912_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_912_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_912_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_912_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_912_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_178_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_178_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_178_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_178_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_913_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_913_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_913_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_913_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_913_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_914_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_914_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_914_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_914_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_914_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_179_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_179_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_179_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_179_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_180_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_180_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_180_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_180_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_915_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_915_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_915_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_915_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_915_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_181_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_181_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_181_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_181_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_182_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_182_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_182_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_182_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_916_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_916_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_916_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_916_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_916_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_183_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_183_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_183_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_183_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_917_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_917_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_917_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_917_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_917_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_918_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_918_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_918_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_918_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_918_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_919_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_919_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_919_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_919_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_919_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_184_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_184_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_184_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_184_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_185_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_185_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_185_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_185_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_920_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_920_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_920_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_920_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_920_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_186_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_186_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_186_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_186_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_921_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_921_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_921_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_921_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_921_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_922_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_922_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_922_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_922_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_922_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_187_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_187_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_187_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_187_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_923_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_923_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_923_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_923_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_923_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_924_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_924_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_924_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_924_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_924_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_925_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_925_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_925_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_925_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_925_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_926_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_926_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_926_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_926_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_926_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_927_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_927_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_927_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_927_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_927_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_928_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_928_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_928_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_928_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_928_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_929_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_929_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_929_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_929_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_929_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_188_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_188_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_188_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_188_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_930_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_930_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_930_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_930_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_930_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_189_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_189_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_189_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_189_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_190_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_190_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_190_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_190_io_co; // @[wallace.scala 57:25]
  wire  res0_0 = io_pp_0[0]; // @[wallace.scala 34:43]
  wire  res0_1 = io_pp_0[1]; // @[wallace.scala 34:43]
  wire  res1_1 = io_pp_1[0]; // @[wallace.scala 34:43]
  wire  res0_62 = HalfAdder_139_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_61 = FullAdder_906_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_60 = HalfAdder_158_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_59 = HalfAdder_140_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_58 = FullAdder_915_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_57 = FullAdder_907_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_56 = HalfAdder_159_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_55 = FullAdder_879_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_54 = HalfAdder_160_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_53 = FullAdder_930_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [9:0] _T_1032 = {res0_62,res0_61,res0_60,res0_59,res0_58,res0_57,res0_56,res0_55,res0_54,res0_53}; // @[Cat.scala 29:58]
  wire  res0_52 = FullAdder_929_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_51 = FullAdder_925_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_50 = HalfAdder_190_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_49 = HalfAdder_189_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_48 = HalfAdder_188_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_47 = FullAdder_926_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_46 = FullAdder_921_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_45 = HalfAdder_182_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_44 = FullAdder_927_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [18:0] _T_1041 = {_T_1032,res0_52,res0_51,res0_50,res0_49,res0_48,res0_47,res0_46,res0_45,res0_44}; // @[Cat.scala 29:58]
  wire  res0_43 = FullAdder_922_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_42 = FullAdder_928_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_41 = HalfAdder_187_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_40 = FullAdder_917_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_39 = HalfAdder_176_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_38 = FullAdder_923_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_37 = FullAdder_918_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_36 = FullAdder_910_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_35 = HalfAdder_177_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [27:0] _T_1050 = {_T_1041,res0_43,res0_42,res0_41,res0_40,res0_39,res0_38,res0_37,res0_36,res0_35}; // @[Cat.scala 29:58]
  wire  res0_34 = FullAdder_900_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_33 = FullAdder_887_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_32 = FullAdder_888_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_31 = FullAdder_911_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_30 = FullAdder_901_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_29 = FullAdder_919_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_28 = FullAdder_924_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_27 = HalfAdder_184_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_26 = HalfAdder_169_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [36:0] _T_1059 = {_T_1050,res0_34,res0_33,res0_32,res0_31,res0_30,res0_29,res0_28,res0_27,res0_26}; // @[Cat.scala 29:58]
  wire  res0_25 = FullAdder_902_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_24 = HalfAdder_170_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_23 = HalfAdder_185_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_22 = FullAdder_913_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_21 = FullAdder_903_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_20 = FullAdder_891_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_19 = FullAdder_874_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_18 = FullAdder_892_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_17 = HalfAdder_154_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [45:0] _T_1068 = {_T_1059,res0_25,res0_24,res0_23,res0_22,res0_21,res0_20,res0_19,res0_18,res0_17}; // @[Cat.scala 29:58]
  wire  res0_16 = HalfAdder_133_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_15 = FullAdder_893_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_14 = FullAdder_914_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_13 = FullAdder_904_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_12 = HalfAdder_179_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_11 = FullAdder_905_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_10 = FullAdder_920_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_9 = HalfAdder_180_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_8 = HalfAdder_171_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [54:0] _T_1077 = {_T_1068,res0_16,res0_15,res0_14,res0_13,res0_12,res0_11,res0_10,res0_9,res0_8}; // @[Cat.scala 29:58]
  wire  res0_7 = FullAdder_894_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_6 = HalfAdder_138_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_5 = HalfAdder_96_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_4 = FullAdder_528_io_co; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_3 = FullAdder_528_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_2 = FullAdder_318_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [62:0] _T_1085 = {_T_1077,res0_7,res0_6,res0_5,res0_4,res0_3,res0_2,res0_1,res0_0}; // @[Cat.scala 29:58]
  wire  res1_62 = FullAdder_906_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_59 = FullAdder_915_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_55 = HalfAdder_160_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_54 = FullAdder_930_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [9:0] _T_1094 = {res1_62,1'h0,1'h0,res1_59,1'h0,1'h0,1'h0,res1_55,res1_54,1'h0}; // @[Cat.scala 29:58]
  wire  res1_51 = HalfAdder_190_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_45 = FullAdder_927_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [18:0] _T_1103 = {_T_1094,1'h0,res1_51,1'h0,1'h0,1'h0,1'h0,1'h0,res1_45,1'h0}; // @[Cat.scala 29:58]
  wire  res1_43 = FullAdder_928_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_39 = FullAdder_923_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_36 = HalfAdder_177_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [27:0] _T_1112 = {_T_1103,res1_43,1'h0,1'h0,1'h0,res1_39,1'h0,1'h0,res1_36,1'h0}; // @[Cat.scala 29:58]
  wire  res1_33 = FullAdder_888_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_32 = FullAdder_911_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_30 = FullAdder_919_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_29 = FullAdder_924_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_26 = FullAdder_902_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [36:0] _T_1121 = {_T_1112,1'h0,res1_33,res1_32,1'h0,res1_30,res1_29,1'h0,1'h0,res1_26}; // @[Cat.scala 29:58]
  wire  res1_25 = HalfAdder_170_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_24 = HalfAdder_185_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_19 = FullAdder_892_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_18 = HalfAdder_154_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [45:0] _T_1130 = {_T_1121,res1_25,res1_24,1'h0,1'h0,1'h0,1'h0,res1_19,res1_18,1'h0}; // @[Cat.scala 29:58]
  wire  res1_16 = FullAdder_893_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_15 = FullAdder_914_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_13 = HalfAdder_179_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_11 = FullAdder_920_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [54:0] _T_1139 = {_T_1130,res1_16,res1_15,1'h0,res1_13,1'h0,res1_11,1'h0,1'h0,1'h0}; // @[Cat.scala 29:58]
  wire  res1_4 = HalfAdder_52_io_s; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [62:0] _T_1147 = {_T_1139,1'h0,1'h0,1'h0,res1_4,1'h0,1'h0,res1_1,1'h0}; // @[Cat.scala 29:58]
  HalfAdder HalfAdder ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_io_a),
    .io_b(HalfAdder_io_b),
    .io_s(HalfAdder_io_s),
    .io_co(HalfAdder_io_co)
  );
  HalfAdder HalfAdder_1 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_1_io_a),
    .io_b(HalfAdder_1_io_b),
    .io_s(HalfAdder_1_io_s),
    .io_co(HalfAdder_1_io_co)
  );
  FullAdder FullAdder ( // @[wallace.scala 67:25]
    .io_a(FullAdder_io_a),
    .io_b(FullAdder_io_b),
    .io_ci(FullAdder_io_ci),
    .io_s(FullAdder_io_s),
    .io_co(FullAdder_io_co)
  );
  FullAdder FullAdder_1 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1_io_a),
    .io_b(FullAdder_1_io_b),
    .io_ci(FullAdder_1_io_ci),
    .io_s(FullAdder_1_io_s),
    .io_co(FullAdder_1_io_co)
  );
  HalfAdder HalfAdder_2 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_2_io_a),
    .io_b(HalfAdder_2_io_b),
    .io_s(HalfAdder_2_io_s),
    .io_co(HalfAdder_2_io_co)
  );
  FullAdder FullAdder_2 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2_io_a),
    .io_b(FullAdder_2_io_b),
    .io_ci(FullAdder_2_io_ci),
    .io_s(FullAdder_2_io_s),
    .io_co(FullAdder_2_io_co)
  );
  FullAdder FullAdder_3 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3_io_a),
    .io_b(FullAdder_3_io_b),
    .io_ci(FullAdder_3_io_ci),
    .io_s(FullAdder_3_io_s),
    .io_co(FullAdder_3_io_co)
  );
  FullAdder FullAdder_4 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_4_io_a),
    .io_b(FullAdder_4_io_b),
    .io_ci(FullAdder_4_io_ci),
    .io_s(FullAdder_4_io_s),
    .io_co(FullAdder_4_io_co)
  );
  FullAdder FullAdder_5 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_5_io_a),
    .io_b(FullAdder_5_io_b),
    .io_ci(FullAdder_5_io_ci),
    .io_s(FullAdder_5_io_s),
    .io_co(FullAdder_5_io_co)
  );
  FullAdder FullAdder_6 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_6_io_a),
    .io_b(FullAdder_6_io_b),
    .io_ci(FullAdder_6_io_ci),
    .io_s(FullAdder_6_io_s),
    .io_co(FullAdder_6_io_co)
  );
  FullAdder FullAdder_7 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_7_io_a),
    .io_b(FullAdder_7_io_b),
    .io_ci(FullAdder_7_io_ci),
    .io_s(FullAdder_7_io_s),
    .io_co(FullAdder_7_io_co)
  );
  FullAdder FullAdder_8 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_8_io_a),
    .io_b(FullAdder_8_io_b),
    .io_ci(FullAdder_8_io_ci),
    .io_s(FullAdder_8_io_s),
    .io_co(FullAdder_8_io_co)
  );
  FullAdder FullAdder_9 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_9_io_a),
    .io_b(FullAdder_9_io_b),
    .io_ci(FullAdder_9_io_ci),
    .io_s(FullAdder_9_io_s),
    .io_co(FullAdder_9_io_co)
  );
  FullAdder FullAdder_10 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_10_io_a),
    .io_b(FullAdder_10_io_b),
    .io_ci(FullAdder_10_io_ci),
    .io_s(FullAdder_10_io_s),
    .io_co(FullAdder_10_io_co)
  );
  FullAdder FullAdder_11 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_11_io_a),
    .io_b(FullAdder_11_io_b),
    .io_ci(FullAdder_11_io_ci),
    .io_s(FullAdder_11_io_s),
    .io_co(FullAdder_11_io_co)
  );
  FullAdder FullAdder_12 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_12_io_a),
    .io_b(FullAdder_12_io_b),
    .io_ci(FullAdder_12_io_ci),
    .io_s(FullAdder_12_io_s),
    .io_co(FullAdder_12_io_co)
  );
  FullAdder FullAdder_13 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_13_io_a),
    .io_b(FullAdder_13_io_b),
    .io_ci(FullAdder_13_io_ci),
    .io_s(FullAdder_13_io_s),
    .io_co(FullAdder_13_io_co)
  );
  FullAdder FullAdder_14 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_14_io_a),
    .io_b(FullAdder_14_io_b),
    .io_ci(FullAdder_14_io_ci),
    .io_s(FullAdder_14_io_s),
    .io_co(FullAdder_14_io_co)
  );
  FullAdder FullAdder_15 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_15_io_a),
    .io_b(FullAdder_15_io_b),
    .io_ci(FullAdder_15_io_ci),
    .io_s(FullAdder_15_io_s),
    .io_co(FullAdder_15_io_co)
  );
  FullAdder FullAdder_16 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_16_io_a),
    .io_b(FullAdder_16_io_b),
    .io_ci(FullAdder_16_io_ci),
    .io_s(FullAdder_16_io_s),
    .io_co(FullAdder_16_io_co)
  );
  HalfAdder HalfAdder_3 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_3_io_a),
    .io_b(HalfAdder_3_io_b),
    .io_s(HalfAdder_3_io_s),
    .io_co(HalfAdder_3_io_co)
  );
  FullAdder FullAdder_17 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_17_io_a),
    .io_b(FullAdder_17_io_b),
    .io_ci(FullAdder_17_io_ci),
    .io_s(FullAdder_17_io_s),
    .io_co(FullAdder_17_io_co)
  );
  FullAdder FullAdder_18 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_18_io_a),
    .io_b(FullAdder_18_io_b),
    .io_ci(FullAdder_18_io_ci),
    .io_s(FullAdder_18_io_s),
    .io_co(FullAdder_18_io_co)
  );
  FullAdder FullAdder_19 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_19_io_a),
    .io_b(FullAdder_19_io_b),
    .io_ci(FullAdder_19_io_ci),
    .io_s(FullAdder_19_io_s),
    .io_co(FullAdder_19_io_co)
  );
  FullAdder FullAdder_20 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_20_io_a),
    .io_b(FullAdder_20_io_b),
    .io_ci(FullAdder_20_io_ci),
    .io_s(FullAdder_20_io_s),
    .io_co(FullAdder_20_io_co)
  );
  FullAdder FullAdder_21 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_21_io_a),
    .io_b(FullAdder_21_io_b),
    .io_ci(FullAdder_21_io_ci),
    .io_s(FullAdder_21_io_s),
    .io_co(FullAdder_21_io_co)
  );
  FullAdder FullAdder_22 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_22_io_a),
    .io_b(FullAdder_22_io_b),
    .io_ci(FullAdder_22_io_ci),
    .io_s(FullAdder_22_io_s),
    .io_co(FullAdder_22_io_co)
  );
  FullAdder FullAdder_23 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_23_io_a),
    .io_b(FullAdder_23_io_b),
    .io_ci(FullAdder_23_io_ci),
    .io_s(FullAdder_23_io_s),
    .io_co(FullAdder_23_io_co)
  );
  FullAdder FullAdder_24 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_24_io_a),
    .io_b(FullAdder_24_io_b),
    .io_ci(FullAdder_24_io_ci),
    .io_s(FullAdder_24_io_s),
    .io_co(FullAdder_24_io_co)
  );
  FullAdder FullAdder_25 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_25_io_a),
    .io_b(FullAdder_25_io_b),
    .io_ci(FullAdder_25_io_ci),
    .io_s(FullAdder_25_io_s),
    .io_co(FullAdder_25_io_co)
  );
  FullAdder FullAdder_26 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_26_io_a),
    .io_b(FullAdder_26_io_b),
    .io_ci(FullAdder_26_io_ci),
    .io_s(FullAdder_26_io_s),
    .io_co(FullAdder_26_io_co)
  );
  FullAdder FullAdder_27 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_27_io_a),
    .io_b(FullAdder_27_io_b),
    .io_ci(FullAdder_27_io_ci),
    .io_s(FullAdder_27_io_s),
    .io_co(FullAdder_27_io_co)
  );
  FullAdder FullAdder_28 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_28_io_a),
    .io_b(FullAdder_28_io_b),
    .io_ci(FullAdder_28_io_ci),
    .io_s(FullAdder_28_io_s),
    .io_co(FullAdder_28_io_co)
  );
  HalfAdder HalfAdder_4 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_4_io_a),
    .io_b(HalfAdder_4_io_b),
    .io_s(HalfAdder_4_io_s),
    .io_co(HalfAdder_4_io_co)
  );
  FullAdder FullAdder_29 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_29_io_a),
    .io_b(FullAdder_29_io_b),
    .io_ci(FullAdder_29_io_ci),
    .io_s(FullAdder_29_io_s),
    .io_co(FullAdder_29_io_co)
  );
  FullAdder FullAdder_30 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_30_io_a),
    .io_b(FullAdder_30_io_b),
    .io_ci(FullAdder_30_io_ci),
    .io_s(FullAdder_30_io_s),
    .io_co(FullAdder_30_io_co)
  );
  FullAdder FullAdder_31 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_31_io_a),
    .io_b(FullAdder_31_io_b),
    .io_ci(FullAdder_31_io_ci),
    .io_s(FullAdder_31_io_s),
    .io_co(FullAdder_31_io_co)
  );
  FullAdder FullAdder_32 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_32_io_a),
    .io_b(FullAdder_32_io_b),
    .io_ci(FullAdder_32_io_ci),
    .io_s(FullAdder_32_io_s),
    .io_co(FullAdder_32_io_co)
  );
  FullAdder FullAdder_33 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_33_io_a),
    .io_b(FullAdder_33_io_b),
    .io_ci(FullAdder_33_io_ci),
    .io_s(FullAdder_33_io_s),
    .io_co(FullAdder_33_io_co)
  );
  FullAdder FullAdder_34 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_34_io_a),
    .io_b(FullAdder_34_io_b),
    .io_ci(FullAdder_34_io_ci),
    .io_s(FullAdder_34_io_s),
    .io_co(FullAdder_34_io_co)
  );
  FullAdder FullAdder_35 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_35_io_a),
    .io_b(FullAdder_35_io_b),
    .io_ci(FullAdder_35_io_ci),
    .io_s(FullAdder_35_io_s),
    .io_co(FullAdder_35_io_co)
  );
  FullAdder FullAdder_36 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_36_io_a),
    .io_b(FullAdder_36_io_b),
    .io_ci(FullAdder_36_io_ci),
    .io_s(FullAdder_36_io_s),
    .io_co(FullAdder_36_io_co)
  );
  FullAdder FullAdder_37 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_37_io_a),
    .io_b(FullAdder_37_io_b),
    .io_ci(FullAdder_37_io_ci),
    .io_s(FullAdder_37_io_s),
    .io_co(FullAdder_37_io_co)
  );
  FullAdder FullAdder_38 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_38_io_a),
    .io_b(FullAdder_38_io_b),
    .io_ci(FullAdder_38_io_ci),
    .io_s(FullAdder_38_io_s),
    .io_co(FullAdder_38_io_co)
  );
  FullAdder FullAdder_39 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_39_io_a),
    .io_b(FullAdder_39_io_b),
    .io_ci(FullAdder_39_io_ci),
    .io_s(FullAdder_39_io_s),
    .io_co(FullAdder_39_io_co)
  );
  FullAdder FullAdder_40 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_40_io_a),
    .io_b(FullAdder_40_io_b),
    .io_ci(FullAdder_40_io_ci),
    .io_s(FullAdder_40_io_s),
    .io_co(FullAdder_40_io_co)
  );
  FullAdder FullAdder_41 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_41_io_a),
    .io_b(FullAdder_41_io_b),
    .io_ci(FullAdder_41_io_ci),
    .io_s(FullAdder_41_io_s),
    .io_co(FullAdder_41_io_co)
  );
  FullAdder FullAdder_42 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_42_io_a),
    .io_b(FullAdder_42_io_b),
    .io_ci(FullAdder_42_io_ci),
    .io_s(FullAdder_42_io_s),
    .io_co(FullAdder_42_io_co)
  );
  FullAdder FullAdder_43 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_43_io_a),
    .io_b(FullAdder_43_io_b),
    .io_ci(FullAdder_43_io_ci),
    .io_s(FullAdder_43_io_s),
    .io_co(FullAdder_43_io_co)
  );
  HalfAdder HalfAdder_5 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_5_io_a),
    .io_b(HalfAdder_5_io_b),
    .io_s(HalfAdder_5_io_s),
    .io_co(HalfAdder_5_io_co)
  );
  FullAdder FullAdder_44 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_44_io_a),
    .io_b(FullAdder_44_io_b),
    .io_ci(FullAdder_44_io_ci),
    .io_s(FullAdder_44_io_s),
    .io_co(FullAdder_44_io_co)
  );
  FullAdder FullAdder_45 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_45_io_a),
    .io_b(FullAdder_45_io_b),
    .io_ci(FullAdder_45_io_ci),
    .io_s(FullAdder_45_io_s),
    .io_co(FullAdder_45_io_co)
  );
  FullAdder FullAdder_46 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_46_io_a),
    .io_b(FullAdder_46_io_b),
    .io_ci(FullAdder_46_io_ci),
    .io_s(FullAdder_46_io_s),
    .io_co(FullAdder_46_io_co)
  );
  FullAdder FullAdder_47 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_47_io_a),
    .io_b(FullAdder_47_io_b),
    .io_ci(FullAdder_47_io_ci),
    .io_s(FullAdder_47_io_s),
    .io_co(FullAdder_47_io_co)
  );
  FullAdder FullAdder_48 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_48_io_a),
    .io_b(FullAdder_48_io_b),
    .io_ci(FullAdder_48_io_ci),
    .io_s(FullAdder_48_io_s),
    .io_co(FullAdder_48_io_co)
  );
  FullAdder FullAdder_49 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_49_io_a),
    .io_b(FullAdder_49_io_b),
    .io_ci(FullAdder_49_io_ci),
    .io_s(FullAdder_49_io_s),
    .io_co(FullAdder_49_io_co)
  );
  FullAdder FullAdder_50 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_50_io_a),
    .io_b(FullAdder_50_io_b),
    .io_ci(FullAdder_50_io_ci),
    .io_s(FullAdder_50_io_s),
    .io_co(FullAdder_50_io_co)
  );
  FullAdder FullAdder_51 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_51_io_a),
    .io_b(FullAdder_51_io_b),
    .io_ci(FullAdder_51_io_ci),
    .io_s(FullAdder_51_io_s),
    .io_co(FullAdder_51_io_co)
  );
  FullAdder FullAdder_52 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_52_io_a),
    .io_b(FullAdder_52_io_b),
    .io_ci(FullAdder_52_io_ci),
    .io_s(FullAdder_52_io_s),
    .io_co(FullAdder_52_io_co)
  );
  FullAdder FullAdder_53 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_53_io_a),
    .io_b(FullAdder_53_io_b),
    .io_ci(FullAdder_53_io_ci),
    .io_s(FullAdder_53_io_s),
    .io_co(FullAdder_53_io_co)
  );
  FullAdder FullAdder_54 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_54_io_a),
    .io_b(FullAdder_54_io_b),
    .io_ci(FullAdder_54_io_ci),
    .io_s(FullAdder_54_io_s),
    .io_co(FullAdder_54_io_co)
  );
  FullAdder FullAdder_55 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_55_io_a),
    .io_b(FullAdder_55_io_b),
    .io_ci(FullAdder_55_io_ci),
    .io_s(FullAdder_55_io_s),
    .io_co(FullAdder_55_io_co)
  );
  FullAdder FullAdder_56 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_56_io_a),
    .io_b(FullAdder_56_io_b),
    .io_ci(FullAdder_56_io_ci),
    .io_s(FullAdder_56_io_s),
    .io_co(FullAdder_56_io_co)
  );
  FullAdder FullAdder_57 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_57_io_a),
    .io_b(FullAdder_57_io_b),
    .io_ci(FullAdder_57_io_ci),
    .io_s(FullAdder_57_io_s),
    .io_co(FullAdder_57_io_co)
  );
  FullAdder FullAdder_58 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_58_io_a),
    .io_b(FullAdder_58_io_b),
    .io_ci(FullAdder_58_io_ci),
    .io_s(FullAdder_58_io_s),
    .io_co(FullAdder_58_io_co)
  );
  FullAdder FullAdder_59 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_59_io_a),
    .io_b(FullAdder_59_io_b),
    .io_ci(FullAdder_59_io_ci),
    .io_s(FullAdder_59_io_s),
    .io_co(FullAdder_59_io_co)
  );
  FullAdder FullAdder_60 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_60_io_a),
    .io_b(FullAdder_60_io_b),
    .io_ci(FullAdder_60_io_ci),
    .io_s(FullAdder_60_io_s),
    .io_co(FullAdder_60_io_co)
  );
  FullAdder FullAdder_61 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_61_io_a),
    .io_b(FullAdder_61_io_b),
    .io_ci(FullAdder_61_io_ci),
    .io_s(FullAdder_61_io_s),
    .io_co(FullAdder_61_io_co)
  );
  FullAdder FullAdder_62 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_62_io_a),
    .io_b(FullAdder_62_io_b),
    .io_ci(FullAdder_62_io_ci),
    .io_s(FullAdder_62_io_s),
    .io_co(FullAdder_62_io_co)
  );
  FullAdder FullAdder_63 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_63_io_a),
    .io_b(FullAdder_63_io_b),
    .io_ci(FullAdder_63_io_ci),
    .io_s(FullAdder_63_io_s),
    .io_co(FullAdder_63_io_co)
  );
  FullAdder FullAdder_64 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_64_io_a),
    .io_b(FullAdder_64_io_b),
    .io_ci(FullAdder_64_io_ci),
    .io_s(FullAdder_64_io_s),
    .io_co(FullAdder_64_io_co)
  );
  FullAdder FullAdder_65 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_65_io_a),
    .io_b(FullAdder_65_io_b),
    .io_ci(FullAdder_65_io_ci),
    .io_s(FullAdder_65_io_s),
    .io_co(FullAdder_65_io_co)
  );
  FullAdder FullAdder_66 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_66_io_a),
    .io_b(FullAdder_66_io_b),
    .io_ci(FullAdder_66_io_ci),
    .io_s(FullAdder_66_io_s),
    .io_co(FullAdder_66_io_co)
  );
  FullAdder FullAdder_67 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_67_io_a),
    .io_b(FullAdder_67_io_b),
    .io_ci(FullAdder_67_io_ci),
    .io_s(FullAdder_67_io_s),
    .io_co(FullAdder_67_io_co)
  );
  FullAdder FullAdder_68 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_68_io_a),
    .io_b(FullAdder_68_io_b),
    .io_ci(FullAdder_68_io_ci),
    .io_s(FullAdder_68_io_s),
    .io_co(FullAdder_68_io_co)
  );
  FullAdder FullAdder_69 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_69_io_a),
    .io_b(FullAdder_69_io_b),
    .io_ci(FullAdder_69_io_ci),
    .io_s(FullAdder_69_io_s),
    .io_co(FullAdder_69_io_co)
  );
  FullAdder FullAdder_70 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_70_io_a),
    .io_b(FullAdder_70_io_b),
    .io_ci(FullAdder_70_io_ci),
    .io_s(FullAdder_70_io_s),
    .io_co(FullAdder_70_io_co)
  );
  FullAdder FullAdder_71 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_71_io_a),
    .io_b(FullAdder_71_io_b),
    .io_ci(FullAdder_71_io_ci),
    .io_s(FullAdder_71_io_s),
    .io_co(FullAdder_71_io_co)
  );
  FullAdder FullAdder_72 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_72_io_a),
    .io_b(FullAdder_72_io_b),
    .io_ci(FullAdder_72_io_ci),
    .io_s(FullAdder_72_io_s),
    .io_co(FullAdder_72_io_co)
  );
  FullAdder FullAdder_73 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_73_io_a),
    .io_b(FullAdder_73_io_b),
    .io_ci(FullAdder_73_io_ci),
    .io_s(FullAdder_73_io_s),
    .io_co(FullAdder_73_io_co)
  );
  FullAdder FullAdder_74 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_74_io_a),
    .io_b(FullAdder_74_io_b),
    .io_ci(FullAdder_74_io_ci),
    .io_s(FullAdder_74_io_s),
    .io_co(FullAdder_74_io_co)
  );
  FullAdder FullAdder_75 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_75_io_a),
    .io_b(FullAdder_75_io_b),
    .io_ci(FullAdder_75_io_ci),
    .io_s(FullAdder_75_io_s),
    .io_co(FullAdder_75_io_co)
  );
  FullAdder FullAdder_76 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_76_io_a),
    .io_b(FullAdder_76_io_b),
    .io_ci(FullAdder_76_io_ci),
    .io_s(FullAdder_76_io_s),
    .io_co(FullAdder_76_io_co)
  );
  FullAdder FullAdder_77 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_77_io_a),
    .io_b(FullAdder_77_io_b),
    .io_ci(FullAdder_77_io_ci),
    .io_s(FullAdder_77_io_s),
    .io_co(FullAdder_77_io_co)
  );
  FullAdder FullAdder_78 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_78_io_a),
    .io_b(FullAdder_78_io_b),
    .io_ci(FullAdder_78_io_ci),
    .io_s(FullAdder_78_io_s),
    .io_co(FullAdder_78_io_co)
  );
  FullAdder FullAdder_79 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_79_io_a),
    .io_b(FullAdder_79_io_b),
    .io_ci(FullAdder_79_io_ci),
    .io_s(FullAdder_79_io_s),
    .io_co(FullAdder_79_io_co)
  );
  FullAdder FullAdder_80 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_80_io_a),
    .io_b(FullAdder_80_io_b),
    .io_ci(FullAdder_80_io_ci),
    .io_s(FullAdder_80_io_s),
    .io_co(FullAdder_80_io_co)
  );
  FullAdder FullAdder_81 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_81_io_a),
    .io_b(FullAdder_81_io_b),
    .io_ci(FullAdder_81_io_ci),
    .io_s(FullAdder_81_io_s),
    .io_co(FullAdder_81_io_co)
  );
  FullAdder FullAdder_82 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_82_io_a),
    .io_b(FullAdder_82_io_b),
    .io_ci(FullAdder_82_io_ci),
    .io_s(FullAdder_82_io_s),
    .io_co(FullAdder_82_io_co)
  );
  HalfAdder HalfAdder_6 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_6_io_a),
    .io_b(HalfAdder_6_io_b),
    .io_s(HalfAdder_6_io_s),
    .io_co(HalfAdder_6_io_co)
  );
  FullAdder FullAdder_83 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_83_io_a),
    .io_b(FullAdder_83_io_b),
    .io_ci(FullAdder_83_io_ci),
    .io_s(FullAdder_83_io_s),
    .io_co(FullAdder_83_io_co)
  );
  FullAdder FullAdder_84 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_84_io_a),
    .io_b(FullAdder_84_io_b),
    .io_ci(FullAdder_84_io_ci),
    .io_s(FullAdder_84_io_s),
    .io_co(FullAdder_84_io_co)
  );
  FullAdder FullAdder_85 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_85_io_a),
    .io_b(FullAdder_85_io_b),
    .io_ci(FullAdder_85_io_ci),
    .io_s(FullAdder_85_io_s),
    .io_co(FullAdder_85_io_co)
  );
  FullAdder FullAdder_86 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_86_io_a),
    .io_b(FullAdder_86_io_b),
    .io_ci(FullAdder_86_io_ci),
    .io_s(FullAdder_86_io_s),
    .io_co(FullAdder_86_io_co)
  );
  FullAdder FullAdder_87 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_87_io_a),
    .io_b(FullAdder_87_io_b),
    .io_ci(FullAdder_87_io_ci),
    .io_s(FullAdder_87_io_s),
    .io_co(FullAdder_87_io_co)
  );
  FullAdder FullAdder_88 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_88_io_a),
    .io_b(FullAdder_88_io_b),
    .io_ci(FullAdder_88_io_ci),
    .io_s(FullAdder_88_io_s),
    .io_co(FullAdder_88_io_co)
  );
  FullAdder FullAdder_89 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_89_io_a),
    .io_b(FullAdder_89_io_b),
    .io_ci(FullAdder_89_io_ci),
    .io_s(FullAdder_89_io_s),
    .io_co(FullAdder_89_io_co)
  );
  FullAdder FullAdder_90 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_90_io_a),
    .io_b(FullAdder_90_io_b),
    .io_ci(FullAdder_90_io_ci),
    .io_s(FullAdder_90_io_s),
    .io_co(FullAdder_90_io_co)
  );
  FullAdder FullAdder_91 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_91_io_a),
    .io_b(FullAdder_91_io_b),
    .io_ci(FullAdder_91_io_ci),
    .io_s(FullAdder_91_io_s),
    .io_co(FullAdder_91_io_co)
  );
  FullAdder FullAdder_92 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_92_io_a),
    .io_b(FullAdder_92_io_b),
    .io_ci(FullAdder_92_io_ci),
    .io_s(FullAdder_92_io_s),
    .io_co(FullAdder_92_io_co)
  );
  FullAdder FullAdder_93 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_93_io_a),
    .io_b(FullAdder_93_io_b),
    .io_ci(FullAdder_93_io_ci),
    .io_s(FullAdder_93_io_s),
    .io_co(FullAdder_93_io_co)
  );
  FullAdder FullAdder_94 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_94_io_a),
    .io_b(FullAdder_94_io_b),
    .io_ci(FullAdder_94_io_ci),
    .io_s(FullAdder_94_io_s),
    .io_co(FullAdder_94_io_co)
  );
  FullAdder FullAdder_95 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_95_io_a),
    .io_b(FullAdder_95_io_b),
    .io_ci(FullAdder_95_io_ci),
    .io_s(FullAdder_95_io_s),
    .io_co(FullAdder_95_io_co)
  );
  FullAdder FullAdder_96 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_96_io_a),
    .io_b(FullAdder_96_io_b),
    .io_ci(FullAdder_96_io_ci),
    .io_s(FullAdder_96_io_s),
    .io_co(FullAdder_96_io_co)
  );
  FullAdder FullAdder_97 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_97_io_a),
    .io_b(FullAdder_97_io_b),
    .io_ci(FullAdder_97_io_ci),
    .io_s(FullAdder_97_io_s),
    .io_co(FullAdder_97_io_co)
  );
  FullAdder FullAdder_98 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_98_io_a),
    .io_b(FullAdder_98_io_b),
    .io_ci(FullAdder_98_io_ci),
    .io_s(FullAdder_98_io_s),
    .io_co(FullAdder_98_io_co)
  );
  FullAdder FullAdder_99 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_99_io_a),
    .io_b(FullAdder_99_io_b),
    .io_ci(FullAdder_99_io_ci),
    .io_s(FullAdder_99_io_s),
    .io_co(FullAdder_99_io_co)
  );
  FullAdder FullAdder_100 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_100_io_a),
    .io_b(FullAdder_100_io_b),
    .io_ci(FullAdder_100_io_ci),
    .io_s(FullAdder_100_io_s),
    .io_co(FullAdder_100_io_co)
  );
  FullAdder FullAdder_101 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_101_io_a),
    .io_b(FullAdder_101_io_b),
    .io_ci(FullAdder_101_io_ci),
    .io_s(FullAdder_101_io_s),
    .io_co(FullAdder_101_io_co)
  );
  FullAdder FullAdder_102 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_102_io_a),
    .io_b(FullAdder_102_io_b),
    .io_ci(FullAdder_102_io_ci),
    .io_s(FullAdder_102_io_s),
    .io_co(FullAdder_102_io_co)
  );
  FullAdder FullAdder_103 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_103_io_a),
    .io_b(FullAdder_103_io_b),
    .io_ci(FullAdder_103_io_ci),
    .io_s(FullAdder_103_io_s),
    .io_co(FullAdder_103_io_co)
  );
  FullAdder FullAdder_104 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_104_io_a),
    .io_b(FullAdder_104_io_b),
    .io_ci(FullAdder_104_io_ci),
    .io_s(FullAdder_104_io_s),
    .io_co(FullAdder_104_io_co)
  );
  FullAdder FullAdder_105 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_105_io_a),
    .io_b(FullAdder_105_io_b),
    .io_ci(FullAdder_105_io_ci),
    .io_s(FullAdder_105_io_s),
    .io_co(FullAdder_105_io_co)
  );
  FullAdder FullAdder_106 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_106_io_a),
    .io_b(FullAdder_106_io_b),
    .io_ci(FullAdder_106_io_ci),
    .io_s(FullAdder_106_io_s),
    .io_co(FullAdder_106_io_co)
  );
  FullAdder FullAdder_107 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_107_io_a),
    .io_b(FullAdder_107_io_b),
    .io_ci(FullAdder_107_io_ci),
    .io_s(FullAdder_107_io_s),
    .io_co(FullAdder_107_io_co)
  );
  FullAdder FullAdder_108 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_108_io_a),
    .io_b(FullAdder_108_io_b),
    .io_ci(FullAdder_108_io_ci),
    .io_s(FullAdder_108_io_s),
    .io_co(FullAdder_108_io_co)
  );
  FullAdder FullAdder_109 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_109_io_a),
    .io_b(FullAdder_109_io_b),
    .io_ci(FullAdder_109_io_ci),
    .io_s(FullAdder_109_io_s),
    .io_co(FullAdder_109_io_co)
  );
  FullAdder FullAdder_110 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_110_io_a),
    .io_b(FullAdder_110_io_b),
    .io_ci(FullAdder_110_io_ci),
    .io_s(FullAdder_110_io_s),
    .io_co(FullAdder_110_io_co)
  );
  FullAdder FullAdder_111 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_111_io_a),
    .io_b(FullAdder_111_io_b),
    .io_ci(FullAdder_111_io_ci),
    .io_s(FullAdder_111_io_s),
    .io_co(FullAdder_111_io_co)
  );
  FullAdder FullAdder_112 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_112_io_a),
    .io_b(FullAdder_112_io_b),
    .io_ci(FullAdder_112_io_ci),
    .io_s(FullAdder_112_io_s),
    .io_co(FullAdder_112_io_co)
  );
  FullAdder FullAdder_113 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_113_io_a),
    .io_b(FullAdder_113_io_b),
    .io_ci(FullAdder_113_io_ci),
    .io_s(FullAdder_113_io_s),
    .io_co(FullAdder_113_io_co)
  );
  FullAdder FullAdder_114 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_114_io_a),
    .io_b(FullAdder_114_io_b),
    .io_ci(FullAdder_114_io_ci),
    .io_s(FullAdder_114_io_s),
    .io_co(FullAdder_114_io_co)
  );
  FullAdder FullAdder_115 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_115_io_a),
    .io_b(FullAdder_115_io_b),
    .io_ci(FullAdder_115_io_ci),
    .io_s(FullAdder_115_io_s),
    .io_co(FullAdder_115_io_co)
  );
  FullAdder FullAdder_116 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_116_io_a),
    .io_b(FullAdder_116_io_b),
    .io_ci(FullAdder_116_io_ci),
    .io_s(FullAdder_116_io_s),
    .io_co(FullAdder_116_io_co)
  );
  FullAdder FullAdder_117 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_117_io_a),
    .io_b(FullAdder_117_io_b),
    .io_ci(FullAdder_117_io_ci),
    .io_s(FullAdder_117_io_s),
    .io_co(FullAdder_117_io_co)
  );
  FullAdder FullAdder_118 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_118_io_a),
    .io_b(FullAdder_118_io_b),
    .io_ci(FullAdder_118_io_ci),
    .io_s(FullAdder_118_io_s),
    .io_co(FullAdder_118_io_co)
  );
  FullAdder FullAdder_119 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_119_io_a),
    .io_b(FullAdder_119_io_b),
    .io_ci(FullAdder_119_io_ci),
    .io_s(FullAdder_119_io_s),
    .io_co(FullAdder_119_io_co)
  );
  FullAdder FullAdder_120 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_120_io_a),
    .io_b(FullAdder_120_io_b),
    .io_ci(FullAdder_120_io_ci),
    .io_s(FullAdder_120_io_s),
    .io_co(FullAdder_120_io_co)
  );
  FullAdder FullAdder_121 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_121_io_a),
    .io_b(FullAdder_121_io_b),
    .io_ci(FullAdder_121_io_ci),
    .io_s(FullAdder_121_io_s),
    .io_co(FullAdder_121_io_co)
  );
  FullAdder FullAdder_122 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_122_io_a),
    .io_b(FullAdder_122_io_b),
    .io_ci(FullAdder_122_io_ci),
    .io_s(FullAdder_122_io_s),
    .io_co(FullAdder_122_io_co)
  );
  FullAdder FullAdder_123 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_123_io_a),
    .io_b(FullAdder_123_io_b),
    .io_ci(FullAdder_123_io_ci),
    .io_s(FullAdder_123_io_s),
    .io_co(FullAdder_123_io_co)
  );
  FullAdder FullAdder_124 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_124_io_a),
    .io_b(FullAdder_124_io_b),
    .io_ci(FullAdder_124_io_ci),
    .io_s(FullAdder_124_io_s),
    .io_co(FullAdder_124_io_co)
  );
  FullAdder FullAdder_125 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_125_io_a),
    .io_b(FullAdder_125_io_b),
    .io_ci(FullAdder_125_io_ci),
    .io_s(FullAdder_125_io_s),
    .io_co(FullAdder_125_io_co)
  );
  FullAdder FullAdder_126 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_126_io_a),
    .io_b(FullAdder_126_io_b),
    .io_ci(FullAdder_126_io_ci),
    .io_s(FullAdder_126_io_s),
    .io_co(FullAdder_126_io_co)
  );
  FullAdder FullAdder_127 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_127_io_a),
    .io_b(FullAdder_127_io_b),
    .io_ci(FullAdder_127_io_ci),
    .io_s(FullAdder_127_io_s),
    .io_co(FullAdder_127_io_co)
  );
  FullAdder FullAdder_128 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_128_io_a),
    .io_b(FullAdder_128_io_b),
    .io_ci(FullAdder_128_io_ci),
    .io_s(FullAdder_128_io_s),
    .io_co(FullAdder_128_io_co)
  );
  FullAdder FullAdder_129 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_129_io_a),
    .io_b(FullAdder_129_io_b),
    .io_ci(FullAdder_129_io_ci),
    .io_s(FullAdder_129_io_s),
    .io_co(FullAdder_129_io_co)
  );
  FullAdder FullAdder_130 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_130_io_a),
    .io_b(FullAdder_130_io_b),
    .io_ci(FullAdder_130_io_ci),
    .io_s(FullAdder_130_io_s),
    .io_co(FullAdder_130_io_co)
  );
  FullAdder FullAdder_131 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_131_io_a),
    .io_b(FullAdder_131_io_b),
    .io_ci(FullAdder_131_io_ci),
    .io_s(FullAdder_131_io_s),
    .io_co(FullAdder_131_io_co)
  );
  FullAdder FullAdder_132 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_132_io_a),
    .io_b(FullAdder_132_io_b),
    .io_ci(FullAdder_132_io_ci),
    .io_s(FullAdder_132_io_s),
    .io_co(FullAdder_132_io_co)
  );
  FullAdder FullAdder_133 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_133_io_a),
    .io_b(FullAdder_133_io_b),
    .io_ci(FullAdder_133_io_ci),
    .io_s(FullAdder_133_io_s),
    .io_co(FullAdder_133_io_co)
  );
  HalfAdder HalfAdder_7 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_7_io_a),
    .io_b(HalfAdder_7_io_b),
    .io_s(HalfAdder_7_io_s),
    .io_co(HalfAdder_7_io_co)
  );
  FullAdder FullAdder_134 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_134_io_a),
    .io_b(FullAdder_134_io_b),
    .io_ci(FullAdder_134_io_ci),
    .io_s(FullAdder_134_io_s),
    .io_co(FullAdder_134_io_co)
  );
  FullAdder FullAdder_135 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_135_io_a),
    .io_b(FullAdder_135_io_b),
    .io_ci(FullAdder_135_io_ci),
    .io_s(FullAdder_135_io_s),
    .io_co(FullAdder_135_io_co)
  );
  FullAdder FullAdder_136 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_136_io_a),
    .io_b(FullAdder_136_io_b),
    .io_ci(FullAdder_136_io_ci),
    .io_s(FullAdder_136_io_s),
    .io_co(FullAdder_136_io_co)
  );
  FullAdder FullAdder_137 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_137_io_a),
    .io_b(FullAdder_137_io_b),
    .io_ci(FullAdder_137_io_ci),
    .io_s(FullAdder_137_io_s),
    .io_co(FullAdder_137_io_co)
  );
  FullAdder FullAdder_138 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_138_io_a),
    .io_b(FullAdder_138_io_b),
    .io_ci(FullAdder_138_io_ci),
    .io_s(FullAdder_138_io_s),
    .io_co(FullAdder_138_io_co)
  );
  FullAdder FullAdder_139 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_139_io_a),
    .io_b(FullAdder_139_io_b),
    .io_ci(FullAdder_139_io_ci),
    .io_s(FullAdder_139_io_s),
    .io_co(FullAdder_139_io_co)
  );
  FullAdder FullAdder_140 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_140_io_a),
    .io_b(FullAdder_140_io_b),
    .io_ci(FullAdder_140_io_ci),
    .io_s(FullAdder_140_io_s),
    .io_co(FullAdder_140_io_co)
  );
  FullAdder FullAdder_141 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_141_io_a),
    .io_b(FullAdder_141_io_b),
    .io_ci(FullAdder_141_io_ci),
    .io_s(FullAdder_141_io_s),
    .io_co(FullAdder_141_io_co)
  );
  FullAdder FullAdder_142 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_142_io_a),
    .io_b(FullAdder_142_io_b),
    .io_ci(FullAdder_142_io_ci),
    .io_s(FullAdder_142_io_s),
    .io_co(FullAdder_142_io_co)
  );
  FullAdder FullAdder_143 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_143_io_a),
    .io_b(FullAdder_143_io_b),
    .io_ci(FullAdder_143_io_ci),
    .io_s(FullAdder_143_io_s),
    .io_co(FullAdder_143_io_co)
  );
  FullAdder FullAdder_144 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_144_io_a),
    .io_b(FullAdder_144_io_b),
    .io_ci(FullAdder_144_io_ci),
    .io_s(FullAdder_144_io_s),
    .io_co(FullAdder_144_io_co)
  );
  FullAdder FullAdder_145 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_145_io_a),
    .io_b(FullAdder_145_io_b),
    .io_ci(FullAdder_145_io_ci),
    .io_s(FullAdder_145_io_s),
    .io_co(FullAdder_145_io_co)
  );
  FullAdder FullAdder_146 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_146_io_a),
    .io_b(FullAdder_146_io_b),
    .io_ci(FullAdder_146_io_ci),
    .io_s(FullAdder_146_io_s),
    .io_co(FullAdder_146_io_co)
  );
  FullAdder FullAdder_147 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_147_io_a),
    .io_b(FullAdder_147_io_b),
    .io_ci(FullAdder_147_io_ci),
    .io_s(FullAdder_147_io_s),
    .io_co(FullAdder_147_io_co)
  );
  FullAdder FullAdder_148 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_148_io_a),
    .io_b(FullAdder_148_io_b),
    .io_ci(FullAdder_148_io_ci),
    .io_s(FullAdder_148_io_s),
    .io_co(FullAdder_148_io_co)
  );
  FullAdder FullAdder_149 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_149_io_a),
    .io_b(FullAdder_149_io_b),
    .io_ci(FullAdder_149_io_ci),
    .io_s(FullAdder_149_io_s),
    .io_co(FullAdder_149_io_co)
  );
  FullAdder FullAdder_150 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_150_io_a),
    .io_b(FullAdder_150_io_b),
    .io_ci(FullAdder_150_io_ci),
    .io_s(FullAdder_150_io_s),
    .io_co(FullAdder_150_io_co)
  );
  FullAdder FullAdder_151 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_151_io_a),
    .io_b(FullAdder_151_io_b),
    .io_ci(FullAdder_151_io_ci),
    .io_s(FullAdder_151_io_s),
    .io_co(FullAdder_151_io_co)
  );
  FullAdder FullAdder_152 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_152_io_a),
    .io_b(FullAdder_152_io_b),
    .io_ci(FullAdder_152_io_ci),
    .io_s(FullAdder_152_io_s),
    .io_co(FullAdder_152_io_co)
  );
  FullAdder FullAdder_153 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_153_io_a),
    .io_b(FullAdder_153_io_b),
    .io_ci(FullAdder_153_io_ci),
    .io_s(FullAdder_153_io_s),
    .io_co(FullAdder_153_io_co)
  );
  FullAdder FullAdder_154 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_154_io_a),
    .io_b(FullAdder_154_io_b),
    .io_ci(FullAdder_154_io_ci),
    .io_s(FullAdder_154_io_s),
    .io_co(FullAdder_154_io_co)
  );
  FullAdder FullAdder_155 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_155_io_a),
    .io_b(FullAdder_155_io_b),
    .io_ci(FullAdder_155_io_ci),
    .io_s(FullAdder_155_io_s),
    .io_co(FullAdder_155_io_co)
  );
  FullAdder FullAdder_156 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_156_io_a),
    .io_b(FullAdder_156_io_b),
    .io_ci(FullAdder_156_io_ci),
    .io_s(FullAdder_156_io_s),
    .io_co(FullAdder_156_io_co)
  );
  FullAdder FullAdder_157 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_157_io_a),
    .io_b(FullAdder_157_io_b),
    .io_ci(FullAdder_157_io_ci),
    .io_s(FullAdder_157_io_s),
    .io_co(FullAdder_157_io_co)
  );
  FullAdder FullAdder_158 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_158_io_a),
    .io_b(FullAdder_158_io_b),
    .io_ci(FullAdder_158_io_ci),
    .io_s(FullAdder_158_io_s),
    .io_co(FullAdder_158_io_co)
  );
  FullAdder FullAdder_159 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_159_io_a),
    .io_b(FullAdder_159_io_b),
    .io_ci(FullAdder_159_io_ci),
    .io_s(FullAdder_159_io_s),
    .io_co(FullAdder_159_io_co)
  );
  FullAdder FullAdder_160 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_160_io_a),
    .io_b(FullAdder_160_io_b),
    .io_ci(FullAdder_160_io_ci),
    .io_s(FullAdder_160_io_s),
    .io_co(FullAdder_160_io_co)
  );
  FullAdder FullAdder_161 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_161_io_a),
    .io_b(FullAdder_161_io_b),
    .io_ci(FullAdder_161_io_ci),
    .io_s(FullAdder_161_io_s),
    .io_co(FullAdder_161_io_co)
  );
  FullAdder FullAdder_162 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_162_io_a),
    .io_b(FullAdder_162_io_b),
    .io_ci(FullAdder_162_io_ci),
    .io_s(FullAdder_162_io_s),
    .io_co(FullAdder_162_io_co)
  );
  FullAdder FullAdder_163 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_163_io_a),
    .io_b(FullAdder_163_io_b),
    .io_ci(FullAdder_163_io_ci),
    .io_s(FullAdder_163_io_s),
    .io_co(FullAdder_163_io_co)
  );
  FullAdder FullAdder_164 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_164_io_a),
    .io_b(FullAdder_164_io_b),
    .io_ci(FullAdder_164_io_ci),
    .io_s(FullAdder_164_io_s),
    .io_co(FullAdder_164_io_co)
  );
  FullAdder FullAdder_165 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_165_io_a),
    .io_b(FullAdder_165_io_b),
    .io_ci(FullAdder_165_io_ci),
    .io_s(FullAdder_165_io_s),
    .io_co(FullAdder_165_io_co)
  );
  FullAdder FullAdder_166 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_166_io_a),
    .io_b(FullAdder_166_io_b),
    .io_ci(FullAdder_166_io_ci),
    .io_s(FullAdder_166_io_s),
    .io_co(FullAdder_166_io_co)
  );
  FullAdder FullAdder_167 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_167_io_a),
    .io_b(FullAdder_167_io_b),
    .io_ci(FullAdder_167_io_ci),
    .io_s(FullAdder_167_io_s),
    .io_co(FullAdder_167_io_co)
  );
  FullAdder FullAdder_168 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_168_io_a),
    .io_b(FullAdder_168_io_b),
    .io_ci(FullAdder_168_io_ci),
    .io_s(FullAdder_168_io_s),
    .io_co(FullAdder_168_io_co)
  );
  FullAdder FullAdder_169 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_169_io_a),
    .io_b(FullAdder_169_io_b),
    .io_ci(FullAdder_169_io_ci),
    .io_s(FullAdder_169_io_s),
    .io_co(FullAdder_169_io_co)
  );
  FullAdder FullAdder_170 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_170_io_a),
    .io_b(FullAdder_170_io_b),
    .io_ci(FullAdder_170_io_ci),
    .io_s(FullAdder_170_io_s),
    .io_co(FullAdder_170_io_co)
  );
  FullAdder FullAdder_171 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_171_io_a),
    .io_b(FullAdder_171_io_b),
    .io_ci(FullAdder_171_io_ci),
    .io_s(FullAdder_171_io_s),
    .io_co(FullAdder_171_io_co)
  );
  FullAdder FullAdder_172 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_172_io_a),
    .io_b(FullAdder_172_io_b),
    .io_ci(FullAdder_172_io_ci),
    .io_s(FullAdder_172_io_s),
    .io_co(FullAdder_172_io_co)
  );
  FullAdder FullAdder_173 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_173_io_a),
    .io_b(FullAdder_173_io_b),
    .io_ci(FullAdder_173_io_ci),
    .io_s(FullAdder_173_io_s),
    .io_co(FullAdder_173_io_co)
  );
  FullAdder FullAdder_174 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_174_io_a),
    .io_b(FullAdder_174_io_b),
    .io_ci(FullAdder_174_io_ci),
    .io_s(FullAdder_174_io_s),
    .io_co(FullAdder_174_io_co)
  );
  FullAdder FullAdder_175 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_175_io_a),
    .io_b(FullAdder_175_io_b),
    .io_ci(FullAdder_175_io_ci),
    .io_s(FullAdder_175_io_s),
    .io_co(FullAdder_175_io_co)
  );
  FullAdder FullAdder_176 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_176_io_a),
    .io_b(FullAdder_176_io_b),
    .io_ci(FullAdder_176_io_ci),
    .io_s(FullAdder_176_io_s),
    .io_co(FullAdder_176_io_co)
  );
  FullAdder FullAdder_177 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_177_io_a),
    .io_b(FullAdder_177_io_b),
    .io_ci(FullAdder_177_io_ci),
    .io_s(FullAdder_177_io_s),
    .io_co(FullAdder_177_io_co)
  );
  FullAdder FullAdder_178 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_178_io_a),
    .io_b(FullAdder_178_io_b),
    .io_ci(FullAdder_178_io_ci),
    .io_s(FullAdder_178_io_s),
    .io_co(FullAdder_178_io_co)
  );
  FullAdder FullAdder_179 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_179_io_a),
    .io_b(FullAdder_179_io_b),
    .io_ci(FullAdder_179_io_ci),
    .io_s(FullAdder_179_io_s),
    .io_co(FullAdder_179_io_co)
  );
  FullAdder FullAdder_180 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_180_io_a),
    .io_b(FullAdder_180_io_b),
    .io_ci(FullAdder_180_io_ci),
    .io_s(FullAdder_180_io_s),
    .io_co(FullAdder_180_io_co)
  );
  FullAdder FullAdder_181 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_181_io_a),
    .io_b(FullAdder_181_io_b),
    .io_ci(FullAdder_181_io_ci),
    .io_s(FullAdder_181_io_s),
    .io_co(FullAdder_181_io_co)
  );
  FullAdder FullAdder_182 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_182_io_a),
    .io_b(FullAdder_182_io_b),
    .io_ci(FullAdder_182_io_ci),
    .io_s(FullAdder_182_io_s),
    .io_co(FullAdder_182_io_co)
  );
  FullAdder FullAdder_183 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_183_io_a),
    .io_b(FullAdder_183_io_b),
    .io_ci(FullAdder_183_io_ci),
    .io_s(FullAdder_183_io_s),
    .io_co(FullAdder_183_io_co)
  );
  FullAdder FullAdder_184 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_184_io_a),
    .io_b(FullAdder_184_io_b),
    .io_ci(FullAdder_184_io_ci),
    .io_s(FullAdder_184_io_s),
    .io_co(FullAdder_184_io_co)
  );
  FullAdder FullAdder_185 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_185_io_a),
    .io_b(FullAdder_185_io_b),
    .io_ci(FullAdder_185_io_ci),
    .io_s(FullAdder_185_io_s),
    .io_co(FullAdder_185_io_co)
  );
  FullAdder FullAdder_186 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_186_io_a),
    .io_b(FullAdder_186_io_b),
    .io_ci(FullAdder_186_io_ci),
    .io_s(FullAdder_186_io_s),
    .io_co(FullAdder_186_io_co)
  );
  FullAdder FullAdder_187 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_187_io_a),
    .io_b(FullAdder_187_io_b),
    .io_ci(FullAdder_187_io_ci),
    .io_s(FullAdder_187_io_s),
    .io_co(FullAdder_187_io_co)
  );
  FullAdder FullAdder_188 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_188_io_a),
    .io_b(FullAdder_188_io_b),
    .io_ci(FullAdder_188_io_ci),
    .io_s(FullAdder_188_io_s),
    .io_co(FullAdder_188_io_co)
  );
  FullAdder FullAdder_189 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_189_io_a),
    .io_b(FullAdder_189_io_b),
    .io_ci(FullAdder_189_io_ci),
    .io_s(FullAdder_189_io_s),
    .io_co(FullAdder_189_io_co)
  );
  FullAdder FullAdder_190 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_190_io_a),
    .io_b(FullAdder_190_io_b),
    .io_ci(FullAdder_190_io_ci),
    .io_s(FullAdder_190_io_s),
    .io_co(FullAdder_190_io_co)
  );
  FullAdder FullAdder_191 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_191_io_a),
    .io_b(FullAdder_191_io_b),
    .io_ci(FullAdder_191_io_ci),
    .io_s(FullAdder_191_io_s),
    .io_co(FullAdder_191_io_co)
  );
  FullAdder FullAdder_192 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_192_io_a),
    .io_b(FullAdder_192_io_b),
    .io_ci(FullAdder_192_io_ci),
    .io_s(FullAdder_192_io_s),
    .io_co(FullAdder_192_io_co)
  );
  HalfAdder HalfAdder_8 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_8_io_a),
    .io_b(HalfAdder_8_io_b),
    .io_s(HalfAdder_8_io_s),
    .io_co(HalfAdder_8_io_co)
  );
  FullAdder FullAdder_193 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_193_io_a),
    .io_b(FullAdder_193_io_b),
    .io_ci(FullAdder_193_io_ci),
    .io_s(FullAdder_193_io_s),
    .io_co(FullAdder_193_io_co)
  );
  FullAdder FullAdder_194 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_194_io_a),
    .io_b(FullAdder_194_io_b),
    .io_ci(FullAdder_194_io_ci),
    .io_s(FullAdder_194_io_s),
    .io_co(FullAdder_194_io_co)
  );
  FullAdder FullAdder_195 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_195_io_a),
    .io_b(FullAdder_195_io_b),
    .io_ci(FullAdder_195_io_ci),
    .io_s(FullAdder_195_io_s),
    .io_co(FullAdder_195_io_co)
  );
  FullAdder FullAdder_196 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_196_io_a),
    .io_b(FullAdder_196_io_b),
    .io_ci(FullAdder_196_io_ci),
    .io_s(FullAdder_196_io_s),
    .io_co(FullAdder_196_io_co)
  );
  FullAdder FullAdder_197 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_197_io_a),
    .io_b(FullAdder_197_io_b),
    .io_ci(FullAdder_197_io_ci),
    .io_s(FullAdder_197_io_s),
    .io_co(FullAdder_197_io_co)
  );
  FullAdder FullAdder_198 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_198_io_a),
    .io_b(FullAdder_198_io_b),
    .io_ci(FullAdder_198_io_ci),
    .io_s(FullAdder_198_io_s),
    .io_co(FullAdder_198_io_co)
  );
  FullAdder FullAdder_199 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_199_io_a),
    .io_b(FullAdder_199_io_b),
    .io_ci(FullAdder_199_io_ci),
    .io_s(FullAdder_199_io_s),
    .io_co(FullAdder_199_io_co)
  );
  FullAdder FullAdder_200 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_200_io_a),
    .io_b(FullAdder_200_io_b),
    .io_ci(FullAdder_200_io_ci),
    .io_s(FullAdder_200_io_s),
    .io_co(FullAdder_200_io_co)
  );
  FullAdder FullAdder_201 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_201_io_a),
    .io_b(FullAdder_201_io_b),
    .io_ci(FullAdder_201_io_ci),
    .io_s(FullAdder_201_io_s),
    .io_co(FullAdder_201_io_co)
  );
  FullAdder FullAdder_202 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_202_io_a),
    .io_b(FullAdder_202_io_b),
    .io_ci(FullAdder_202_io_ci),
    .io_s(FullAdder_202_io_s),
    .io_co(FullAdder_202_io_co)
  );
  FullAdder FullAdder_203 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_203_io_a),
    .io_b(FullAdder_203_io_b),
    .io_ci(FullAdder_203_io_ci),
    .io_s(FullAdder_203_io_s),
    .io_co(FullAdder_203_io_co)
  );
  FullAdder FullAdder_204 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_204_io_a),
    .io_b(FullAdder_204_io_b),
    .io_ci(FullAdder_204_io_ci),
    .io_s(FullAdder_204_io_s),
    .io_co(FullAdder_204_io_co)
  );
  FullAdder FullAdder_205 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_205_io_a),
    .io_b(FullAdder_205_io_b),
    .io_ci(FullAdder_205_io_ci),
    .io_s(FullAdder_205_io_s),
    .io_co(FullAdder_205_io_co)
  );
  FullAdder FullAdder_206 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_206_io_a),
    .io_b(FullAdder_206_io_b),
    .io_ci(FullAdder_206_io_ci),
    .io_s(FullAdder_206_io_s),
    .io_co(FullAdder_206_io_co)
  );
  FullAdder FullAdder_207 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_207_io_a),
    .io_b(FullAdder_207_io_b),
    .io_ci(FullAdder_207_io_ci),
    .io_s(FullAdder_207_io_s),
    .io_co(FullAdder_207_io_co)
  );
  FullAdder FullAdder_208 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_208_io_a),
    .io_b(FullAdder_208_io_b),
    .io_ci(FullAdder_208_io_ci),
    .io_s(FullAdder_208_io_s),
    .io_co(FullAdder_208_io_co)
  );
  FullAdder FullAdder_209 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_209_io_a),
    .io_b(FullAdder_209_io_b),
    .io_ci(FullAdder_209_io_ci),
    .io_s(FullAdder_209_io_s),
    .io_co(FullAdder_209_io_co)
  );
  FullAdder FullAdder_210 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_210_io_a),
    .io_b(FullAdder_210_io_b),
    .io_ci(FullAdder_210_io_ci),
    .io_s(FullAdder_210_io_s),
    .io_co(FullAdder_210_io_co)
  );
  FullAdder FullAdder_211 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_211_io_a),
    .io_b(FullAdder_211_io_b),
    .io_ci(FullAdder_211_io_ci),
    .io_s(FullAdder_211_io_s),
    .io_co(FullAdder_211_io_co)
  );
  FullAdder FullAdder_212 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_212_io_a),
    .io_b(FullAdder_212_io_b),
    .io_ci(FullAdder_212_io_ci),
    .io_s(FullAdder_212_io_s),
    .io_co(FullAdder_212_io_co)
  );
  FullAdder FullAdder_213 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_213_io_a),
    .io_b(FullAdder_213_io_b),
    .io_ci(FullAdder_213_io_ci),
    .io_s(FullAdder_213_io_s),
    .io_co(FullAdder_213_io_co)
  );
  FullAdder FullAdder_214 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_214_io_a),
    .io_b(FullAdder_214_io_b),
    .io_ci(FullAdder_214_io_ci),
    .io_s(FullAdder_214_io_s),
    .io_co(FullAdder_214_io_co)
  );
  FullAdder FullAdder_215 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_215_io_a),
    .io_b(FullAdder_215_io_b),
    .io_ci(FullAdder_215_io_ci),
    .io_s(FullAdder_215_io_s),
    .io_co(FullAdder_215_io_co)
  );
  FullAdder FullAdder_216 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_216_io_a),
    .io_b(FullAdder_216_io_b),
    .io_ci(FullAdder_216_io_ci),
    .io_s(FullAdder_216_io_s),
    .io_co(FullAdder_216_io_co)
  );
  FullAdder FullAdder_217 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_217_io_a),
    .io_b(FullAdder_217_io_b),
    .io_ci(FullAdder_217_io_ci),
    .io_s(FullAdder_217_io_s),
    .io_co(FullAdder_217_io_co)
  );
  FullAdder FullAdder_218 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_218_io_a),
    .io_b(FullAdder_218_io_b),
    .io_ci(FullAdder_218_io_ci),
    .io_s(FullAdder_218_io_s),
    .io_co(FullAdder_218_io_co)
  );
  HalfAdder HalfAdder_9 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_9_io_a),
    .io_b(HalfAdder_9_io_b),
    .io_s(HalfAdder_9_io_s),
    .io_co(HalfAdder_9_io_co)
  );
  FullAdder FullAdder_219 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_219_io_a),
    .io_b(FullAdder_219_io_b),
    .io_ci(FullAdder_219_io_ci),
    .io_s(FullAdder_219_io_s),
    .io_co(FullAdder_219_io_co)
  );
  FullAdder FullAdder_220 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_220_io_a),
    .io_b(FullAdder_220_io_b),
    .io_ci(FullAdder_220_io_ci),
    .io_s(FullAdder_220_io_s),
    .io_co(FullAdder_220_io_co)
  );
  FullAdder FullAdder_221 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_221_io_a),
    .io_b(FullAdder_221_io_b),
    .io_ci(FullAdder_221_io_ci),
    .io_s(FullAdder_221_io_s),
    .io_co(FullAdder_221_io_co)
  );
  FullAdder FullAdder_222 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_222_io_a),
    .io_b(FullAdder_222_io_b),
    .io_ci(FullAdder_222_io_ci),
    .io_s(FullAdder_222_io_s),
    .io_co(FullAdder_222_io_co)
  );
  FullAdder FullAdder_223 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_223_io_a),
    .io_b(FullAdder_223_io_b),
    .io_ci(FullAdder_223_io_ci),
    .io_s(FullAdder_223_io_s),
    .io_co(FullAdder_223_io_co)
  );
  FullAdder FullAdder_224 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_224_io_a),
    .io_b(FullAdder_224_io_b),
    .io_ci(FullAdder_224_io_ci),
    .io_s(FullAdder_224_io_s),
    .io_co(FullAdder_224_io_co)
  );
  FullAdder FullAdder_225 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_225_io_a),
    .io_b(FullAdder_225_io_b),
    .io_ci(FullAdder_225_io_ci),
    .io_s(FullAdder_225_io_s),
    .io_co(FullAdder_225_io_co)
  );
  FullAdder FullAdder_226 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_226_io_a),
    .io_b(FullAdder_226_io_b),
    .io_ci(FullAdder_226_io_ci),
    .io_s(FullAdder_226_io_s),
    .io_co(FullAdder_226_io_co)
  );
  FullAdder FullAdder_227 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_227_io_a),
    .io_b(FullAdder_227_io_b),
    .io_ci(FullAdder_227_io_ci),
    .io_s(FullAdder_227_io_s),
    .io_co(FullAdder_227_io_co)
  );
  FullAdder FullAdder_228 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_228_io_a),
    .io_b(FullAdder_228_io_b),
    .io_ci(FullAdder_228_io_ci),
    .io_s(FullAdder_228_io_s),
    .io_co(FullAdder_228_io_co)
  );
  FullAdder FullAdder_229 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_229_io_a),
    .io_b(FullAdder_229_io_b),
    .io_ci(FullAdder_229_io_ci),
    .io_s(FullAdder_229_io_s),
    .io_co(FullAdder_229_io_co)
  );
  FullAdder FullAdder_230 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_230_io_a),
    .io_b(FullAdder_230_io_b),
    .io_ci(FullAdder_230_io_ci),
    .io_s(FullAdder_230_io_s),
    .io_co(FullAdder_230_io_co)
  );
  FullAdder FullAdder_231 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_231_io_a),
    .io_b(FullAdder_231_io_b),
    .io_ci(FullAdder_231_io_ci),
    .io_s(FullAdder_231_io_s),
    .io_co(FullAdder_231_io_co)
  );
  FullAdder FullAdder_232 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_232_io_a),
    .io_b(FullAdder_232_io_b),
    .io_ci(FullAdder_232_io_ci),
    .io_s(FullAdder_232_io_s),
    .io_co(FullAdder_232_io_co)
  );
  FullAdder FullAdder_233 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_233_io_a),
    .io_b(FullAdder_233_io_b),
    .io_ci(FullAdder_233_io_ci),
    .io_s(FullAdder_233_io_s),
    .io_co(FullAdder_233_io_co)
  );
  FullAdder FullAdder_234 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_234_io_a),
    .io_b(FullAdder_234_io_b),
    .io_ci(FullAdder_234_io_ci),
    .io_s(FullAdder_234_io_s),
    .io_co(FullAdder_234_io_co)
  );
  FullAdder FullAdder_235 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_235_io_a),
    .io_b(FullAdder_235_io_b),
    .io_ci(FullAdder_235_io_ci),
    .io_s(FullAdder_235_io_s),
    .io_co(FullAdder_235_io_co)
  );
  FullAdder FullAdder_236 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_236_io_a),
    .io_b(FullAdder_236_io_b),
    .io_ci(FullAdder_236_io_ci),
    .io_s(FullAdder_236_io_s),
    .io_co(FullAdder_236_io_co)
  );
  FullAdder FullAdder_237 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_237_io_a),
    .io_b(FullAdder_237_io_b),
    .io_ci(FullAdder_237_io_ci),
    .io_s(FullAdder_237_io_s),
    .io_co(FullAdder_237_io_co)
  );
  FullAdder FullAdder_238 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_238_io_a),
    .io_b(FullAdder_238_io_b),
    .io_ci(FullAdder_238_io_ci),
    .io_s(FullAdder_238_io_s),
    .io_co(FullAdder_238_io_co)
  );
  FullAdder FullAdder_239 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_239_io_a),
    .io_b(FullAdder_239_io_b),
    .io_ci(FullAdder_239_io_ci),
    .io_s(FullAdder_239_io_s),
    .io_co(FullAdder_239_io_co)
  );
  FullAdder FullAdder_240 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_240_io_a),
    .io_b(FullAdder_240_io_b),
    .io_ci(FullAdder_240_io_ci),
    .io_s(FullAdder_240_io_s),
    .io_co(FullAdder_240_io_co)
  );
  FullAdder FullAdder_241 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_241_io_a),
    .io_b(FullAdder_241_io_b),
    .io_ci(FullAdder_241_io_ci),
    .io_s(FullAdder_241_io_s),
    .io_co(FullAdder_241_io_co)
  );
  FullAdder FullAdder_242 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_242_io_a),
    .io_b(FullAdder_242_io_b),
    .io_ci(FullAdder_242_io_ci),
    .io_s(FullAdder_242_io_s),
    .io_co(FullAdder_242_io_co)
  );
  FullAdder FullAdder_243 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_243_io_a),
    .io_b(FullAdder_243_io_b),
    .io_ci(FullAdder_243_io_ci),
    .io_s(FullAdder_243_io_s),
    .io_co(FullAdder_243_io_co)
  );
  FullAdder FullAdder_244 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_244_io_a),
    .io_b(FullAdder_244_io_b),
    .io_ci(FullAdder_244_io_ci),
    .io_s(FullAdder_244_io_s),
    .io_co(FullAdder_244_io_co)
  );
  FullAdder FullAdder_245 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_245_io_a),
    .io_b(FullAdder_245_io_b),
    .io_ci(FullAdder_245_io_ci),
    .io_s(FullAdder_245_io_s),
    .io_co(FullAdder_245_io_co)
  );
  FullAdder FullAdder_246 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_246_io_a),
    .io_b(FullAdder_246_io_b),
    .io_ci(FullAdder_246_io_ci),
    .io_s(FullAdder_246_io_s),
    .io_co(FullAdder_246_io_co)
  );
  FullAdder FullAdder_247 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_247_io_a),
    .io_b(FullAdder_247_io_b),
    .io_ci(FullAdder_247_io_ci),
    .io_s(FullAdder_247_io_s),
    .io_co(FullAdder_247_io_co)
  );
  FullAdder FullAdder_248 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_248_io_a),
    .io_b(FullAdder_248_io_b),
    .io_ci(FullAdder_248_io_ci),
    .io_s(FullAdder_248_io_s),
    .io_co(FullAdder_248_io_co)
  );
  FullAdder FullAdder_249 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_249_io_a),
    .io_b(FullAdder_249_io_b),
    .io_ci(FullAdder_249_io_ci),
    .io_s(FullAdder_249_io_s),
    .io_co(FullAdder_249_io_co)
  );
  FullAdder FullAdder_250 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_250_io_a),
    .io_b(FullAdder_250_io_b),
    .io_ci(FullAdder_250_io_ci),
    .io_s(FullAdder_250_io_s),
    .io_co(FullAdder_250_io_co)
  );
  FullAdder FullAdder_251 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_251_io_a),
    .io_b(FullAdder_251_io_b),
    .io_ci(FullAdder_251_io_ci),
    .io_s(FullAdder_251_io_s),
    .io_co(FullAdder_251_io_co)
  );
  FullAdder FullAdder_252 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_252_io_a),
    .io_b(FullAdder_252_io_b),
    .io_ci(FullAdder_252_io_ci),
    .io_s(FullAdder_252_io_s),
    .io_co(FullAdder_252_io_co)
  );
  FullAdder FullAdder_253 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_253_io_a),
    .io_b(FullAdder_253_io_b),
    .io_ci(FullAdder_253_io_ci),
    .io_s(FullAdder_253_io_s),
    .io_co(FullAdder_253_io_co)
  );
  FullAdder FullAdder_254 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_254_io_a),
    .io_b(FullAdder_254_io_b),
    .io_ci(FullAdder_254_io_ci),
    .io_s(FullAdder_254_io_s),
    .io_co(FullAdder_254_io_co)
  );
  FullAdder FullAdder_255 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_255_io_a),
    .io_b(FullAdder_255_io_b),
    .io_ci(FullAdder_255_io_ci),
    .io_s(FullAdder_255_io_s),
    .io_co(FullAdder_255_io_co)
  );
  FullAdder FullAdder_256 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_256_io_a),
    .io_b(FullAdder_256_io_b),
    .io_ci(FullAdder_256_io_ci),
    .io_s(FullAdder_256_io_s),
    .io_co(FullAdder_256_io_co)
  );
  FullAdder FullAdder_257 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_257_io_a),
    .io_b(FullAdder_257_io_b),
    .io_ci(FullAdder_257_io_ci),
    .io_s(FullAdder_257_io_s),
    .io_co(FullAdder_257_io_co)
  );
  FullAdder FullAdder_258 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_258_io_a),
    .io_b(FullAdder_258_io_b),
    .io_ci(FullAdder_258_io_ci),
    .io_s(FullAdder_258_io_s),
    .io_co(FullAdder_258_io_co)
  );
  FullAdder FullAdder_259 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_259_io_a),
    .io_b(FullAdder_259_io_b),
    .io_ci(FullAdder_259_io_ci),
    .io_s(FullAdder_259_io_s),
    .io_co(FullAdder_259_io_co)
  );
  FullAdder FullAdder_260 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_260_io_a),
    .io_b(FullAdder_260_io_b),
    .io_ci(FullAdder_260_io_ci),
    .io_s(FullAdder_260_io_s),
    .io_co(FullAdder_260_io_co)
  );
  FullAdder FullAdder_261 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_261_io_a),
    .io_b(FullAdder_261_io_b),
    .io_ci(FullAdder_261_io_ci),
    .io_s(FullAdder_261_io_s),
    .io_co(FullAdder_261_io_co)
  );
  FullAdder FullAdder_262 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_262_io_a),
    .io_b(FullAdder_262_io_b),
    .io_ci(FullAdder_262_io_ci),
    .io_s(FullAdder_262_io_s),
    .io_co(FullAdder_262_io_co)
  );
  FullAdder FullAdder_263 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_263_io_a),
    .io_b(FullAdder_263_io_b),
    .io_ci(FullAdder_263_io_ci),
    .io_s(FullAdder_263_io_s),
    .io_co(FullAdder_263_io_co)
  );
  FullAdder FullAdder_264 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_264_io_a),
    .io_b(FullAdder_264_io_b),
    .io_ci(FullAdder_264_io_ci),
    .io_s(FullAdder_264_io_s),
    .io_co(FullAdder_264_io_co)
  );
  FullAdder FullAdder_265 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_265_io_a),
    .io_b(FullAdder_265_io_b),
    .io_ci(FullAdder_265_io_ci),
    .io_s(FullAdder_265_io_s),
    .io_co(FullAdder_265_io_co)
  );
  FullAdder FullAdder_266 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_266_io_a),
    .io_b(FullAdder_266_io_b),
    .io_ci(FullAdder_266_io_ci),
    .io_s(FullAdder_266_io_s),
    .io_co(FullAdder_266_io_co)
  );
  FullAdder FullAdder_267 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_267_io_a),
    .io_b(FullAdder_267_io_b),
    .io_ci(FullAdder_267_io_ci),
    .io_s(FullAdder_267_io_s),
    .io_co(FullAdder_267_io_co)
  );
  FullAdder FullAdder_268 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_268_io_a),
    .io_b(FullAdder_268_io_b),
    .io_ci(FullAdder_268_io_ci),
    .io_s(FullAdder_268_io_s),
    .io_co(FullAdder_268_io_co)
  );
  FullAdder FullAdder_269 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_269_io_a),
    .io_b(FullAdder_269_io_b),
    .io_ci(FullAdder_269_io_ci),
    .io_s(FullAdder_269_io_s),
    .io_co(FullAdder_269_io_co)
  );
  FullAdder FullAdder_270 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_270_io_a),
    .io_b(FullAdder_270_io_b),
    .io_ci(FullAdder_270_io_ci),
    .io_s(FullAdder_270_io_s),
    .io_co(FullAdder_270_io_co)
  );
  FullAdder FullAdder_271 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_271_io_a),
    .io_b(FullAdder_271_io_b),
    .io_ci(FullAdder_271_io_ci),
    .io_s(FullAdder_271_io_s),
    .io_co(FullAdder_271_io_co)
  );
  FullAdder FullAdder_272 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_272_io_a),
    .io_b(FullAdder_272_io_b),
    .io_ci(FullAdder_272_io_ci),
    .io_s(FullAdder_272_io_s),
    .io_co(FullAdder_272_io_co)
  );
  FullAdder FullAdder_273 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_273_io_a),
    .io_b(FullAdder_273_io_b),
    .io_ci(FullAdder_273_io_ci),
    .io_s(FullAdder_273_io_s),
    .io_co(FullAdder_273_io_co)
  );
  FullAdder FullAdder_274 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_274_io_a),
    .io_b(FullAdder_274_io_b),
    .io_ci(FullAdder_274_io_ci),
    .io_s(FullAdder_274_io_s),
    .io_co(FullAdder_274_io_co)
  );
  FullAdder FullAdder_275 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_275_io_a),
    .io_b(FullAdder_275_io_b),
    .io_ci(FullAdder_275_io_ci),
    .io_s(FullAdder_275_io_s),
    .io_co(FullAdder_275_io_co)
  );
  FullAdder FullAdder_276 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_276_io_a),
    .io_b(FullAdder_276_io_b),
    .io_ci(FullAdder_276_io_ci),
    .io_s(FullAdder_276_io_s),
    .io_co(FullAdder_276_io_co)
  );
  FullAdder FullAdder_277 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_277_io_a),
    .io_b(FullAdder_277_io_b),
    .io_ci(FullAdder_277_io_ci),
    .io_s(FullAdder_277_io_s),
    .io_co(FullAdder_277_io_co)
  );
  FullAdder FullAdder_278 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_278_io_a),
    .io_b(FullAdder_278_io_b),
    .io_ci(FullAdder_278_io_ci),
    .io_s(FullAdder_278_io_s),
    .io_co(FullAdder_278_io_co)
  );
  HalfAdder HalfAdder_10 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_10_io_a),
    .io_b(HalfAdder_10_io_b),
    .io_s(HalfAdder_10_io_s),
    .io_co(HalfAdder_10_io_co)
  );
  FullAdder FullAdder_279 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_279_io_a),
    .io_b(FullAdder_279_io_b),
    .io_ci(FullAdder_279_io_ci),
    .io_s(FullAdder_279_io_s),
    .io_co(FullAdder_279_io_co)
  );
  FullAdder FullAdder_280 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_280_io_a),
    .io_b(FullAdder_280_io_b),
    .io_ci(FullAdder_280_io_ci),
    .io_s(FullAdder_280_io_s),
    .io_co(FullAdder_280_io_co)
  );
  FullAdder FullAdder_281 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_281_io_a),
    .io_b(FullAdder_281_io_b),
    .io_ci(FullAdder_281_io_ci),
    .io_s(FullAdder_281_io_s),
    .io_co(FullAdder_281_io_co)
  );
  FullAdder FullAdder_282 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_282_io_a),
    .io_b(FullAdder_282_io_b),
    .io_ci(FullAdder_282_io_ci),
    .io_s(FullAdder_282_io_s),
    .io_co(FullAdder_282_io_co)
  );
  FullAdder FullAdder_283 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_283_io_a),
    .io_b(FullAdder_283_io_b),
    .io_ci(FullAdder_283_io_ci),
    .io_s(FullAdder_283_io_s),
    .io_co(FullAdder_283_io_co)
  );
  FullAdder FullAdder_284 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_284_io_a),
    .io_b(FullAdder_284_io_b),
    .io_ci(FullAdder_284_io_ci),
    .io_s(FullAdder_284_io_s),
    .io_co(FullAdder_284_io_co)
  );
  FullAdder FullAdder_285 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_285_io_a),
    .io_b(FullAdder_285_io_b),
    .io_ci(FullAdder_285_io_ci),
    .io_s(FullAdder_285_io_s),
    .io_co(FullAdder_285_io_co)
  );
  FullAdder FullAdder_286 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_286_io_a),
    .io_b(FullAdder_286_io_b),
    .io_ci(FullAdder_286_io_ci),
    .io_s(FullAdder_286_io_s),
    .io_co(FullAdder_286_io_co)
  );
  FullAdder FullAdder_287 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_287_io_a),
    .io_b(FullAdder_287_io_b),
    .io_ci(FullAdder_287_io_ci),
    .io_s(FullAdder_287_io_s),
    .io_co(FullAdder_287_io_co)
  );
  FullAdder FullAdder_288 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_288_io_a),
    .io_b(FullAdder_288_io_b),
    .io_ci(FullAdder_288_io_ci),
    .io_s(FullAdder_288_io_s),
    .io_co(FullAdder_288_io_co)
  );
  FullAdder FullAdder_289 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_289_io_a),
    .io_b(FullAdder_289_io_b),
    .io_ci(FullAdder_289_io_ci),
    .io_s(FullAdder_289_io_s),
    .io_co(FullAdder_289_io_co)
  );
  FullAdder FullAdder_290 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_290_io_a),
    .io_b(FullAdder_290_io_b),
    .io_ci(FullAdder_290_io_ci),
    .io_s(FullAdder_290_io_s),
    .io_co(FullAdder_290_io_co)
  );
  FullAdder FullAdder_291 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_291_io_a),
    .io_b(FullAdder_291_io_b),
    .io_ci(FullAdder_291_io_ci),
    .io_s(FullAdder_291_io_s),
    .io_co(FullAdder_291_io_co)
  );
  FullAdder FullAdder_292 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_292_io_a),
    .io_b(FullAdder_292_io_b),
    .io_ci(FullAdder_292_io_ci),
    .io_s(FullAdder_292_io_s),
    .io_co(FullAdder_292_io_co)
  );
  FullAdder FullAdder_293 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_293_io_a),
    .io_b(FullAdder_293_io_b),
    .io_ci(FullAdder_293_io_ci),
    .io_s(FullAdder_293_io_s),
    .io_co(FullAdder_293_io_co)
  );
  FullAdder FullAdder_294 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_294_io_a),
    .io_b(FullAdder_294_io_b),
    .io_ci(FullAdder_294_io_ci),
    .io_s(FullAdder_294_io_s),
    .io_co(FullAdder_294_io_co)
  );
  FullAdder FullAdder_295 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_295_io_a),
    .io_b(FullAdder_295_io_b),
    .io_ci(FullAdder_295_io_ci),
    .io_s(FullAdder_295_io_s),
    .io_co(FullAdder_295_io_co)
  );
  FullAdder FullAdder_296 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_296_io_a),
    .io_b(FullAdder_296_io_b),
    .io_ci(FullAdder_296_io_ci),
    .io_s(FullAdder_296_io_s),
    .io_co(FullAdder_296_io_co)
  );
  FullAdder FullAdder_297 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_297_io_a),
    .io_b(FullAdder_297_io_b),
    .io_ci(FullAdder_297_io_ci),
    .io_s(FullAdder_297_io_s),
    .io_co(FullAdder_297_io_co)
  );
  FullAdder FullAdder_298 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_298_io_a),
    .io_b(FullAdder_298_io_b),
    .io_ci(FullAdder_298_io_ci),
    .io_s(FullAdder_298_io_s),
    .io_co(FullAdder_298_io_co)
  );
  FullAdder FullAdder_299 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_299_io_a),
    .io_b(FullAdder_299_io_b),
    .io_ci(FullAdder_299_io_ci),
    .io_s(FullAdder_299_io_s),
    .io_co(FullAdder_299_io_co)
  );
  FullAdder FullAdder_300 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_300_io_a),
    .io_b(FullAdder_300_io_b),
    .io_ci(FullAdder_300_io_ci),
    .io_s(FullAdder_300_io_s),
    .io_co(FullAdder_300_io_co)
  );
  FullAdder FullAdder_301 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_301_io_a),
    .io_b(FullAdder_301_io_b),
    .io_ci(FullAdder_301_io_ci),
    .io_s(FullAdder_301_io_s),
    .io_co(FullAdder_301_io_co)
  );
  FullAdder FullAdder_302 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_302_io_a),
    .io_b(FullAdder_302_io_b),
    .io_ci(FullAdder_302_io_ci),
    .io_s(FullAdder_302_io_s),
    .io_co(FullAdder_302_io_co)
  );
  FullAdder FullAdder_303 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_303_io_a),
    .io_b(FullAdder_303_io_b),
    .io_ci(FullAdder_303_io_ci),
    .io_s(FullAdder_303_io_s),
    .io_co(FullAdder_303_io_co)
  );
  HalfAdder HalfAdder_11 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_11_io_a),
    .io_b(HalfAdder_11_io_b),
    .io_s(HalfAdder_11_io_s),
    .io_co(HalfAdder_11_io_co)
  );
  FullAdder FullAdder_304 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_304_io_a),
    .io_b(FullAdder_304_io_b),
    .io_ci(FullAdder_304_io_ci),
    .io_s(FullAdder_304_io_s),
    .io_co(FullAdder_304_io_co)
  );
  FullAdder FullAdder_305 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_305_io_a),
    .io_b(FullAdder_305_io_b),
    .io_ci(FullAdder_305_io_ci),
    .io_s(FullAdder_305_io_s),
    .io_co(FullAdder_305_io_co)
  );
  FullAdder FullAdder_306 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_306_io_a),
    .io_b(FullAdder_306_io_b),
    .io_ci(FullAdder_306_io_ci),
    .io_s(FullAdder_306_io_s),
    .io_co(FullAdder_306_io_co)
  );
  FullAdder FullAdder_307 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_307_io_a),
    .io_b(FullAdder_307_io_b),
    .io_ci(FullAdder_307_io_ci),
    .io_s(FullAdder_307_io_s),
    .io_co(FullAdder_307_io_co)
  );
  FullAdder FullAdder_308 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_308_io_a),
    .io_b(FullAdder_308_io_b),
    .io_ci(FullAdder_308_io_ci),
    .io_s(FullAdder_308_io_s),
    .io_co(FullAdder_308_io_co)
  );
  FullAdder FullAdder_309 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_309_io_a),
    .io_b(FullAdder_309_io_b),
    .io_ci(FullAdder_309_io_ci),
    .io_s(FullAdder_309_io_s),
    .io_co(FullAdder_309_io_co)
  );
  FullAdder FullAdder_310 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_310_io_a),
    .io_b(FullAdder_310_io_b),
    .io_ci(FullAdder_310_io_ci),
    .io_s(FullAdder_310_io_s),
    .io_co(FullAdder_310_io_co)
  );
  FullAdder FullAdder_311 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_311_io_a),
    .io_b(FullAdder_311_io_b),
    .io_ci(FullAdder_311_io_ci),
    .io_s(FullAdder_311_io_s),
    .io_co(FullAdder_311_io_co)
  );
  HalfAdder HalfAdder_12 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_12_io_a),
    .io_b(HalfAdder_12_io_b),
    .io_s(HalfAdder_12_io_s),
    .io_co(HalfAdder_12_io_co)
  );
  FullAdder FullAdder_312 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_312_io_a),
    .io_b(FullAdder_312_io_b),
    .io_ci(FullAdder_312_io_ci),
    .io_s(FullAdder_312_io_s),
    .io_co(FullAdder_312_io_co)
  );
  FullAdder FullAdder_313 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_313_io_a),
    .io_b(FullAdder_313_io_b),
    .io_ci(FullAdder_313_io_ci),
    .io_s(FullAdder_313_io_s),
    .io_co(FullAdder_313_io_co)
  );
  FullAdder FullAdder_314 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_314_io_a),
    .io_b(FullAdder_314_io_b),
    .io_ci(FullAdder_314_io_ci),
    .io_s(FullAdder_314_io_s),
    .io_co(FullAdder_314_io_co)
  );
  FullAdder FullAdder_315 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_315_io_a),
    .io_b(FullAdder_315_io_b),
    .io_ci(FullAdder_315_io_ci),
    .io_s(FullAdder_315_io_s),
    .io_co(FullAdder_315_io_co)
  );
  FullAdder FullAdder_316 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_316_io_a),
    .io_b(FullAdder_316_io_b),
    .io_ci(FullAdder_316_io_ci),
    .io_s(FullAdder_316_io_s),
    .io_co(FullAdder_316_io_co)
  );
  HalfAdder HalfAdder_13 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_13_io_a),
    .io_b(HalfAdder_13_io_b),
    .io_s(HalfAdder_13_io_s),
    .io_co(HalfAdder_13_io_co)
  );
  FullAdder FullAdder_317 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_317_io_a),
    .io_b(FullAdder_317_io_b),
    .io_ci(FullAdder_317_io_ci),
    .io_s(FullAdder_317_io_s),
    .io_co(FullAdder_317_io_co)
  );
  FullAdder FullAdder_318 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_318_io_a),
    .io_b(FullAdder_318_io_b),
    .io_ci(FullAdder_318_io_ci),
    .io_s(FullAdder_318_io_s),
    .io_co(FullAdder_318_io_co)
  );
  HalfAdder HalfAdder_14 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_14_io_a),
    .io_b(HalfAdder_14_io_b),
    .io_s(HalfAdder_14_io_s),
    .io_co(HalfAdder_14_io_co)
  );
  HalfAdder HalfAdder_15 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_15_io_a),
    .io_b(HalfAdder_15_io_b),
    .io_s(HalfAdder_15_io_s),
    .io_co(HalfAdder_15_io_co)
  );
  HalfAdder HalfAdder_16 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_16_io_a),
    .io_b(HalfAdder_16_io_b),
    .io_s(HalfAdder_16_io_s),
    .io_co(HalfAdder_16_io_co)
  );
  FullAdder FullAdder_319 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_319_io_a),
    .io_b(FullAdder_319_io_b),
    .io_ci(FullAdder_319_io_ci),
    .io_s(FullAdder_319_io_s),
    .io_co(FullAdder_319_io_co)
  );
  FullAdder FullAdder_320 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_320_io_a),
    .io_b(FullAdder_320_io_b),
    .io_ci(FullAdder_320_io_ci),
    .io_s(FullAdder_320_io_s),
    .io_co(FullAdder_320_io_co)
  );
  FullAdder FullAdder_321 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_321_io_a),
    .io_b(FullAdder_321_io_b),
    .io_ci(FullAdder_321_io_ci),
    .io_s(FullAdder_321_io_s),
    .io_co(FullAdder_321_io_co)
  );
  FullAdder FullAdder_322 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_322_io_a),
    .io_b(FullAdder_322_io_b),
    .io_ci(FullAdder_322_io_ci),
    .io_s(FullAdder_322_io_s),
    .io_co(FullAdder_322_io_co)
  );
  HalfAdder HalfAdder_17 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_17_io_a),
    .io_b(HalfAdder_17_io_b),
    .io_s(HalfAdder_17_io_s),
    .io_co(HalfAdder_17_io_co)
  );
  FullAdder FullAdder_323 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_323_io_a),
    .io_b(FullAdder_323_io_b),
    .io_ci(FullAdder_323_io_ci),
    .io_s(FullAdder_323_io_s),
    .io_co(FullAdder_323_io_co)
  );
  FullAdder FullAdder_324 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_324_io_a),
    .io_b(FullAdder_324_io_b),
    .io_ci(FullAdder_324_io_ci),
    .io_s(FullAdder_324_io_s),
    .io_co(FullAdder_324_io_co)
  );
  FullAdder FullAdder_325 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_325_io_a),
    .io_b(FullAdder_325_io_b),
    .io_ci(FullAdder_325_io_ci),
    .io_s(FullAdder_325_io_s),
    .io_co(FullAdder_325_io_co)
  );
  FullAdder FullAdder_326 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_326_io_a),
    .io_b(FullAdder_326_io_b),
    .io_ci(FullAdder_326_io_ci),
    .io_s(FullAdder_326_io_s),
    .io_co(FullAdder_326_io_co)
  );
  FullAdder FullAdder_327 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_327_io_a),
    .io_b(FullAdder_327_io_b),
    .io_ci(FullAdder_327_io_ci),
    .io_s(FullAdder_327_io_s),
    .io_co(FullAdder_327_io_co)
  );
  FullAdder FullAdder_328 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_328_io_a),
    .io_b(FullAdder_328_io_b),
    .io_ci(FullAdder_328_io_ci),
    .io_s(FullAdder_328_io_s),
    .io_co(FullAdder_328_io_co)
  );
  HalfAdder HalfAdder_18 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_18_io_a),
    .io_b(HalfAdder_18_io_b),
    .io_s(HalfAdder_18_io_s),
    .io_co(HalfAdder_18_io_co)
  );
  FullAdder FullAdder_329 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_329_io_a),
    .io_b(FullAdder_329_io_b),
    .io_ci(FullAdder_329_io_ci),
    .io_s(FullAdder_329_io_s),
    .io_co(FullAdder_329_io_co)
  );
  FullAdder FullAdder_330 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_330_io_a),
    .io_b(FullAdder_330_io_b),
    .io_ci(FullAdder_330_io_ci),
    .io_s(FullAdder_330_io_s),
    .io_co(FullAdder_330_io_co)
  );
  HalfAdder HalfAdder_19 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_19_io_a),
    .io_b(HalfAdder_19_io_b),
    .io_s(HalfAdder_19_io_s),
    .io_co(HalfAdder_19_io_co)
  );
  FullAdder FullAdder_331 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_331_io_a),
    .io_b(FullAdder_331_io_b),
    .io_ci(FullAdder_331_io_ci),
    .io_s(FullAdder_331_io_s),
    .io_co(FullAdder_331_io_co)
  );
  FullAdder FullAdder_332 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_332_io_a),
    .io_b(FullAdder_332_io_b),
    .io_ci(FullAdder_332_io_ci),
    .io_s(FullAdder_332_io_s),
    .io_co(FullAdder_332_io_co)
  );
  HalfAdder HalfAdder_20 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_20_io_a),
    .io_b(HalfAdder_20_io_b),
    .io_s(HalfAdder_20_io_s),
    .io_co(HalfAdder_20_io_co)
  );
  FullAdder FullAdder_333 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_333_io_a),
    .io_b(FullAdder_333_io_b),
    .io_ci(FullAdder_333_io_ci),
    .io_s(FullAdder_333_io_s),
    .io_co(FullAdder_333_io_co)
  );
  FullAdder FullAdder_334 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_334_io_a),
    .io_b(FullAdder_334_io_b),
    .io_ci(FullAdder_334_io_ci),
    .io_s(FullAdder_334_io_s),
    .io_co(FullAdder_334_io_co)
  );
  FullAdder FullAdder_335 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_335_io_a),
    .io_b(FullAdder_335_io_b),
    .io_ci(FullAdder_335_io_ci),
    .io_s(FullAdder_335_io_s),
    .io_co(FullAdder_335_io_co)
  );
  FullAdder FullAdder_336 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_336_io_a),
    .io_b(FullAdder_336_io_b),
    .io_ci(FullAdder_336_io_ci),
    .io_s(FullAdder_336_io_s),
    .io_co(FullAdder_336_io_co)
  );
  FullAdder FullAdder_337 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_337_io_a),
    .io_b(FullAdder_337_io_b),
    .io_ci(FullAdder_337_io_ci),
    .io_s(FullAdder_337_io_s),
    .io_co(FullAdder_337_io_co)
  );
  FullAdder FullAdder_338 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_338_io_a),
    .io_b(FullAdder_338_io_b),
    .io_ci(FullAdder_338_io_ci),
    .io_s(FullAdder_338_io_s),
    .io_co(FullAdder_338_io_co)
  );
  FullAdder FullAdder_339 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_339_io_a),
    .io_b(FullAdder_339_io_b),
    .io_ci(FullAdder_339_io_ci),
    .io_s(FullAdder_339_io_s),
    .io_co(FullAdder_339_io_co)
  );
  FullAdder FullAdder_340 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_340_io_a),
    .io_b(FullAdder_340_io_b),
    .io_ci(FullAdder_340_io_ci),
    .io_s(FullAdder_340_io_s),
    .io_co(FullAdder_340_io_co)
  );
  FullAdder FullAdder_341 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_341_io_a),
    .io_b(FullAdder_341_io_b),
    .io_ci(FullAdder_341_io_ci),
    .io_s(FullAdder_341_io_s),
    .io_co(FullAdder_341_io_co)
  );
  FullAdder FullAdder_342 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_342_io_a),
    .io_b(FullAdder_342_io_b),
    .io_ci(FullAdder_342_io_ci),
    .io_s(FullAdder_342_io_s),
    .io_co(FullAdder_342_io_co)
  );
  FullAdder FullAdder_343 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_343_io_a),
    .io_b(FullAdder_343_io_b),
    .io_ci(FullAdder_343_io_ci),
    .io_s(FullAdder_343_io_s),
    .io_co(FullAdder_343_io_co)
  );
  FullAdder FullAdder_344 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_344_io_a),
    .io_b(FullAdder_344_io_b),
    .io_ci(FullAdder_344_io_ci),
    .io_s(FullAdder_344_io_s),
    .io_co(FullAdder_344_io_co)
  );
  FullAdder FullAdder_345 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_345_io_a),
    .io_b(FullAdder_345_io_b),
    .io_ci(FullAdder_345_io_ci),
    .io_s(FullAdder_345_io_s),
    .io_co(FullAdder_345_io_co)
  );
  FullAdder FullAdder_346 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_346_io_a),
    .io_b(FullAdder_346_io_b),
    .io_ci(FullAdder_346_io_ci),
    .io_s(FullAdder_346_io_s),
    .io_co(FullAdder_346_io_co)
  );
  FullAdder FullAdder_347 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_347_io_a),
    .io_b(FullAdder_347_io_b),
    .io_ci(FullAdder_347_io_ci),
    .io_s(FullAdder_347_io_s),
    .io_co(FullAdder_347_io_co)
  );
  FullAdder FullAdder_348 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_348_io_a),
    .io_b(FullAdder_348_io_b),
    .io_ci(FullAdder_348_io_ci),
    .io_s(FullAdder_348_io_s),
    .io_co(FullAdder_348_io_co)
  );
  FullAdder FullAdder_349 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_349_io_a),
    .io_b(FullAdder_349_io_b),
    .io_ci(FullAdder_349_io_ci),
    .io_s(FullAdder_349_io_s),
    .io_co(FullAdder_349_io_co)
  );
  FullAdder FullAdder_350 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_350_io_a),
    .io_b(FullAdder_350_io_b),
    .io_ci(FullAdder_350_io_ci),
    .io_s(FullAdder_350_io_s),
    .io_co(FullAdder_350_io_co)
  );
  FullAdder FullAdder_351 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_351_io_a),
    .io_b(FullAdder_351_io_b),
    .io_ci(FullAdder_351_io_ci),
    .io_s(FullAdder_351_io_s),
    .io_co(FullAdder_351_io_co)
  );
  FullAdder FullAdder_352 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_352_io_a),
    .io_b(FullAdder_352_io_b),
    .io_ci(FullAdder_352_io_ci),
    .io_s(FullAdder_352_io_s),
    .io_co(FullAdder_352_io_co)
  );
  FullAdder FullAdder_353 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_353_io_a),
    .io_b(FullAdder_353_io_b),
    .io_ci(FullAdder_353_io_ci),
    .io_s(FullAdder_353_io_s),
    .io_co(FullAdder_353_io_co)
  );
  FullAdder FullAdder_354 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_354_io_a),
    .io_b(FullAdder_354_io_b),
    .io_ci(FullAdder_354_io_ci),
    .io_s(FullAdder_354_io_s),
    .io_co(FullAdder_354_io_co)
  );
  FullAdder FullAdder_355 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_355_io_a),
    .io_b(FullAdder_355_io_b),
    .io_ci(FullAdder_355_io_ci),
    .io_s(FullAdder_355_io_s),
    .io_co(FullAdder_355_io_co)
  );
  FullAdder FullAdder_356 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_356_io_a),
    .io_b(FullAdder_356_io_b),
    .io_ci(FullAdder_356_io_ci),
    .io_s(FullAdder_356_io_s),
    .io_co(FullAdder_356_io_co)
  );
  FullAdder FullAdder_357 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_357_io_a),
    .io_b(FullAdder_357_io_b),
    .io_ci(FullAdder_357_io_ci),
    .io_s(FullAdder_357_io_s),
    .io_co(FullAdder_357_io_co)
  );
  FullAdder FullAdder_358 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_358_io_a),
    .io_b(FullAdder_358_io_b),
    .io_ci(FullAdder_358_io_ci),
    .io_s(FullAdder_358_io_s),
    .io_co(FullAdder_358_io_co)
  );
  FullAdder FullAdder_359 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_359_io_a),
    .io_b(FullAdder_359_io_b),
    .io_ci(FullAdder_359_io_ci),
    .io_s(FullAdder_359_io_s),
    .io_co(FullAdder_359_io_co)
  );
  FullAdder FullAdder_360 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_360_io_a),
    .io_b(FullAdder_360_io_b),
    .io_ci(FullAdder_360_io_ci),
    .io_s(FullAdder_360_io_s),
    .io_co(FullAdder_360_io_co)
  );
  FullAdder FullAdder_361 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_361_io_a),
    .io_b(FullAdder_361_io_b),
    .io_ci(FullAdder_361_io_ci),
    .io_s(FullAdder_361_io_s),
    .io_co(FullAdder_361_io_co)
  );
  FullAdder FullAdder_362 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_362_io_a),
    .io_b(FullAdder_362_io_b),
    .io_ci(FullAdder_362_io_ci),
    .io_s(FullAdder_362_io_s),
    .io_co(FullAdder_362_io_co)
  );
  FullAdder FullAdder_363 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_363_io_a),
    .io_b(FullAdder_363_io_b),
    .io_ci(FullAdder_363_io_ci),
    .io_s(FullAdder_363_io_s),
    .io_co(FullAdder_363_io_co)
  );
  FullAdder FullAdder_364 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_364_io_a),
    .io_b(FullAdder_364_io_b),
    .io_ci(FullAdder_364_io_ci),
    .io_s(FullAdder_364_io_s),
    .io_co(FullAdder_364_io_co)
  );
  FullAdder FullAdder_365 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_365_io_a),
    .io_b(FullAdder_365_io_b),
    .io_ci(FullAdder_365_io_ci),
    .io_s(FullAdder_365_io_s),
    .io_co(FullAdder_365_io_co)
  );
  FullAdder FullAdder_366 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_366_io_a),
    .io_b(FullAdder_366_io_b),
    .io_ci(FullAdder_366_io_ci),
    .io_s(FullAdder_366_io_s),
    .io_co(FullAdder_366_io_co)
  );
  HalfAdder HalfAdder_21 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_21_io_a),
    .io_b(HalfAdder_21_io_b),
    .io_s(HalfAdder_21_io_s),
    .io_co(HalfAdder_21_io_co)
  );
  FullAdder FullAdder_367 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_367_io_a),
    .io_b(FullAdder_367_io_b),
    .io_ci(FullAdder_367_io_ci),
    .io_s(FullAdder_367_io_s),
    .io_co(FullAdder_367_io_co)
  );
  FullAdder FullAdder_368 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_368_io_a),
    .io_b(FullAdder_368_io_b),
    .io_ci(FullAdder_368_io_ci),
    .io_s(FullAdder_368_io_s),
    .io_co(FullAdder_368_io_co)
  );
  FullAdder FullAdder_369 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_369_io_a),
    .io_b(FullAdder_369_io_b),
    .io_ci(FullAdder_369_io_ci),
    .io_s(FullAdder_369_io_s),
    .io_co(FullAdder_369_io_co)
  );
  FullAdder FullAdder_370 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_370_io_a),
    .io_b(FullAdder_370_io_b),
    .io_ci(FullAdder_370_io_ci),
    .io_s(FullAdder_370_io_s),
    .io_co(FullAdder_370_io_co)
  );
  FullAdder FullAdder_371 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_371_io_a),
    .io_b(FullAdder_371_io_b),
    .io_ci(FullAdder_371_io_ci),
    .io_s(FullAdder_371_io_s),
    .io_co(FullAdder_371_io_co)
  );
  FullAdder FullAdder_372 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_372_io_a),
    .io_b(FullAdder_372_io_b),
    .io_ci(FullAdder_372_io_ci),
    .io_s(FullAdder_372_io_s),
    .io_co(FullAdder_372_io_co)
  );
  FullAdder FullAdder_373 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_373_io_a),
    .io_b(FullAdder_373_io_b),
    .io_ci(FullAdder_373_io_ci),
    .io_s(FullAdder_373_io_s),
    .io_co(FullAdder_373_io_co)
  );
  FullAdder FullAdder_374 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_374_io_a),
    .io_b(FullAdder_374_io_b),
    .io_ci(FullAdder_374_io_ci),
    .io_s(FullAdder_374_io_s),
    .io_co(FullAdder_374_io_co)
  );
  FullAdder FullAdder_375 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_375_io_a),
    .io_b(FullAdder_375_io_b),
    .io_ci(FullAdder_375_io_ci),
    .io_s(FullAdder_375_io_s),
    .io_co(FullAdder_375_io_co)
  );
  FullAdder FullAdder_376 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_376_io_a),
    .io_b(FullAdder_376_io_b),
    .io_ci(FullAdder_376_io_ci),
    .io_s(FullAdder_376_io_s),
    .io_co(FullAdder_376_io_co)
  );
  FullAdder FullAdder_377 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_377_io_a),
    .io_b(FullAdder_377_io_b),
    .io_ci(FullAdder_377_io_ci),
    .io_s(FullAdder_377_io_s),
    .io_co(FullAdder_377_io_co)
  );
  FullAdder FullAdder_378 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_378_io_a),
    .io_b(FullAdder_378_io_b),
    .io_ci(FullAdder_378_io_ci),
    .io_s(FullAdder_378_io_s),
    .io_co(FullAdder_378_io_co)
  );
  FullAdder FullAdder_379 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_379_io_a),
    .io_b(FullAdder_379_io_b),
    .io_ci(FullAdder_379_io_ci),
    .io_s(FullAdder_379_io_s),
    .io_co(FullAdder_379_io_co)
  );
  FullAdder FullAdder_380 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_380_io_a),
    .io_b(FullAdder_380_io_b),
    .io_ci(FullAdder_380_io_ci),
    .io_s(FullAdder_380_io_s),
    .io_co(FullAdder_380_io_co)
  );
  FullAdder FullAdder_381 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_381_io_a),
    .io_b(FullAdder_381_io_b),
    .io_ci(FullAdder_381_io_ci),
    .io_s(FullAdder_381_io_s),
    .io_co(FullAdder_381_io_co)
  );
  FullAdder FullAdder_382 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_382_io_a),
    .io_b(FullAdder_382_io_b),
    .io_ci(FullAdder_382_io_ci),
    .io_s(FullAdder_382_io_s),
    .io_co(FullAdder_382_io_co)
  );
  FullAdder FullAdder_383 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_383_io_a),
    .io_b(FullAdder_383_io_b),
    .io_ci(FullAdder_383_io_ci),
    .io_s(FullAdder_383_io_s),
    .io_co(FullAdder_383_io_co)
  );
  FullAdder FullAdder_384 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_384_io_a),
    .io_b(FullAdder_384_io_b),
    .io_ci(FullAdder_384_io_ci),
    .io_s(FullAdder_384_io_s),
    .io_co(FullAdder_384_io_co)
  );
  FullAdder FullAdder_385 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_385_io_a),
    .io_b(FullAdder_385_io_b),
    .io_ci(FullAdder_385_io_ci),
    .io_s(FullAdder_385_io_s),
    .io_co(FullAdder_385_io_co)
  );
  FullAdder FullAdder_386 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_386_io_a),
    .io_b(FullAdder_386_io_b),
    .io_ci(FullAdder_386_io_ci),
    .io_s(FullAdder_386_io_s),
    .io_co(FullAdder_386_io_co)
  );
  HalfAdder HalfAdder_22 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_22_io_a),
    .io_b(HalfAdder_22_io_b),
    .io_s(HalfAdder_22_io_s),
    .io_co(HalfAdder_22_io_co)
  );
  FullAdder FullAdder_387 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_387_io_a),
    .io_b(FullAdder_387_io_b),
    .io_ci(FullAdder_387_io_ci),
    .io_s(FullAdder_387_io_s),
    .io_co(FullAdder_387_io_co)
  );
  FullAdder FullAdder_388 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_388_io_a),
    .io_b(FullAdder_388_io_b),
    .io_ci(FullAdder_388_io_ci),
    .io_s(FullAdder_388_io_s),
    .io_co(FullAdder_388_io_co)
  );
  FullAdder FullAdder_389 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_389_io_a),
    .io_b(FullAdder_389_io_b),
    .io_ci(FullAdder_389_io_ci),
    .io_s(FullAdder_389_io_s),
    .io_co(FullAdder_389_io_co)
  );
  FullAdder FullAdder_390 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_390_io_a),
    .io_b(FullAdder_390_io_b),
    .io_ci(FullAdder_390_io_ci),
    .io_s(FullAdder_390_io_s),
    .io_co(FullAdder_390_io_co)
  );
  FullAdder FullAdder_391 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_391_io_a),
    .io_b(FullAdder_391_io_b),
    .io_ci(FullAdder_391_io_ci),
    .io_s(FullAdder_391_io_s),
    .io_co(FullAdder_391_io_co)
  );
  FullAdder FullAdder_392 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_392_io_a),
    .io_b(FullAdder_392_io_b),
    .io_ci(FullAdder_392_io_ci),
    .io_s(FullAdder_392_io_s),
    .io_co(FullAdder_392_io_co)
  );
  FullAdder FullAdder_393 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_393_io_a),
    .io_b(FullAdder_393_io_b),
    .io_ci(FullAdder_393_io_ci),
    .io_s(FullAdder_393_io_s),
    .io_co(FullAdder_393_io_co)
  );
  FullAdder FullAdder_394 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_394_io_a),
    .io_b(FullAdder_394_io_b),
    .io_ci(FullAdder_394_io_ci),
    .io_s(FullAdder_394_io_s),
    .io_co(FullAdder_394_io_co)
  );
  FullAdder FullAdder_395 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_395_io_a),
    .io_b(FullAdder_395_io_b),
    .io_ci(FullAdder_395_io_ci),
    .io_s(FullAdder_395_io_s),
    .io_co(FullAdder_395_io_co)
  );
  FullAdder FullAdder_396 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_396_io_a),
    .io_b(FullAdder_396_io_b),
    .io_ci(FullAdder_396_io_ci),
    .io_s(FullAdder_396_io_s),
    .io_co(FullAdder_396_io_co)
  );
  FullAdder FullAdder_397 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_397_io_a),
    .io_b(FullAdder_397_io_b),
    .io_ci(FullAdder_397_io_ci),
    .io_s(FullAdder_397_io_s),
    .io_co(FullAdder_397_io_co)
  );
  FullAdder FullAdder_398 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_398_io_a),
    .io_b(FullAdder_398_io_b),
    .io_ci(FullAdder_398_io_ci),
    .io_s(FullAdder_398_io_s),
    .io_co(FullAdder_398_io_co)
  );
  FullAdder FullAdder_399 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_399_io_a),
    .io_b(FullAdder_399_io_b),
    .io_ci(FullAdder_399_io_ci),
    .io_s(FullAdder_399_io_s),
    .io_co(FullAdder_399_io_co)
  );
  FullAdder FullAdder_400 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_400_io_a),
    .io_b(FullAdder_400_io_b),
    .io_ci(FullAdder_400_io_ci),
    .io_s(FullAdder_400_io_s),
    .io_co(FullAdder_400_io_co)
  );
  FullAdder FullAdder_401 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_401_io_a),
    .io_b(FullAdder_401_io_b),
    .io_ci(FullAdder_401_io_ci),
    .io_s(FullAdder_401_io_s),
    .io_co(FullAdder_401_io_co)
  );
  FullAdder FullAdder_402 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_402_io_a),
    .io_b(FullAdder_402_io_b),
    .io_ci(FullAdder_402_io_ci),
    .io_s(FullAdder_402_io_s),
    .io_co(FullAdder_402_io_co)
  );
  FullAdder FullAdder_403 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_403_io_a),
    .io_b(FullAdder_403_io_b),
    .io_ci(FullAdder_403_io_ci),
    .io_s(FullAdder_403_io_s),
    .io_co(FullAdder_403_io_co)
  );
  FullAdder FullAdder_404 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_404_io_a),
    .io_b(FullAdder_404_io_b),
    .io_ci(FullAdder_404_io_ci),
    .io_s(FullAdder_404_io_s),
    .io_co(FullAdder_404_io_co)
  );
  HalfAdder HalfAdder_23 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_23_io_a),
    .io_b(HalfAdder_23_io_b),
    .io_s(HalfAdder_23_io_s),
    .io_co(HalfAdder_23_io_co)
  );
  FullAdder FullAdder_405 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_405_io_a),
    .io_b(FullAdder_405_io_b),
    .io_ci(FullAdder_405_io_ci),
    .io_s(FullAdder_405_io_s),
    .io_co(FullAdder_405_io_co)
  );
  FullAdder FullAdder_406 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_406_io_a),
    .io_b(FullAdder_406_io_b),
    .io_ci(FullAdder_406_io_ci),
    .io_s(FullAdder_406_io_s),
    .io_co(FullAdder_406_io_co)
  );
  FullAdder FullAdder_407 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_407_io_a),
    .io_b(FullAdder_407_io_b),
    .io_ci(FullAdder_407_io_ci),
    .io_s(FullAdder_407_io_s),
    .io_co(FullAdder_407_io_co)
  );
  FullAdder FullAdder_408 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_408_io_a),
    .io_b(FullAdder_408_io_b),
    .io_ci(FullAdder_408_io_ci),
    .io_s(FullAdder_408_io_s),
    .io_co(FullAdder_408_io_co)
  );
  FullAdder FullAdder_409 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_409_io_a),
    .io_b(FullAdder_409_io_b),
    .io_ci(FullAdder_409_io_ci),
    .io_s(FullAdder_409_io_s),
    .io_co(FullAdder_409_io_co)
  );
  FullAdder FullAdder_410 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_410_io_a),
    .io_b(FullAdder_410_io_b),
    .io_ci(FullAdder_410_io_ci),
    .io_s(FullAdder_410_io_s),
    .io_co(FullAdder_410_io_co)
  );
  HalfAdder HalfAdder_24 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_24_io_a),
    .io_b(HalfAdder_24_io_b),
    .io_s(HalfAdder_24_io_s),
    .io_co(HalfAdder_24_io_co)
  );
  FullAdder FullAdder_411 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_411_io_a),
    .io_b(FullAdder_411_io_b),
    .io_ci(FullAdder_411_io_ci),
    .io_s(FullAdder_411_io_s),
    .io_co(FullAdder_411_io_co)
  );
  FullAdder FullAdder_412 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_412_io_a),
    .io_b(FullAdder_412_io_b),
    .io_ci(FullAdder_412_io_ci),
    .io_s(FullAdder_412_io_s),
    .io_co(FullAdder_412_io_co)
  );
  FullAdder FullAdder_413 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_413_io_a),
    .io_b(FullAdder_413_io_b),
    .io_ci(FullAdder_413_io_ci),
    .io_s(FullAdder_413_io_s),
    .io_co(FullAdder_413_io_co)
  );
  FullAdder FullAdder_414 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_414_io_a),
    .io_b(FullAdder_414_io_b),
    .io_ci(FullAdder_414_io_ci),
    .io_s(FullAdder_414_io_s),
    .io_co(FullAdder_414_io_co)
  );
  FullAdder FullAdder_415 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_415_io_a),
    .io_b(FullAdder_415_io_b),
    .io_ci(FullAdder_415_io_ci),
    .io_s(FullAdder_415_io_s),
    .io_co(FullAdder_415_io_co)
  );
  FullAdder FullAdder_416 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_416_io_a),
    .io_b(FullAdder_416_io_b),
    .io_ci(FullAdder_416_io_ci),
    .io_s(FullAdder_416_io_s),
    .io_co(FullAdder_416_io_co)
  );
  FullAdder FullAdder_417 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_417_io_a),
    .io_b(FullAdder_417_io_b),
    .io_ci(FullAdder_417_io_ci),
    .io_s(FullAdder_417_io_s),
    .io_co(FullAdder_417_io_co)
  );
  FullAdder FullAdder_418 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_418_io_a),
    .io_b(FullAdder_418_io_b),
    .io_ci(FullAdder_418_io_ci),
    .io_s(FullAdder_418_io_s),
    .io_co(FullAdder_418_io_co)
  );
  FullAdder FullAdder_419 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_419_io_a),
    .io_b(FullAdder_419_io_b),
    .io_ci(FullAdder_419_io_ci),
    .io_s(FullAdder_419_io_s),
    .io_co(FullAdder_419_io_co)
  );
  FullAdder FullAdder_420 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_420_io_a),
    .io_b(FullAdder_420_io_b),
    .io_ci(FullAdder_420_io_ci),
    .io_s(FullAdder_420_io_s),
    .io_co(FullAdder_420_io_co)
  );
  FullAdder FullAdder_421 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_421_io_a),
    .io_b(FullAdder_421_io_b),
    .io_ci(FullAdder_421_io_ci),
    .io_s(FullAdder_421_io_s),
    .io_co(FullAdder_421_io_co)
  );
  FullAdder FullAdder_422 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_422_io_a),
    .io_b(FullAdder_422_io_b),
    .io_ci(FullAdder_422_io_ci),
    .io_s(FullAdder_422_io_s),
    .io_co(FullAdder_422_io_co)
  );
  FullAdder FullAdder_423 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_423_io_a),
    .io_b(FullAdder_423_io_b),
    .io_ci(FullAdder_423_io_ci),
    .io_s(FullAdder_423_io_s),
    .io_co(FullAdder_423_io_co)
  );
  FullAdder FullAdder_424 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_424_io_a),
    .io_b(FullAdder_424_io_b),
    .io_ci(FullAdder_424_io_ci),
    .io_s(FullAdder_424_io_s),
    .io_co(FullAdder_424_io_co)
  );
  FullAdder FullAdder_425 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_425_io_a),
    .io_b(FullAdder_425_io_b),
    .io_ci(FullAdder_425_io_ci),
    .io_s(FullAdder_425_io_s),
    .io_co(FullAdder_425_io_co)
  );
  FullAdder FullAdder_426 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_426_io_a),
    .io_b(FullAdder_426_io_b),
    .io_ci(FullAdder_426_io_ci),
    .io_s(FullAdder_426_io_s),
    .io_co(FullAdder_426_io_co)
  );
  FullAdder FullAdder_427 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_427_io_a),
    .io_b(FullAdder_427_io_b),
    .io_ci(FullAdder_427_io_ci),
    .io_s(FullAdder_427_io_s),
    .io_co(FullAdder_427_io_co)
  );
  FullAdder FullAdder_428 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_428_io_a),
    .io_b(FullAdder_428_io_b),
    .io_ci(FullAdder_428_io_ci),
    .io_s(FullAdder_428_io_s),
    .io_co(FullAdder_428_io_co)
  );
  FullAdder FullAdder_429 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_429_io_a),
    .io_b(FullAdder_429_io_b),
    .io_ci(FullAdder_429_io_ci),
    .io_s(FullAdder_429_io_s),
    .io_co(FullAdder_429_io_co)
  );
  FullAdder FullAdder_430 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_430_io_a),
    .io_b(FullAdder_430_io_b),
    .io_ci(FullAdder_430_io_ci),
    .io_s(FullAdder_430_io_s),
    .io_co(FullAdder_430_io_co)
  );
  FullAdder FullAdder_431 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_431_io_a),
    .io_b(FullAdder_431_io_b),
    .io_ci(FullAdder_431_io_ci),
    .io_s(FullAdder_431_io_s),
    .io_co(FullAdder_431_io_co)
  );
  FullAdder FullAdder_432 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_432_io_a),
    .io_b(FullAdder_432_io_b),
    .io_ci(FullAdder_432_io_ci),
    .io_s(FullAdder_432_io_s),
    .io_co(FullAdder_432_io_co)
  );
  FullAdder FullAdder_433 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_433_io_a),
    .io_b(FullAdder_433_io_b),
    .io_ci(FullAdder_433_io_ci),
    .io_s(FullAdder_433_io_s),
    .io_co(FullAdder_433_io_co)
  );
  FullAdder FullAdder_434 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_434_io_a),
    .io_b(FullAdder_434_io_b),
    .io_ci(FullAdder_434_io_ci),
    .io_s(FullAdder_434_io_s),
    .io_co(FullAdder_434_io_co)
  );
  FullAdder FullAdder_435 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_435_io_a),
    .io_b(FullAdder_435_io_b),
    .io_ci(FullAdder_435_io_ci),
    .io_s(FullAdder_435_io_s),
    .io_co(FullAdder_435_io_co)
  );
  FullAdder FullAdder_436 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_436_io_a),
    .io_b(FullAdder_436_io_b),
    .io_ci(FullAdder_436_io_ci),
    .io_s(FullAdder_436_io_s),
    .io_co(FullAdder_436_io_co)
  );
  FullAdder FullAdder_437 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_437_io_a),
    .io_b(FullAdder_437_io_b),
    .io_ci(FullAdder_437_io_ci),
    .io_s(FullAdder_437_io_s),
    .io_co(FullAdder_437_io_co)
  );
  FullAdder FullAdder_438 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_438_io_a),
    .io_b(FullAdder_438_io_b),
    .io_ci(FullAdder_438_io_ci),
    .io_s(FullAdder_438_io_s),
    .io_co(FullAdder_438_io_co)
  );
  FullAdder FullAdder_439 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_439_io_a),
    .io_b(FullAdder_439_io_b),
    .io_ci(FullAdder_439_io_ci),
    .io_s(FullAdder_439_io_s),
    .io_co(FullAdder_439_io_co)
  );
  FullAdder FullAdder_440 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_440_io_a),
    .io_b(FullAdder_440_io_b),
    .io_ci(FullAdder_440_io_ci),
    .io_s(FullAdder_440_io_s),
    .io_co(FullAdder_440_io_co)
  );
  FullAdder FullAdder_441 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_441_io_a),
    .io_b(FullAdder_441_io_b),
    .io_ci(FullAdder_441_io_ci),
    .io_s(FullAdder_441_io_s),
    .io_co(FullAdder_441_io_co)
  );
  FullAdder FullAdder_442 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_442_io_a),
    .io_b(FullAdder_442_io_b),
    .io_ci(FullAdder_442_io_ci),
    .io_s(FullAdder_442_io_s),
    .io_co(FullAdder_442_io_co)
  );
  FullAdder FullAdder_443 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_443_io_a),
    .io_b(FullAdder_443_io_b),
    .io_ci(FullAdder_443_io_ci),
    .io_s(FullAdder_443_io_s),
    .io_co(FullAdder_443_io_co)
  );
  FullAdder FullAdder_444 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_444_io_a),
    .io_b(FullAdder_444_io_b),
    .io_ci(FullAdder_444_io_ci),
    .io_s(FullAdder_444_io_s),
    .io_co(FullAdder_444_io_co)
  );
  FullAdder FullAdder_445 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_445_io_a),
    .io_b(FullAdder_445_io_b),
    .io_ci(FullAdder_445_io_ci),
    .io_s(FullAdder_445_io_s),
    .io_co(FullAdder_445_io_co)
  );
  FullAdder FullAdder_446 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_446_io_a),
    .io_b(FullAdder_446_io_b),
    .io_ci(FullAdder_446_io_ci),
    .io_s(FullAdder_446_io_s),
    .io_co(FullAdder_446_io_co)
  );
  FullAdder FullAdder_447 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_447_io_a),
    .io_b(FullAdder_447_io_b),
    .io_ci(FullAdder_447_io_ci),
    .io_s(FullAdder_447_io_s),
    .io_co(FullAdder_447_io_co)
  );
  FullAdder FullAdder_448 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_448_io_a),
    .io_b(FullAdder_448_io_b),
    .io_ci(FullAdder_448_io_ci),
    .io_s(FullAdder_448_io_s),
    .io_co(FullAdder_448_io_co)
  );
  FullAdder FullAdder_449 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_449_io_a),
    .io_b(FullAdder_449_io_b),
    .io_ci(FullAdder_449_io_ci),
    .io_s(FullAdder_449_io_s),
    .io_co(FullAdder_449_io_co)
  );
  FullAdder FullAdder_450 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_450_io_a),
    .io_b(FullAdder_450_io_b),
    .io_ci(FullAdder_450_io_ci),
    .io_s(FullAdder_450_io_s),
    .io_co(FullAdder_450_io_co)
  );
  FullAdder FullAdder_451 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_451_io_a),
    .io_b(FullAdder_451_io_b),
    .io_ci(FullAdder_451_io_ci),
    .io_s(FullAdder_451_io_s),
    .io_co(FullAdder_451_io_co)
  );
  FullAdder FullAdder_452 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_452_io_a),
    .io_b(FullAdder_452_io_b),
    .io_ci(FullAdder_452_io_ci),
    .io_s(FullAdder_452_io_s),
    .io_co(FullAdder_452_io_co)
  );
  FullAdder FullAdder_453 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_453_io_a),
    .io_b(FullAdder_453_io_b),
    .io_ci(FullAdder_453_io_ci),
    .io_s(FullAdder_453_io_s),
    .io_co(FullAdder_453_io_co)
  );
  FullAdder FullAdder_454 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_454_io_a),
    .io_b(FullAdder_454_io_b),
    .io_ci(FullAdder_454_io_ci),
    .io_s(FullAdder_454_io_s),
    .io_co(FullAdder_454_io_co)
  );
  FullAdder FullAdder_455 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_455_io_a),
    .io_b(FullAdder_455_io_b),
    .io_ci(FullAdder_455_io_ci),
    .io_s(FullAdder_455_io_s),
    .io_co(FullAdder_455_io_co)
  );
  FullAdder FullAdder_456 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_456_io_a),
    .io_b(FullAdder_456_io_b),
    .io_ci(FullAdder_456_io_ci),
    .io_s(FullAdder_456_io_s),
    .io_co(FullAdder_456_io_co)
  );
  FullAdder FullAdder_457 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_457_io_a),
    .io_b(FullAdder_457_io_b),
    .io_ci(FullAdder_457_io_ci),
    .io_s(FullAdder_457_io_s),
    .io_co(FullAdder_457_io_co)
  );
  FullAdder FullAdder_458 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_458_io_a),
    .io_b(FullAdder_458_io_b),
    .io_ci(FullAdder_458_io_ci),
    .io_s(FullAdder_458_io_s),
    .io_co(FullAdder_458_io_co)
  );
  FullAdder FullAdder_459 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_459_io_a),
    .io_b(FullAdder_459_io_b),
    .io_ci(FullAdder_459_io_ci),
    .io_s(FullAdder_459_io_s),
    .io_co(FullAdder_459_io_co)
  );
  FullAdder FullAdder_460 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_460_io_a),
    .io_b(FullAdder_460_io_b),
    .io_ci(FullAdder_460_io_ci),
    .io_s(FullAdder_460_io_s),
    .io_co(FullAdder_460_io_co)
  );
  FullAdder FullAdder_461 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_461_io_a),
    .io_b(FullAdder_461_io_b),
    .io_ci(FullAdder_461_io_ci),
    .io_s(FullAdder_461_io_s),
    .io_co(FullAdder_461_io_co)
  );
  FullAdder FullAdder_462 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_462_io_a),
    .io_b(FullAdder_462_io_b),
    .io_ci(FullAdder_462_io_ci),
    .io_s(FullAdder_462_io_s),
    .io_co(FullAdder_462_io_co)
  );
  FullAdder FullAdder_463 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_463_io_a),
    .io_b(FullAdder_463_io_b),
    .io_ci(FullAdder_463_io_ci),
    .io_s(FullAdder_463_io_s),
    .io_co(FullAdder_463_io_co)
  );
  FullAdder FullAdder_464 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_464_io_a),
    .io_b(FullAdder_464_io_b),
    .io_ci(FullAdder_464_io_ci),
    .io_s(FullAdder_464_io_s),
    .io_co(FullAdder_464_io_co)
  );
  FullAdder FullAdder_465 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_465_io_a),
    .io_b(FullAdder_465_io_b),
    .io_ci(FullAdder_465_io_ci),
    .io_s(FullAdder_465_io_s),
    .io_co(FullAdder_465_io_co)
  );
  FullAdder FullAdder_466 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_466_io_a),
    .io_b(FullAdder_466_io_b),
    .io_ci(FullAdder_466_io_ci),
    .io_s(FullAdder_466_io_s),
    .io_co(FullAdder_466_io_co)
  );
  HalfAdder HalfAdder_25 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_25_io_a),
    .io_b(HalfAdder_25_io_b),
    .io_s(HalfAdder_25_io_s),
    .io_co(HalfAdder_25_io_co)
  );
  FullAdder FullAdder_467 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_467_io_a),
    .io_b(FullAdder_467_io_b),
    .io_ci(FullAdder_467_io_ci),
    .io_s(FullAdder_467_io_s),
    .io_co(FullAdder_467_io_co)
  );
  FullAdder FullAdder_468 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_468_io_a),
    .io_b(FullAdder_468_io_b),
    .io_ci(FullAdder_468_io_ci),
    .io_s(FullAdder_468_io_s),
    .io_co(FullAdder_468_io_co)
  );
  FullAdder FullAdder_469 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_469_io_a),
    .io_b(FullAdder_469_io_b),
    .io_ci(FullAdder_469_io_ci),
    .io_s(FullAdder_469_io_s),
    .io_co(FullAdder_469_io_co)
  );
  FullAdder FullAdder_470 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_470_io_a),
    .io_b(FullAdder_470_io_b),
    .io_ci(FullAdder_470_io_ci),
    .io_s(FullAdder_470_io_s),
    .io_co(FullAdder_470_io_co)
  );
  FullAdder FullAdder_471 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_471_io_a),
    .io_b(FullAdder_471_io_b),
    .io_ci(FullAdder_471_io_ci),
    .io_s(FullAdder_471_io_s),
    .io_co(FullAdder_471_io_co)
  );
  HalfAdder HalfAdder_26 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_26_io_a),
    .io_b(HalfAdder_26_io_b),
    .io_s(HalfAdder_26_io_s),
    .io_co(HalfAdder_26_io_co)
  );
  FullAdder FullAdder_472 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_472_io_a),
    .io_b(FullAdder_472_io_b),
    .io_ci(FullAdder_472_io_ci),
    .io_s(FullAdder_472_io_s),
    .io_co(FullAdder_472_io_co)
  );
  FullAdder FullAdder_473 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_473_io_a),
    .io_b(FullAdder_473_io_b),
    .io_ci(FullAdder_473_io_ci),
    .io_s(FullAdder_473_io_s),
    .io_co(FullAdder_473_io_co)
  );
  FullAdder FullAdder_474 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_474_io_a),
    .io_b(FullAdder_474_io_b),
    .io_ci(FullAdder_474_io_ci),
    .io_s(FullAdder_474_io_s),
    .io_co(FullAdder_474_io_co)
  );
  FullAdder FullAdder_475 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_475_io_a),
    .io_b(FullAdder_475_io_b),
    .io_ci(FullAdder_475_io_ci),
    .io_s(FullAdder_475_io_s),
    .io_co(FullAdder_475_io_co)
  );
  FullAdder FullAdder_476 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_476_io_a),
    .io_b(FullAdder_476_io_b),
    .io_ci(FullAdder_476_io_ci),
    .io_s(FullAdder_476_io_s),
    .io_co(FullAdder_476_io_co)
  );
  FullAdder FullAdder_477 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_477_io_a),
    .io_b(FullAdder_477_io_b),
    .io_ci(FullAdder_477_io_ci),
    .io_s(FullAdder_477_io_s),
    .io_co(FullAdder_477_io_co)
  );
  FullAdder FullAdder_478 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_478_io_a),
    .io_b(FullAdder_478_io_b),
    .io_ci(FullAdder_478_io_ci),
    .io_s(FullAdder_478_io_s),
    .io_co(FullAdder_478_io_co)
  );
  FullAdder FullAdder_479 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_479_io_a),
    .io_b(FullAdder_479_io_b),
    .io_ci(FullAdder_479_io_ci),
    .io_s(FullAdder_479_io_s),
    .io_co(FullAdder_479_io_co)
  );
  FullAdder FullAdder_480 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_480_io_a),
    .io_b(FullAdder_480_io_b),
    .io_ci(FullAdder_480_io_ci),
    .io_s(FullAdder_480_io_s),
    .io_co(FullAdder_480_io_co)
  );
  FullAdder FullAdder_481 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_481_io_a),
    .io_b(FullAdder_481_io_b),
    .io_ci(FullAdder_481_io_ci),
    .io_s(FullAdder_481_io_s),
    .io_co(FullAdder_481_io_co)
  );
  FullAdder FullAdder_482 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_482_io_a),
    .io_b(FullAdder_482_io_b),
    .io_ci(FullAdder_482_io_ci),
    .io_s(FullAdder_482_io_s),
    .io_co(FullAdder_482_io_co)
  );
  FullAdder FullAdder_483 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_483_io_a),
    .io_b(FullAdder_483_io_b),
    .io_ci(FullAdder_483_io_ci),
    .io_s(FullAdder_483_io_s),
    .io_co(FullAdder_483_io_co)
  );
  FullAdder FullAdder_484 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_484_io_a),
    .io_b(FullAdder_484_io_b),
    .io_ci(FullAdder_484_io_ci),
    .io_s(FullAdder_484_io_s),
    .io_co(FullAdder_484_io_co)
  );
  FullAdder FullAdder_485 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_485_io_a),
    .io_b(FullAdder_485_io_b),
    .io_ci(FullAdder_485_io_ci),
    .io_s(FullAdder_485_io_s),
    .io_co(FullAdder_485_io_co)
  );
  FullAdder FullAdder_486 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_486_io_a),
    .io_b(FullAdder_486_io_b),
    .io_ci(FullAdder_486_io_ci),
    .io_s(FullAdder_486_io_s),
    .io_co(FullAdder_486_io_co)
  );
  FullAdder FullAdder_487 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_487_io_a),
    .io_b(FullAdder_487_io_b),
    .io_ci(FullAdder_487_io_ci),
    .io_s(FullAdder_487_io_s),
    .io_co(FullAdder_487_io_co)
  );
  FullAdder FullAdder_488 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_488_io_a),
    .io_b(FullAdder_488_io_b),
    .io_ci(FullAdder_488_io_ci),
    .io_s(FullAdder_488_io_s),
    .io_co(FullAdder_488_io_co)
  );
  FullAdder FullAdder_489 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_489_io_a),
    .io_b(FullAdder_489_io_b),
    .io_ci(FullAdder_489_io_ci),
    .io_s(FullAdder_489_io_s),
    .io_co(FullAdder_489_io_co)
  );
  FullAdder FullAdder_490 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_490_io_a),
    .io_b(FullAdder_490_io_b),
    .io_ci(FullAdder_490_io_ci),
    .io_s(FullAdder_490_io_s),
    .io_co(FullAdder_490_io_co)
  );
  FullAdder FullAdder_491 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_491_io_a),
    .io_b(FullAdder_491_io_b),
    .io_ci(FullAdder_491_io_ci),
    .io_s(FullAdder_491_io_s),
    .io_co(FullAdder_491_io_co)
  );
  FullAdder FullAdder_492 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_492_io_a),
    .io_b(FullAdder_492_io_b),
    .io_ci(FullAdder_492_io_ci),
    .io_s(FullAdder_492_io_s),
    .io_co(FullAdder_492_io_co)
  );
  FullAdder FullAdder_493 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_493_io_a),
    .io_b(FullAdder_493_io_b),
    .io_ci(FullAdder_493_io_ci),
    .io_s(FullAdder_493_io_s),
    .io_co(FullAdder_493_io_co)
  );
  FullAdder FullAdder_494 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_494_io_a),
    .io_b(FullAdder_494_io_b),
    .io_ci(FullAdder_494_io_ci),
    .io_s(FullAdder_494_io_s),
    .io_co(FullAdder_494_io_co)
  );
  FullAdder FullAdder_495 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_495_io_a),
    .io_b(FullAdder_495_io_b),
    .io_ci(FullAdder_495_io_ci),
    .io_s(FullAdder_495_io_s),
    .io_co(FullAdder_495_io_co)
  );
  FullAdder FullAdder_496 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_496_io_a),
    .io_b(FullAdder_496_io_b),
    .io_ci(FullAdder_496_io_ci),
    .io_s(FullAdder_496_io_s),
    .io_co(FullAdder_496_io_co)
  );
  FullAdder FullAdder_497 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_497_io_a),
    .io_b(FullAdder_497_io_b),
    .io_ci(FullAdder_497_io_ci),
    .io_s(FullAdder_497_io_s),
    .io_co(FullAdder_497_io_co)
  );
  FullAdder FullAdder_498 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_498_io_a),
    .io_b(FullAdder_498_io_b),
    .io_ci(FullAdder_498_io_ci),
    .io_s(FullAdder_498_io_s),
    .io_co(FullAdder_498_io_co)
  );
  FullAdder FullAdder_499 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_499_io_a),
    .io_b(FullAdder_499_io_b),
    .io_ci(FullAdder_499_io_ci),
    .io_s(FullAdder_499_io_s),
    .io_co(FullAdder_499_io_co)
  );
  FullAdder FullAdder_500 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_500_io_a),
    .io_b(FullAdder_500_io_b),
    .io_ci(FullAdder_500_io_ci),
    .io_s(FullAdder_500_io_s),
    .io_co(FullAdder_500_io_co)
  );
  FullAdder FullAdder_501 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_501_io_a),
    .io_b(FullAdder_501_io_b),
    .io_ci(FullAdder_501_io_ci),
    .io_s(FullAdder_501_io_s),
    .io_co(FullAdder_501_io_co)
  );
  FullAdder FullAdder_502 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_502_io_a),
    .io_b(FullAdder_502_io_b),
    .io_ci(FullAdder_502_io_ci),
    .io_s(FullAdder_502_io_s),
    .io_co(FullAdder_502_io_co)
  );
  FullAdder FullAdder_503 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_503_io_a),
    .io_b(FullAdder_503_io_b),
    .io_ci(FullAdder_503_io_ci),
    .io_s(FullAdder_503_io_s),
    .io_co(FullAdder_503_io_co)
  );
  FullAdder FullAdder_504 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_504_io_a),
    .io_b(FullAdder_504_io_b),
    .io_ci(FullAdder_504_io_ci),
    .io_s(FullAdder_504_io_s),
    .io_co(FullAdder_504_io_co)
  );
  FullAdder FullAdder_505 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_505_io_a),
    .io_b(FullAdder_505_io_b),
    .io_ci(FullAdder_505_io_ci),
    .io_s(FullAdder_505_io_s),
    .io_co(FullAdder_505_io_co)
  );
  HalfAdder HalfAdder_27 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_27_io_a),
    .io_b(HalfAdder_27_io_b),
    .io_s(HalfAdder_27_io_s),
    .io_co(HalfAdder_27_io_co)
  );
  FullAdder FullAdder_506 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_506_io_a),
    .io_b(FullAdder_506_io_b),
    .io_ci(FullAdder_506_io_ci),
    .io_s(FullAdder_506_io_s),
    .io_co(FullAdder_506_io_co)
  );
  FullAdder FullAdder_507 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_507_io_a),
    .io_b(FullAdder_507_io_b),
    .io_ci(FullAdder_507_io_ci),
    .io_s(FullAdder_507_io_s),
    .io_co(FullAdder_507_io_co)
  );
  FullAdder FullAdder_508 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_508_io_a),
    .io_b(FullAdder_508_io_b),
    .io_ci(FullAdder_508_io_ci),
    .io_s(FullAdder_508_io_s),
    .io_co(FullAdder_508_io_co)
  );
  FullAdder FullAdder_509 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_509_io_a),
    .io_b(FullAdder_509_io_b),
    .io_ci(FullAdder_509_io_ci),
    .io_s(FullAdder_509_io_s),
    .io_co(FullAdder_509_io_co)
  );
  FullAdder FullAdder_510 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_510_io_a),
    .io_b(FullAdder_510_io_b),
    .io_ci(FullAdder_510_io_ci),
    .io_s(FullAdder_510_io_s),
    .io_co(FullAdder_510_io_co)
  );
  FullAdder FullAdder_511 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_511_io_a),
    .io_b(FullAdder_511_io_b),
    .io_ci(FullAdder_511_io_ci),
    .io_s(FullAdder_511_io_s),
    .io_co(FullAdder_511_io_co)
  );
  FullAdder FullAdder_512 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_512_io_a),
    .io_b(FullAdder_512_io_b),
    .io_ci(FullAdder_512_io_ci),
    .io_s(FullAdder_512_io_s),
    .io_co(FullAdder_512_io_co)
  );
  FullAdder FullAdder_513 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_513_io_a),
    .io_b(FullAdder_513_io_b),
    .io_ci(FullAdder_513_io_ci),
    .io_s(FullAdder_513_io_s),
    .io_co(FullAdder_513_io_co)
  );
  FullAdder FullAdder_514 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_514_io_a),
    .io_b(FullAdder_514_io_b),
    .io_ci(FullAdder_514_io_ci),
    .io_s(FullAdder_514_io_s),
    .io_co(FullAdder_514_io_co)
  );
  FullAdder FullAdder_515 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_515_io_a),
    .io_b(FullAdder_515_io_b),
    .io_ci(FullAdder_515_io_ci),
    .io_s(FullAdder_515_io_s),
    .io_co(FullAdder_515_io_co)
  );
  FullAdder FullAdder_516 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_516_io_a),
    .io_b(FullAdder_516_io_b),
    .io_ci(FullAdder_516_io_ci),
    .io_s(FullAdder_516_io_s),
    .io_co(FullAdder_516_io_co)
  );
  FullAdder FullAdder_517 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_517_io_a),
    .io_b(FullAdder_517_io_b),
    .io_ci(FullAdder_517_io_ci),
    .io_s(FullAdder_517_io_s),
    .io_co(FullAdder_517_io_co)
  );
  FullAdder FullAdder_518 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_518_io_a),
    .io_b(FullAdder_518_io_b),
    .io_ci(FullAdder_518_io_ci),
    .io_s(FullAdder_518_io_s),
    .io_co(FullAdder_518_io_co)
  );
  FullAdder FullAdder_519 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_519_io_a),
    .io_b(FullAdder_519_io_b),
    .io_ci(FullAdder_519_io_ci),
    .io_s(FullAdder_519_io_s),
    .io_co(FullAdder_519_io_co)
  );
  HalfAdder HalfAdder_28 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_28_io_a),
    .io_b(HalfAdder_28_io_b),
    .io_s(HalfAdder_28_io_s),
    .io_co(HalfAdder_28_io_co)
  );
  FullAdder FullAdder_520 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_520_io_a),
    .io_b(FullAdder_520_io_b),
    .io_ci(FullAdder_520_io_ci),
    .io_s(FullAdder_520_io_s),
    .io_co(FullAdder_520_io_co)
  );
  FullAdder FullAdder_521 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_521_io_a),
    .io_b(FullAdder_521_io_b),
    .io_ci(FullAdder_521_io_ci),
    .io_s(FullAdder_521_io_s),
    .io_co(FullAdder_521_io_co)
  );
  FullAdder FullAdder_522 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_522_io_a),
    .io_b(FullAdder_522_io_b),
    .io_ci(FullAdder_522_io_ci),
    .io_s(FullAdder_522_io_s),
    .io_co(FullAdder_522_io_co)
  );
  FullAdder FullAdder_523 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_523_io_a),
    .io_b(FullAdder_523_io_b),
    .io_ci(FullAdder_523_io_ci),
    .io_s(FullAdder_523_io_s),
    .io_co(FullAdder_523_io_co)
  );
  FullAdder FullAdder_524 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_524_io_a),
    .io_b(FullAdder_524_io_b),
    .io_ci(FullAdder_524_io_ci),
    .io_s(FullAdder_524_io_s),
    .io_co(FullAdder_524_io_co)
  );
  FullAdder FullAdder_525 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_525_io_a),
    .io_b(FullAdder_525_io_b),
    .io_ci(FullAdder_525_io_ci),
    .io_s(FullAdder_525_io_s),
    .io_co(FullAdder_525_io_co)
  );
  FullAdder FullAdder_526 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_526_io_a),
    .io_b(FullAdder_526_io_b),
    .io_ci(FullAdder_526_io_ci),
    .io_s(FullAdder_526_io_s),
    .io_co(FullAdder_526_io_co)
  );
  HalfAdder HalfAdder_29 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_29_io_a),
    .io_b(HalfAdder_29_io_b),
    .io_s(HalfAdder_29_io_s),
    .io_co(HalfAdder_29_io_co)
  );
  FullAdder FullAdder_527 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_527_io_a),
    .io_b(FullAdder_527_io_b),
    .io_ci(FullAdder_527_io_ci),
    .io_s(FullAdder_527_io_s),
    .io_co(FullAdder_527_io_co)
  );
  HalfAdder HalfAdder_30 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_30_io_a),
    .io_b(HalfAdder_30_io_b),
    .io_s(HalfAdder_30_io_s),
    .io_co(HalfAdder_30_io_co)
  );
  HalfAdder HalfAdder_31 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_31_io_a),
    .io_b(HalfAdder_31_io_b),
    .io_s(HalfAdder_31_io_s),
    .io_co(HalfAdder_31_io_co)
  );
  HalfAdder HalfAdder_32 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_32_io_a),
    .io_b(HalfAdder_32_io_b),
    .io_s(HalfAdder_32_io_s),
    .io_co(HalfAdder_32_io_co)
  );
  HalfAdder HalfAdder_33 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_33_io_a),
    .io_b(HalfAdder_33_io_b),
    .io_s(HalfAdder_33_io_s),
    .io_co(HalfAdder_33_io_co)
  );
  FullAdder FullAdder_528 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_528_io_a),
    .io_b(FullAdder_528_io_b),
    .io_ci(FullAdder_528_io_ci),
    .io_s(FullAdder_528_io_s),
    .io_co(FullAdder_528_io_co)
  );
  HalfAdder HalfAdder_34 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_34_io_a),
    .io_b(HalfAdder_34_io_b),
    .io_s(HalfAdder_34_io_s),
    .io_co(HalfAdder_34_io_co)
  );
  HalfAdder HalfAdder_35 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_35_io_a),
    .io_b(HalfAdder_35_io_b),
    .io_s(HalfAdder_35_io_s),
    .io_co(HalfAdder_35_io_co)
  );
  HalfAdder HalfAdder_36 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_36_io_a),
    .io_b(HalfAdder_36_io_b),
    .io_s(HalfAdder_36_io_s),
    .io_co(HalfAdder_36_io_co)
  );
  FullAdder FullAdder_529 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_529_io_a),
    .io_b(FullAdder_529_io_b),
    .io_ci(FullAdder_529_io_ci),
    .io_s(FullAdder_529_io_s),
    .io_co(FullAdder_529_io_co)
  );
  FullAdder FullAdder_530 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_530_io_a),
    .io_b(FullAdder_530_io_b),
    .io_ci(FullAdder_530_io_ci),
    .io_s(FullAdder_530_io_s),
    .io_co(FullAdder_530_io_co)
  );
  FullAdder FullAdder_531 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_531_io_a),
    .io_b(FullAdder_531_io_b),
    .io_ci(FullAdder_531_io_ci),
    .io_s(FullAdder_531_io_s),
    .io_co(FullAdder_531_io_co)
  );
  FullAdder FullAdder_532 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_532_io_a),
    .io_b(FullAdder_532_io_b),
    .io_ci(FullAdder_532_io_ci),
    .io_s(FullAdder_532_io_s),
    .io_co(FullAdder_532_io_co)
  );
  FullAdder FullAdder_533 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_533_io_a),
    .io_b(FullAdder_533_io_b),
    .io_ci(FullAdder_533_io_ci),
    .io_s(FullAdder_533_io_s),
    .io_co(FullAdder_533_io_co)
  );
  FullAdder FullAdder_534 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_534_io_a),
    .io_b(FullAdder_534_io_b),
    .io_ci(FullAdder_534_io_ci),
    .io_s(FullAdder_534_io_s),
    .io_co(FullAdder_534_io_co)
  );
  HalfAdder HalfAdder_37 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_37_io_a),
    .io_b(HalfAdder_37_io_b),
    .io_s(HalfAdder_37_io_s),
    .io_co(HalfAdder_37_io_co)
  );
  FullAdder FullAdder_535 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_535_io_a),
    .io_b(FullAdder_535_io_b),
    .io_ci(FullAdder_535_io_ci),
    .io_s(FullAdder_535_io_s),
    .io_co(FullAdder_535_io_co)
  );
  FullAdder FullAdder_536 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_536_io_a),
    .io_b(FullAdder_536_io_b),
    .io_ci(FullAdder_536_io_ci),
    .io_s(FullAdder_536_io_s),
    .io_co(FullAdder_536_io_co)
  );
  FullAdder FullAdder_537 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_537_io_a),
    .io_b(FullAdder_537_io_b),
    .io_ci(FullAdder_537_io_ci),
    .io_s(FullAdder_537_io_s),
    .io_co(FullAdder_537_io_co)
  );
  FullAdder FullAdder_538 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_538_io_a),
    .io_b(FullAdder_538_io_b),
    .io_ci(FullAdder_538_io_ci),
    .io_s(FullAdder_538_io_s),
    .io_co(FullAdder_538_io_co)
  );
  FullAdder FullAdder_539 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_539_io_a),
    .io_b(FullAdder_539_io_b),
    .io_ci(FullAdder_539_io_ci),
    .io_s(FullAdder_539_io_s),
    .io_co(FullAdder_539_io_co)
  );
  FullAdder FullAdder_540 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_540_io_a),
    .io_b(FullAdder_540_io_b),
    .io_ci(FullAdder_540_io_ci),
    .io_s(FullAdder_540_io_s),
    .io_co(FullAdder_540_io_co)
  );
  FullAdder FullAdder_541 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_541_io_a),
    .io_b(FullAdder_541_io_b),
    .io_ci(FullAdder_541_io_ci),
    .io_s(FullAdder_541_io_s),
    .io_co(FullAdder_541_io_co)
  );
  FullAdder FullAdder_542 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_542_io_a),
    .io_b(FullAdder_542_io_b),
    .io_ci(FullAdder_542_io_ci),
    .io_s(FullAdder_542_io_s),
    .io_co(FullAdder_542_io_co)
  );
  FullAdder FullAdder_543 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_543_io_a),
    .io_b(FullAdder_543_io_b),
    .io_ci(FullAdder_543_io_ci),
    .io_s(FullAdder_543_io_s),
    .io_co(FullAdder_543_io_co)
  );
  FullAdder FullAdder_544 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_544_io_a),
    .io_b(FullAdder_544_io_b),
    .io_ci(FullAdder_544_io_ci),
    .io_s(FullAdder_544_io_s),
    .io_co(FullAdder_544_io_co)
  );
  FullAdder FullAdder_545 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_545_io_a),
    .io_b(FullAdder_545_io_b),
    .io_ci(FullAdder_545_io_ci),
    .io_s(FullAdder_545_io_s),
    .io_co(FullAdder_545_io_co)
  );
  FullAdder FullAdder_546 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_546_io_a),
    .io_b(FullAdder_546_io_b),
    .io_ci(FullAdder_546_io_ci),
    .io_s(FullAdder_546_io_s),
    .io_co(FullAdder_546_io_co)
  );
  HalfAdder HalfAdder_38 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_38_io_a),
    .io_b(HalfAdder_38_io_b),
    .io_s(HalfAdder_38_io_s),
    .io_co(HalfAdder_38_io_co)
  );
  FullAdder FullAdder_547 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_547_io_a),
    .io_b(FullAdder_547_io_b),
    .io_ci(FullAdder_547_io_ci),
    .io_s(FullAdder_547_io_s),
    .io_co(FullAdder_547_io_co)
  );
  FullAdder FullAdder_548 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_548_io_a),
    .io_b(FullAdder_548_io_b),
    .io_ci(FullAdder_548_io_ci),
    .io_s(FullAdder_548_io_s),
    .io_co(FullAdder_548_io_co)
  );
  HalfAdder HalfAdder_39 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_39_io_a),
    .io_b(HalfAdder_39_io_b),
    .io_s(HalfAdder_39_io_s),
    .io_co(HalfAdder_39_io_co)
  );
  FullAdder FullAdder_549 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_549_io_a),
    .io_b(FullAdder_549_io_b),
    .io_ci(FullAdder_549_io_ci),
    .io_s(FullAdder_549_io_s),
    .io_co(FullAdder_549_io_co)
  );
  FullAdder FullAdder_550 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_550_io_a),
    .io_b(FullAdder_550_io_b),
    .io_ci(FullAdder_550_io_ci),
    .io_s(FullAdder_550_io_s),
    .io_co(FullAdder_550_io_co)
  );
  HalfAdder HalfAdder_40 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_40_io_a),
    .io_b(HalfAdder_40_io_b),
    .io_s(HalfAdder_40_io_s),
    .io_co(HalfAdder_40_io_co)
  );
  FullAdder FullAdder_551 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_551_io_a),
    .io_b(FullAdder_551_io_b),
    .io_ci(FullAdder_551_io_ci),
    .io_s(FullAdder_551_io_s),
    .io_co(FullAdder_551_io_co)
  );
  FullAdder FullAdder_552 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_552_io_a),
    .io_b(FullAdder_552_io_b),
    .io_ci(FullAdder_552_io_ci),
    .io_s(FullAdder_552_io_s),
    .io_co(FullAdder_552_io_co)
  );
  HalfAdder HalfAdder_41 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_41_io_a),
    .io_b(HalfAdder_41_io_b),
    .io_s(HalfAdder_41_io_s),
    .io_co(HalfAdder_41_io_co)
  );
  FullAdder FullAdder_553 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_553_io_a),
    .io_b(FullAdder_553_io_b),
    .io_ci(FullAdder_553_io_ci),
    .io_s(FullAdder_553_io_s),
    .io_co(FullAdder_553_io_co)
  );
  FullAdder FullAdder_554 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_554_io_a),
    .io_b(FullAdder_554_io_b),
    .io_ci(FullAdder_554_io_ci),
    .io_s(FullAdder_554_io_s),
    .io_co(FullAdder_554_io_co)
  );
  FullAdder FullAdder_555 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_555_io_a),
    .io_b(FullAdder_555_io_b),
    .io_ci(FullAdder_555_io_ci),
    .io_s(FullAdder_555_io_s),
    .io_co(FullAdder_555_io_co)
  );
  FullAdder FullAdder_556 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_556_io_a),
    .io_b(FullAdder_556_io_b),
    .io_ci(FullAdder_556_io_ci),
    .io_s(FullAdder_556_io_s),
    .io_co(FullAdder_556_io_co)
  );
  FullAdder FullAdder_557 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_557_io_a),
    .io_b(FullAdder_557_io_b),
    .io_ci(FullAdder_557_io_ci),
    .io_s(FullAdder_557_io_s),
    .io_co(FullAdder_557_io_co)
  );
  FullAdder FullAdder_558 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_558_io_a),
    .io_b(FullAdder_558_io_b),
    .io_ci(FullAdder_558_io_ci),
    .io_s(FullAdder_558_io_s),
    .io_co(FullAdder_558_io_co)
  );
  FullAdder FullAdder_559 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_559_io_a),
    .io_b(FullAdder_559_io_b),
    .io_ci(FullAdder_559_io_ci),
    .io_s(FullAdder_559_io_s),
    .io_co(FullAdder_559_io_co)
  );
  FullAdder FullAdder_560 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_560_io_a),
    .io_b(FullAdder_560_io_b),
    .io_ci(FullAdder_560_io_ci),
    .io_s(FullAdder_560_io_s),
    .io_co(FullAdder_560_io_co)
  );
  FullAdder FullAdder_561 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_561_io_a),
    .io_b(FullAdder_561_io_b),
    .io_ci(FullAdder_561_io_ci),
    .io_s(FullAdder_561_io_s),
    .io_co(FullAdder_561_io_co)
  );
  FullAdder FullAdder_562 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_562_io_a),
    .io_b(FullAdder_562_io_b),
    .io_ci(FullAdder_562_io_ci),
    .io_s(FullAdder_562_io_s),
    .io_co(FullAdder_562_io_co)
  );
  FullAdder FullAdder_563 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_563_io_a),
    .io_b(FullAdder_563_io_b),
    .io_ci(FullAdder_563_io_ci),
    .io_s(FullAdder_563_io_s),
    .io_co(FullAdder_563_io_co)
  );
  FullAdder FullAdder_564 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_564_io_a),
    .io_b(FullAdder_564_io_b),
    .io_ci(FullAdder_564_io_ci),
    .io_s(FullAdder_564_io_s),
    .io_co(FullAdder_564_io_co)
  );
  HalfAdder HalfAdder_42 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_42_io_a),
    .io_b(HalfAdder_42_io_b),
    .io_s(HalfAdder_42_io_s),
    .io_co(HalfAdder_42_io_co)
  );
  FullAdder FullAdder_565 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_565_io_a),
    .io_b(FullAdder_565_io_b),
    .io_ci(FullAdder_565_io_ci),
    .io_s(FullAdder_565_io_s),
    .io_co(FullAdder_565_io_co)
  );
  FullAdder FullAdder_566 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_566_io_a),
    .io_b(FullAdder_566_io_b),
    .io_ci(FullAdder_566_io_ci),
    .io_s(FullAdder_566_io_s),
    .io_co(FullAdder_566_io_co)
  );
  FullAdder FullAdder_567 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_567_io_a),
    .io_b(FullAdder_567_io_b),
    .io_ci(FullAdder_567_io_ci),
    .io_s(FullAdder_567_io_s),
    .io_co(FullAdder_567_io_co)
  );
  HalfAdder HalfAdder_43 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_43_io_a),
    .io_b(HalfAdder_43_io_b),
    .io_s(HalfAdder_43_io_s),
    .io_co(HalfAdder_43_io_co)
  );
  FullAdder FullAdder_568 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_568_io_a),
    .io_b(FullAdder_568_io_b),
    .io_ci(FullAdder_568_io_ci),
    .io_s(FullAdder_568_io_s),
    .io_co(FullAdder_568_io_co)
  );
  FullAdder FullAdder_569 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_569_io_a),
    .io_b(FullAdder_569_io_b),
    .io_ci(FullAdder_569_io_ci),
    .io_s(FullAdder_569_io_s),
    .io_co(FullAdder_569_io_co)
  );
  FullAdder FullAdder_570 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_570_io_a),
    .io_b(FullAdder_570_io_b),
    .io_ci(FullAdder_570_io_ci),
    .io_s(FullAdder_570_io_s),
    .io_co(FullAdder_570_io_co)
  );
  FullAdder FullAdder_571 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_571_io_a),
    .io_b(FullAdder_571_io_b),
    .io_ci(FullAdder_571_io_ci),
    .io_s(FullAdder_571_io_s),
    .io_co(FullAdder_571_io_co)
  );
  FullAdder FullAdder_572 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_572_io_a),
    .io_b(FullAdder_572_io_b),
    .io_ci(FullAdder_572_io_ci),
    .io_s(FullAdder_572_io_s),
    .io_co(FullAdder_572_io_co)
  );
  FullAdder FullAdder_573 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_573_io_a),
    .io_b(FullAdder_573_io_b),
    .io_ci(FullAdder_573_io_ci),
    .io_s(FullAdder_573_io_s),
    .io_co(FullAdder_573_io_co)
  );
  FullAdder FullAdder_574 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_574_io_a),
    .io_b(FullAdder_574_io_b),
    .io_ci(FullAdder_574_io_ci),
    .io_s(FullAdder_574_io_s),
    .io_co(FullAdder_574_io_co)
  );
  FullAdder FullAdder_575 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_575_io_a),
    .io_b(FullAdder_575_io_b),
    .io_ci(FullAdder_575_io_ci),
    .io_s(FullAdder_575_io_s),
    .io_co(FullAdder_575_io_co)
  );
  FullAdder FullAdder_576 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_576_io_a),
    .io_b(FullAdder_576_io_b),
    .io_ci(FullAdder_576_io_ci),
    .io_s(FullAdder_576_io_s),
    .io_co(FullAdder_576_io_co)
  );
  FullAdder FullAdder_577 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_577_io_a),
    .io_b(FullAdder_577_io_b),
    .io_ci(FullAdder_577_io_ci),
    .io_s(FullAdder_577_io_s),
    .io_co(FullAdder_577_io_co)
  );
  FullAdder FullAdder_578 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_578_io_a),
    .io_b(FullAdder_578_io_b),
    .io_ci(FullAdder_578_io_ci),
    .io_s(FullAdder_578_io_s),
    .io_co(FullAdder_578_io_co)
  );
  FullAdder FullAdder_579 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_579_io_a),
    .io_b(FullAdder_579_io_b),
    .io_ci(FullAdder_579_io_ci),
    .io_s(FullAdder_579_io_s),
    .io_co(FullAdder_579_io_co)
  );
  FullAdder FullAdder_580 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_580_io_a),
    .io_b(FullAdder_580_io_b),
    .io_ci(FullAdder_580_io_ci),
    .io_s(FullAdder_580_io_s),
    .io_co(FullAdder_580_io_co)
  );
  FullAdder FullAdder_581 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_581_io_a),
    .io_b(FullAdder_581_io_b),
    .io_ci(FullAdder_581_io_ci),
    .io_s(FullAdder_581_io_s),
    .io_co(FullAdder_581_io_co)
  );
  FullAdder FullAdder_582 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_582_io_a),
    .io_b(FullAdder_582_io_b),
    .io_ci(FullAdder_582_io_ci),
    .io_s(FullAdder_582_io_s),
    .io_co(FullAdder_582_io_co)
  );
  FullAdder FullAdder_583 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_583_io_a),
    .io_b(FullAdder_583_io_b),
    .io_ci(FullAdder_583_io_ci),
    .io_s(FullAdder_583_io_s),
    .io_co(FullAdder_583_io_co)
  );
  FullAdder FullAdder_584 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_584_io_a),
    .io_b(FullAdder_584_io_b),
    .io_ci(FullAdder_584_io_ci),
    .io_s(FullAdder_584_io_s),
    .io_co(FullAdder_584_io_co)
  );
  FullAdder FullAdder_585 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_585_io_a),
    .io_b(FullAdder_585_io_b),
    .io_ci(FullAdder_585_io_ci),
    .io_s(FullAdder_585_io_s),
    .io_co(FullAdder_585_io_co)
  );
  FullAdder FullAdder_586 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_586_io_a),
    .io_b(FullAdder_586_io_b),
    .io_ci(FullAdder_586_io_ci),
    .io_s(FullAdder_586_io_s),
    .io_co(FullAdder_586_io_co)
  );
  FullAdder FullAdder_587 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_587_io_a),
    .io_b(FullAdder_587_io_b),
    .io_ci(FullAdder_587_io_ci),
    .io_s(FullAdder_587_io_s),
    .io_co(FullAdder_587_io_co)
  );
  HalfAdder HalfAdder_44 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_44_io_a),
    .io_b(HalfAdder_44_io_b),
    .io_s(HalfAdder_44_io_s),
    .io_co(HalfAdder_44_io_co)
  );
  FullAdder FullAdder_588 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_588_io_a),
    .io_b(FullAdder_588_io_b),
    .io_ci(FullAdder_588_io_ci),
    .io_s(FullAdder_588_io_s),
    .io_co(FullAdder_588_io_co)
  );
  FullAdder FullAdder_589 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_589_io_a),
    .io_b(FullAdder_589_io_b),
    .io_ci(FullAdder_589_io_ci),
    .io_s(FullAdder_589_io_s),
    .io_co(FullAdder_589_io_co)
  );
  FullAdder FullAdder_590 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_590_io_a),
    .io_b(FullAdder_590_io_b),
    .io_ci(FullAdder_590_io_ci),
    .io_s(FullAdder_590_io_s),
    .io_co(FullAdder_590_io_co)
  );
  FullAdder FullAdder_591 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_591_io_a),
    .io_b(FullAdder_591_io_b),
    .io_ci(FullAdder_591_io_ci),
    .io_s(FullAdder_591_io_s),
    .io_co(FullAdder_591_io_co)
  );
  FullAdder FullAdder_592 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_592_io_a),
    .io_b(FullAdder_592_io_b),
    .io_ci(FullAdder_592_io_ci),
    .io_s(FullAdder_592_io_s),
    .io_co(FullAdder_592_io_co)
  );
  FullAdder FullAdder_593 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_593_io_a),
    .io_b(FullAdder_593_io_b),
    .io_ci(FullAdder_593_io_ci),
    .io_s(FullAdder_593_io_s),
    .io_co(FullAdder_593_io_co)
  );
  FullAdder FullAdder_594 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_594_io_a),
    .io_b(FullAdder_594_io_b),
    .io_ci(FullAdder_594_io_ci),
    .io_s(FullAdder_594_io_s),
    .io_co(FullAdder_594_io_co)
  );
  FullAdder FullAdder_595 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_595_io_a),
    .io_b(FullAdder_595_io_b),
    .io_ci(FullAdder_595_io_ci),
    .io_s(FullAdder_595_io_s),
    .io_co(FullAdder_595_io_co)
  );
  FullAdder FullAdder_596 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_596_io_a),
    .io_b(FullAdder_596_io_b),
    .io_ci(FullAdder_596_io_ci),
    .io_s(FullAdder_596_io_s),
    .io_co(FullAdder_596_io_co)
  );
  FullAdder FullAdder_597 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_597_io_a),
    .io_b(FullAdder_597_io_b),
    .io_ci(FullAdder_597_io_ci),
    .io_s(FullAdder_597_io_s),
    .io_co(FullAdder_597_io_co)
  );
  FullAdder FullAdder_598 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_598_io_a),
    .io_b(FullAdder_598_io_b),
    .io_ci(FullAdder_598_io_ci),
    .io_s(FullAdder_598_io_s),
    .io_co(FullAdder_598_io_co)
  );
  FullAdder FullAdder_599 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_599_io_a),
    .io_b(FullAdder_599_io_b),
    .io_ci(FullAdder_599_io_ci),
    .io_s(FullAdder_599_io_s),
    .io_co(FullAdder_599_io_co)
  );
  FullAdder FullAdder_600 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_600_io_a),
    .io_b(FullAdder_600_io_b),
    .io_ci(FullAdder_600_io_ci),
    .io_s(FullAdder_600_io_s),
    .io_co(FullAdder_600_io_co)
  );
  HalfAdder HalfAdder_45 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_45_io_a),
    .io_b(HalfAdder_45_io_b),
    .io_s(HalfAdder_45_io_s),
    .io_co(HalfAdder_45_io_co)
  );
  FullAdder FullAdder_601 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_601_io_a),
    .io_b(FullAdder_601_io_b),
    .io_ci(FullAdder_601_io_ci),
    .io_s(FullAdder_601_io_s),
    .io_co(FullAdder_601_io_co)
  );
  FullAdder FullAdder_602 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_602_io_a),
    .io_b(FullAdder_602_io_b),
    .io_ci(FullAdder_602_io_ci),
    .io_s(FullAdder_602_io_s),
    .io_co(FullAdder_602_io_co)
  );
  FullAdder FullAdder_603 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_603_io_a),
    .io_b(FullAdder_603_io_b),
    .io_ci(FullAdder_603_io_ci),
    .io_s(FullAdder_603_io_s),
    .io_co(FullAdder_603_io_co)
  );
  FullAdder FullAdder_604 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_604_io_a),
    .io_b(FullAdder_604_io_b),
    .io_ci(FullAdder_604_io_ci),
    .io_s(FullAdder_604_io_s),
    .io_co(FullAdder_604_io_co)
  );
  FullAdder FullAdder_605 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_605_io_a),
    .io_b(FullAdder_605_io_b),
    .io_ci(FullAdder_605_io_ci),
    .io_s(FullAdder_605_io_s),
    .io_co(FullAdder_605_io_co)
  );
  FullAdder FullAdder_606 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_606_io_a),
    .io_b(FullAdder_606_io_b),
    .io_ci(FullAdder_606_io_ci),
    .io_s(FullAdder_606_io_s),
    .io_co(FullAdder_606_io_co)
  );
  FullAdder FullAdder_607 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_607_io_a),
    .io_b(FullAdder_607_io_b),
    .io_ci(FullAdder_607_io_ci),
    .io_s(FullAdder_607_io_s),
    .io_co(FullAdder_607_io_co)
  );
  FullAdder FullAdder_608 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_608_io_a),
    .io_b(FullAdder_608_io_b),
    .io_ci(FullAdder_608_io_ci),
    .io_s(FullAdder_608_io_s),
    .io_co(FullAdder_608_io_co)
  );
  FullAdder FullAdder_609 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_609_io_a),
    .io_b(FullAdder_609_io_b),
    .io_ci(FullAdder_609_io_ci),
    .io_s(FullAdder_609_io_s),
    .io_co(FullAdder_609_io_co)
  );
  FullAdder FullAdder_610 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_610_io_a),
    .io_b(FullAdder_610_io_b),
    .io_ci(FullAdder_610_io_ci),
    .io_s(FullAdder_610_io_s),
    .io_co(FullAdder_610_io_co)
  );
  FullAdder FullAdder_611 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_611_io_a),
    .io_b(FullAdder_611_io_b),
    .io_ci(FullAdder_611_io_ci),
    .io_s(FullAdder_611_io_s),
    .io_co(FullAdder_611_io_co)
  );
  FullAdder FullAdder_612 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_612_io_a),
    .io_b(FullAdder_612_io_b),
    .io_ci(FullAdder_612_io_ci),
    .io_s(FullAdder_612_io_s),
    .io_co(FullAdder_612_io_co)
  );
  FullAdder FullAdder_613 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_613_io_a),
    .io_b(FullAdder_613_io_b),
    .io_ci(FullAdder_613_io_ci),
    .io_s(FullAdder_613_io_s),
    .io_co(FullAdder_613_io_co)
  );
  FullAdder FullAdder_614 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_614_io_a),
    .io_b(FullAdder_614_io_b),
    .io_ci(FullAdder_614_io_ci),
    .io_s(FullAdder_614_io_s),
    .io_co(FullAdder_614_io_co)
  );
  FullAdder FullAdder_615 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_615_io_a),
    .io_b(FullAdder_615_io_b),
    .io_ci(FullAdder_615_io_ci),
    .io_s(FullAdder_615_io_s),
    .io_co(FullAdder_615_io_co)
  );
  FullAdder FullAdder_616 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_616_io_a),
    .io_b(FullAdder_616_io_b),
    .io_ci(FullAdder_616_io_ci),
    .io_s(FullAdder_616_io_s),
    .io_co(FullAdder_616_io_co)
  );
  FullAdder FullAdder_617 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_617_io_a),
    .io_b(FullAdder_617_io_b),
    .io_ci(FullAdder_617_io_ci),
    .io_s(FullAdder_617_io_s),
    .io_co(FullAdder_617_io_co)
  );
  FullAdder FullAdder_618 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_618_io_a),
    .io_b(FullAdder_618_io_b),
    .io_ci(FullAdder_618_io_ci),
    .io_s(FullAdder_618_io_s),
    .io_co(FullAdder_618_io_co)
  );
  FullAdder FullAdder_619 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_619_io_a),
    .io_b(FullAdder_619_io_b),
    .io_ci(FullAdder_619_io_ci),
    .io_s(FullAdder_619_io_s),
    .io_co(FullAdder_619_io_co)
  );
  FullAdder FullAdder_620 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_620_io_a),
    .io_b(FullAdder_620_io_b),
    .io_ci(FullAdder_620_io_ci),
    .io_s(FullAdder_620_io_s),
    .io_co(FullAdder_620_io_co)
  );
  FullAdder FullAdder_621 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_621_io_a),
    .io_b(FullAdder_621_io_b),
    .io_ci(FullAdder_621_io_ci),
    .io_s(FullAdder_621_io_s),
    .io_co(FullAdder_621_io_co)
  );
  FullAdder FullAdder_622 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_622_io_a),
    .io_b(FullAdder_622_io_b),
    .io_ci(FullAdder_622_io_ci),
    .io_s(FullAdder_622_io_s),
    .io_co(FullAdder_622_io_co)
  );
  FullAdder FullAdder_623 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_623_io_a),
    .io_b(FullAdder_623_io_b),
    .io_ci(FullAdder_623_io_ci),
    .io_s(FullAdder_623_io_s),
    .io_co(FullAdder_623_io_co)
  );
  FullAdder FullAdder_624 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_624_io_a),
    .io_b(FullAdder_624_io_b),
    .io_ci(FullAdder_624_io_ci),
    .io_s(FullAdder_624_io_s),
    .io_co(FullAdder_624_io_co)
  );
  FullAdder FullAdder_625 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_625_io_a),
    .io_b(FullAdder_625_io_b),
    .io_ci(FullAdder_625_io_ci),
    .io_s(FullAdder_625_io_s),
    .io_co(FullAdder_625_io_co)
  );
  FullAdder FullAdder_626 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_626_io_a),
    .io_b(FullAdder_626_io_b),
    .io_ci(FullAdder_626_io_ci),
    .io_s(FullAdder_626_io_s),
    .io_co(FullAdder_626_io_co)
  );
  FullAdder FullAdder_627 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_627_io_a),
    .io_b(FullAdder_627_io_b),
    .io_ci(FullAdder_627_io_ci),
    .io_s(FullAdder_627_io_s),
    .io_co(FullAdder_627_io_co)
  );
  FullAdder FullAdder_628 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_628_io_a),
    .io_b(FullAdder_628_io_b),
    .io_ci(FullAdder_628_io_ci),
    .io_s(FullAdder_628_io_s),
    .io_co(FullAdder_628_io_co)
  );
  FullAdder FullAdder_629 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_629_io_a),
    .io_b(FullAdder_629_io_b),
    .io_ci(FullAdder_629_io_ci),
    .io_s(FullAdder_629_io_s),
    .io_co(FullAdder_629_io_co)
  );
  FullAdder FullAdder_630 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_630_io_a),
    .io_b(FullAdder_630_io_b),
    .io_ci(FullAdder_630_io_ci),
    .io_s(FullAdder_630_io_s),
    .io_co(FullAdder_630_io_co)
  );
  FullAdder FullAdder_631 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_631_io_a),
    .io_b(FullAdder_631_io_b),
    .io_ci(FullAdder_631_io_ci),
    .io_s(FullAdder_631_io_s),
    .io_co(FullAdder_631_io_co)
  );
  FullAdder FullAdder_632 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_632_io_a),
    .io_b(FullAdder_632_io_b),
    .io_ci(FullAdder_632_io_ci),
    .io_s(FullAdder_632_io_s),
    .io_co(FullAdder_632_io_co)
  );
  HalfAdder HalfAdder_46 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_46_io_a),
    .io_b(HalfAdder_46_io_b),
    .io_s(HalfAdder_46_io_s),
    .io_co(HalfAdder_46_io_co)
  );
  FullAdder FullAdder_633 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_633_io_a),
    .io_b(FullAdder_633_io_b),
    .io_ci(FullAdder_633_io_ci),
    .io_s(FullAdder_633_io_s),
    .io_co(FullAdder_633_io_co)
  );
  FullAdder FullAdder_634 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_634_io_a),
    .io_b(FullAdder_634_io_b),
    .io_ci(FullAdder_634_io_ci),
    .io_s(FullAdder_634_io_s),
    .io_co(FullAdder_634_io_co)
  );
  FullAdder FullAdder_635 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_635_io_a),
    .io_b(FullAdder_635_io_b),
    .io_ci(FullAdder_635_io_ci),
    .io_s(FullAdder_635_io_s),
    .io_co(FullAdder_635_io_co)
  );
  FullAdder FullAdder_636 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_636_io_a),
    .io_b(FullAdder_636_io_b),
    .io_ci(FullAdder_636_io_ci),
    .io_s(FullAdder_636_io_s),
    .io_co(FullAdder_636_io_co)
  );
  FullAdder FullAdder_637 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_637_io_a),
    .io_b(FullAdder_637_io_b),
    .io_ci(FullAdder_637_io_ci),
    .io_s(FullAdder_637_io_s),
    .io_co(FullAdder_637_io_co)
  );
  FullAdder FullAdder_638 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_638_io_a),
    .io_b(FullAdder_638_io_b),
    .io_ci(FullAdder_638_io_ci),
    .io_s(FullAdder_638_io_s),
    .io_co(FullAdder_638_io_co)
  );
  FullAdder FullAdder_639 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_639_io_a),
    .io_b(FullAdder_639_io_b),
    .io_ci(FullAdder_639_io_ci),
    .io_s(FullAdder_639_io_s),
    .io_co(FullAdder_639_io_co)
  );
  FullAdder FullAdder_640 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_640_io_a),
    .io_b(FullAdder_640_io_b),
    .io_ci(FullAdder_640_io_ci),
    .io_s(FullAdder_640_io_s),
    .io_co(FullAdder_640_io_co)
  );
  FullAdder FullAdder_641 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_641_io_a),
    .io_b(FullAdder_641_io_b),
    .io_ci(FullAdder_641_io_ci),
    .io_s(FullAdder_641_io_s),
    .io_co(FullAdder_641_io_co)
  );
  FullAdder FullAdder_642 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_642_io_a),
    .io_b(FullAdder_642_io_b),
    .io_ci(FullAdder_642_io_ci),
    .io_s(FullAdder_642_io_s),
    .io_co(FullAdder_642_io_co)
  );
  FullAdder FullAdder_643 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_643_io_a),
    .io_b(FullAdder_643_io_b),
    .io_ci(FullAdder_643_io_ci),
    .io_s(FullAdder_643_io_s),
    .io_co(FullAdder_643_io_co)
  );
  FullAdder FullAdder_644 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_644_io_a),
    .io_b(FullAdder_644_io_b),
    .io_ci(FullAdder_644_io_ci),
    .io_s(FullAdder_644_io_s),
    .io_co(FullAdder_644_io_co)
  );
  FullAdder FullAdder_645 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_645_io_a),
    .io_b(FullAdder_645_io_b),
    .io_ci(FullAdder_645_io_ci),
    .io_s(FullAdder_645_io_s),
    .io_co(FullAdder_645_io_co)
  );
  FullAdder FullAdder_646 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_646_io_a),
    .io_b(FullAdder_646_io_b),
    .io_ci(FullAdder_646_io_ci),
    .io_s(FullAdder_646_io_s),
    .io_co(FullAdder_646_io_co)
  );
  FullAdder FullAdder_647 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_647_io_a),
    .io_b(FullAdder_647_io_b),
    .io_ci(FullAdder_647_io_ci),
    .io_s(FullAdder_647_io_s),
    .io_co(FullAdder_647_io_co)
  );
  FullAdder FullAdder_648 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_648_io_a),
    .io_b(FullAdder_648_io_b),
    .io_ci(FullAdder_648_io_ci),
    .io_s(FullAdder_648_io_s),
    .io_co(FullAdder_648_io_co)
  );
  FullAdder FullAdder_649 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_649_io_a),
    .io_b(FullAdder_649_io_b),
    .io_ci(FullAdder_649_io_ci),
    .io_s(FullAdder_649_io_s),
    .io_co(FullAdder_649_io_co)
  );
  FullAdder FullAdder_650 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_650_io_a),
    .io_b(FullAdder_650_io_b),
    .io_ci(FullAdder_650_io_ci),
    .io_s(FullAdder_650_io_s),
    .io_co(FullAdder_650_io_co)
  );
  FullAdder FullAdder_651 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_651_io_a),
    .io_b(FullAdder_651_io_b),
    .io_ci(FullAdder_651_io_ci),
    .io_s(FullAdder_651_io_s),
    .io_co(FullAdder_651_io_co)
  );
  FullAdder FullAdder_652 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_652_io_a),
    .io_b(FullAdder_652_io_b),
    .io_ci(FullAdder_652_io_ci),
    .io_s(FullAdder_652_io_s),
    .io_co(FullAdder_652_io_co)
  );
  HalfAdder HalfAdder_47 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_47_io_a),
    .io_b(HalfAdder_47_io_b),
    .io_s(HalfAdder_47_io_s),
    .io_co(HalfAdder_47_io_co)
  );
  FullAdder FullAdder_653 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_653_io_a),
    .io_b(FullAdder_653_io_b),
    .io_ci(FullAdder_653_io_ci),
    .io_s(FullAdder_653_io_s),
    .io_co(FullAdder_653_io_co)
  );
  FullAdder FullAdder_654 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_654_io_a),
    .io_b(FullAdder_654_io_b),
    .io_ci(FullAdder_654_io_ci),
    .io_s(FullAdder_654_io_s),
    .io_co(FullAdder_654_io_co)
  );
  FullAdder FullAdder_655 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_655_io_a),
    .io_b(FullAdder_655_io_b),
    .io_ci(FullAdder_655_io_ci),
    .io_s(FullAdder_655_io_s),
    .io_co(FullAdder_655_io_co)
  );
  FullAdder FullAdder_656 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_656_io_a),
    .io_b(FullAdder_656_io_b),
    .io_ci(FullAdder_656_io_ci),
    .io_s(FullAdder_656_io_s),
    .io_co(FullAdder_656_io_co)
  );
  FullAdder FullAdder_657 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_657_io_a),
    .io_b(FullAdder_657_io_b),
    .io_ci(FullAdder_657_io_ci),
    .io_s(FullAdder_657_io_s),
    .io_co(FullAdder_657_io_co)
  );
  FullAdder FullAdder_658 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_658_io_a),
    .io_b(FullAdder_658_io_b),
    .io_ci(FullAdder_658_io_ci),
    .io_s(FullAdder_658_io_s),
    .io_co(FullAdder_658_io_co)
  );
  FullAdder FullAdder_659 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_659_io_a),
    .io_b(FullAdder_659_io_b),
    .io_ci(FullAdder_659_io_ci),
    .io_s(FullAdder_659_io_s),
    .io_co(FullAdder_659_io_co)
  );
  FullAdder FullAdder_660 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_660_io_a),
    .io_b(FullAdder_660_io_b),
    .io_ci(FullAdder_660_io_ci),
    .io_s(FullAdder_660_io_s),
    .io_co(FullAdder_660_io_co)
  );
  FullAdder FullAdder_661 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_661_io_a),
    .io_b(FullAdder_661_io_b),
    .io_ci(FullAdder_661_io_ci),
    .io_s(FullAdder_661_io_s),
    .io_co(FullAdder_661_io_co)
  );
  FullAdder FullAdder_662 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_662_io_a),
    .io_b(FullAdder_662_io_b),
    .io_ci(FullAdder_662_io_ci),
    .io_s(FullAdder_662_io_s),
    .io_co(FullAdder_662_io_co)
  );
  FullAdder FullAdder_663 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_663_io_a),
    .io_b(FullAdder_663_io_b),
    .io_ci(FullAdder_663_io_ci),
    .io_s(FullAdder_663_io_s),
    .io_co(FullAdder_663_io_co)
  );
  HalfAdder HalfAdder_48 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_48_io_a),
    .io_b(HalfAdder_48_io_b),
    .io_s(HalfAdder_48_io_s),
    .io_co(HalfAdder_48_io_co)
  );
  FullAdder FullAdder_664 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_664_io_a),
    .io_b(FullAdder_664_io_b),
    .io_ci(FullAdder_664_io_ci),
    .io_s(FullAdder_664_io_s),
    .io_co(FullAdder_664_io_co)
  );
  HalfAdder HalfAdder_49 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_49_io_a),
    .io_b(HalfAdder_49_io_b),
    .io_s(HalfAdder_49_io_s),
    .io_co(HalfAdder_49_io_co)
  );
  FullAdder FullAdder_665 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_665_io_a),
    .io_b(FullAdder_665_io_b),
    .io_ci(FullAdder_665_io_ci),
    .io_s(FullAdder_665_io_s),
    .io_co(FullAdder_665_io_co)
  );
  HalfAdder HalfAdder_50 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_50_io_a),
    .io_b(HalfAdder_50_io_b),
    .io_s(HalfAdder_50_io_s),
    .io_co(HalfAdder_50_io_co)
  );
  FullAdder FullAdder_666 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_666_io_a),
    .io_b(FullAdder_666_io_b),
    .io_ci(FullAdder_666_io_ci),
    .io_s(FullAdder_666_io_s),
    .io_co(FullAdder_666_io_co)
  );
  FullAdder FullAdder_667 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_667_io_a),
    .io_b(FullAdder_667_io_b),
    .io_ci(FullAdder_667_io_ci),
    .io_s(FullAdder_667_io_s),
    .io_co(FullAdder_667_io_co)
  );
  FullAdder FullAdder_668 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_668_io_a),
    .io_b(FullAdder_668_io_b),
    .io_ci(FullAdder_668_io_ci),
    .io_s(FullAdder_668_io_s),
    .io_co(FullAdder_668_io_co)
  );
  HalfAdder HalfAdder_51 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_51_io_a),
    .io_b(HalfAdder_51_io_b),
    .io_s(HalfAdder_51_io_s),
    .io_co(HalfAdder_51_io_co)
  );
  HalfAdder HalfAdder_52 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_52_io_a),
    .io_b(HalfAdder_52_io_b),
    .io_s(HalfAdder_52_io_s),
    .io_co(HalfAdder_52_io_co)
  );
  HalfAdder HalfAdder_53 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_53_io_a),
    .io_b(HalfAdder_53_io_b),
    .io_s(HalfAdder_53_io_s),
    .io_co(HalfAdder_53_io_co)
  );
  HalfAdder HalfAdder_54 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_54_io_a),
    .io_b(HalfAdder_54_io_b),
    .io_s(HalfAdder_54_io_s),
    .io_co(HalfAdder_54_io_co)
  );
  HalfAdder HalfAdder_55 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_55_io_a),
    .io_b(HalfAdder_55_io_b),
    .io_s(HalfAdder_55_io_s),
    .io_co(HalfAdder_55_io_co)
  );
  HalfAdder HalfAdder_56 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_56_io_a),
    .io_b(HalfAdder_56_io_b),
    .io_s(HalfAdder_56_io_s),
    .io_co(HalfAdder_56_io_co)
  );
  FullAdder FullAdder_669 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_669_io_a),
    .io_b(FullAdder_669_io_b),
    .io_ci(FullAdder_669_io_ci),
    .io_s(FullAdder_669_io_s),
    .io_co(FullAdder_669_io_co)
  );
  FullAdder FullAdder_670 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_670_io_a),
    .io_b(FullAdder_670_io_b),
    .io_ci(FullAdder_670_io_ci),
    .io_s(FullAdder_670_io_s),
    .io_co(FullAdder_670_io_co)
  );
  FullAdder FullAdder_671 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_671_io_a),
    .io_b(FullAdder_671_io_b),
    .io_ci(FullAdder_671_io_ci),
    .io_s(FullAdder_671_io_s),
    .io_co(FullAdder_671_io_co)
  );
  FullAdder FullAdder_672 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_672_io_a),
    .io_b(FullAdder_672_io_b),
    .io_ci(FullAdder_672_io_ci),
    .io_s(FullAdder_672_io_s),
    .io_co(FullAdder_672_io_co)
  );
  FullAdder FullAdder_673 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_673_io_a),
    .io_b(FullAdder_673_io_b),
    .io_ci(FullAdder_673_io_ci),
    .io_s(FullAdder_673_io_s),
    .io_co(FullAdder_673_io_co)
  );
  FullAdder FullAdder_674 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_674_io_a),
    .io_b(FullAdder_674_io_b),
    .io_ci(FullAdder_674_io_ci),
    .io_s(FullAdder_674_io_s),
    .io_co(FullAdder_674_io_co)
  );
  FullAdder FullAdder_675 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_675_io_a),
    .io_b(FullAdder_675_io_b),
    .io_ci(FullAdder_675_io_ci),
    .io_s(FullAdder_675_io_s),
    .io_co(FullAdder_675_io_co)
  );
  FullAdder FullAdder_676 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_676_io_a),
    .io_b(FullAdder_676_io_b),
    .io_ci(FullAdder_676_io_ci),
    .io_s(FullAdder_676_io_s),
    .io_co(FullAdder_676_io_co)
  );
  HalfAdder HalfAdder_57 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_57_io_a),
    .io_b(HalfAdder_57_io_b),
    .io_s(HalfAdder_57_io_s),
    .io_co(HalfAdder_57_io_co)
  );
  HalfAdder HalfAdder_58 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_58_io_a),
    .io_b(HalfAdder_58_io_b),
    .io_s(HalfAdder_58_io_s),
    .io_co(HalfAdder_58_io_co)
  );
  HalfAdder HalfAdder_59 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_59_io_a),
    .io_b(HalfAdder_59_io_b),
    .io_s(HalfAdder_59_io_s),
    .io_co(HalfAdder_59_io_co)
  );
  HalfAdder HalfAdder_60 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_60_io_a),
    .io_b(HalfAdder_60_io_b),
    .io_s(HalfAdder_60_io_s),
    .io_co(HalfAdder_60_io_co)
  );
  FullAdder FullAdder_677 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_677_io_a),
    .io_b(FullAdder_677_io_b),
    .io_ci(FullAdder_677_io_ci),
    .io_s(FullAdder_677_io_s),
    .io_co(FullAdder_677_io_co)
  );
  FullAdder FullAdder_678 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_678_io_a),
    .io_b(FullAdder_678_io_b),
    .io_ci(FullAdder_678_io_ci),
    .io_s(FullAdder_678_io_s),
    .io_co(FullAdder_678_io_co)
  );
  FullAdder FullAdder_679 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_679_io_a),
    .io_b(FullAdder_679_io_b),
    .io_ci(FullAdder_679_io_ci),
    .io_s(FullAdder_679_io_s),
    .io_co(FullAdder_679_io_co)
  );
  FullAdder FullAdder_680 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_680_io_a),
    .io_b(FullAdder_680_io_b),
    .io_ci(FullAdder_680_io_ci),
    .io_s(FullAdder_680_io_s),
    .io_co(FullAdder_680_io_co)
  );
  FullAdder FullAdder_681 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_681_io_a),
    .io_b(FullAdder_681_io_b),
    .io_ci(FullAdder_681_io_ci),
    .io_s(FullAdder_681_io_s),
    .io_co(FullAdder_681_io_co)
  );
  FullAdder FullAdder_682 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_682_io_a),
    .io_b(FullAdder_682_io_b),
    .io_ci(FullAdder_682_io_ci),
    .io_s(FullAdder_682_io_s),
    .io_co(FullAdder_682_io_co)
  );
  FullAdder FullAdder_683 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_683_io_a),
    .io_b(FullAdder_683_io_b),
    .io_ci(FullAdder_683_io_ci),
    .io_s(FullAdder_683_io_s),
    .io_co(FullAdder_683_io_co)
  );
  FullAdder FullAdder_684 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_684_io_a),
    .io_b(FullAdder_684_io_b),
    .io_ci(FullAdder_684_io_ci),
    .io_s(FullAdder_684_io_s),
    .io_co(FullAdder_684_io_co)
  );
  FullAdder FullAdder_685 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_685_io_a),
    .io_b(FullAdder_685_io_b),
    .io_ci(FullAdder_685_io_ci),
    .io_s(FullAdder_685_io_s),
    .io_co(FullAdder_685_io_co)
  );
  FullAdder FullAdder_686 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_686_io_a),
    .io_b(FullAdder_686_io_b),
    .io_ci(FullAdder_686_io_ci),
    .io_s(FullAdder_686_io_s),
    .io_co(FullAdder_686_io_co)
  );
  FullAdder FullAdder_687 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_687_io_a),
    .io_b(FullAdder_687_io_b),
    .io_ci(FullAdder_687_io_ci),
    .io_s(FullAdder_687_io_s),
    .io_co(FullAdder_687_io_co)
  );
  FullAdder FullAdder_688 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_688_io_a),
    .io_b(FullAdder_688_io_b),
    .io_ci(FullAdder_688_io_ci),
    .io_s(FullAdder_688_io_s),
    .io_co(FullAdder_688_io_co)
  );
  FullAdder FullAdder_689 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_689_io_a),
    .io_b(FullAdder_689_io_b),
    .io_ci(FullAdder_689_io_ci),
    .io_s(FullAdder_689_io_s),
    .io_co(FullAdder_689_io_co)
  );
  FullAdder FullAdder_690 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_690_io_a),
    .io_b(FullAdder_690_io_b),
    .io_ci(FullAdder_690_io_ci),
    .io_s(FullAdder_690_io_s),
    .io_co(FullAdder_690_io_co)
  );
  FullAdder FullAdder_691 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_691_io_a),
    .io_b(FullAdder_691_io_b),
    .io_ci(FullAdder_691_io_ci),
    .io_s(FullAdder_691_io_s),
    .io_co(FullAdder_691_io_co)
  );
  HalfAdder HalfAdder_61 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_61_io_a),
    .io_b(HalfAdder_61_io_b),
    .io_s(HalfAdder_61_io_s),
    .io_co(HalfAdder_61_io_co)
  );
  HalfAdder HalfAdder_62 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_62_io_a),
    .io_b(HalfAdder_62_io_b),
    .io_s(HalfAdder_62_io_s),
    .io_co(HalfAdder_62_io_co)
  );
  FullAdder FullAdder_692 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_692_io_a),
    .io_b(FullAdder_692_io_b),
    .io_ci(FullAdder_692_io_ci),
    .io_s(FullAdder_692_io_s),
    .io_co(FullAdder_692_io_co)
  );
  FullAdder FullAdder_693 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_693_io_a),
    .io_b(FullAdder_693_io_b),
    .io_ci(FullAdder_693_io_ci),
    .io_s(FullAdder_693_io_s),
    .io_co(FullAdder_693_io_co)
  );
  FullAdder FullAdder_694 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_694_io_a),
    .io_b(FullAdder_694_io_b),
    .io_ci(FullAdder_694_io_ci),
    .io_s(FullAdder_694_io_s),
    .io_co(FullAdder_694_io_co)
  );
  FullAdder FullAdder_695 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_695_io_a),
    .io_b(FullAdder_695_io_b),
    .io_ci(FullAdder_695_io_ci),
    .io_s(FullAdder_695_io_s),
    .io_co(FullAdder_695_io_co)
  );
  HalfAdder HalfAdder_63 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_63_io_a),
    .io_b(HalfAdder_63_io_b),
    .io_s(HalfAdder_63_io_s),
    .io_co(HalfAdder_63_io_co)
  );
  FullAdder FullAdder_696 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_696_io_a),
    .io_b(FullAdder_696_io_b),
    .io_ci(FullAdder_696_io_ci),
    .io_s(FullAdder_696_io_s),
    .io_co(FullAdder_696_io_co)
  );
  FullAdder FullAdder_697 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_697_io_a),
    .io_b(FullAdder_697_io_b),
    .io_ci(FullAdder_697_io_ci),
    .io_s(FullAdder_697_io_s),
    .io_co(FullAdder_697_io_co)
  );
  FullAdder FullAdder_698 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_698_io_a),
    .io_b(FullAdder_698_io_b),
    .io_ci(FullAdder_698_io_ci),
    .io_s(FullAdder_698_io_s),
    .io_co(FullAdder_698_io_co)
  );
  FullAdder FullAdder_699 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_699_io_a),
    .io_b(FullAdder_699_io_b),
    .io_ci(FullAdder_699_io_ci),
    .io_s(FullAdder_699_io_s),
    .io_co(FullAdder_699_io_co)
  );
  FullAdder FullAdder_700 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_700_io_a),
    .io_b(FullAdder_700_io_b),
    .io_ci(FullAdder_700_io_ci),
    .io_s(FullAdder_700_io_s),
    .io_co(FullAdder_700_io_co)
  );
  FullAdder FullAdder_701 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_701_io_a),
    .io_b(FullAdder_701_io_b),
    .io_ci(FullAdder_701_io_ci),
    .io_s(FullAdder_701_io_s),
    .io_co(FullAdder_701_io_co)
  );
  FullAdder FullAdder_702 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_702_io_a),
    .io_b(FullAdder_702_io_b),
    .io_ci(FullAdder_702_io_ci),
    .io_s(FullAdder_702_io_s),
    .io_co(FullAdder_702_io_co)
  );
  FullAdder FullAdder_703 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_703_io_a),
    .io_b(FullAdder_703_io_b),
    .io_ci(FullAdder_703_io_ci),
    .io_s(FullAdder_703_io_s),
    .io_co(FullAdder_703_io_co)
  );
  FullAdder FullAdder_704 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_704_io_a),
    .io_b(FullAdder_704_io_b),
    .io_ci(FullAdder_704_io_ci),
    .io_s(FullAdder_704_io_s),
    .io_co(FullAdder_704_io_co)
  );
  FullAdder FullAdder_705 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_705_io_a),
    .io_b(FullAdder_705_io_b),
    .io_ci(FullAdder_705_io_ci),
    .io_s(FullAdder_705_io_s),
    .io_co(FullAdder_705_io_co)
  );
  FullAdder FullAdder_706 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_706_io_a),
    .io_b(FullAdder_706_io_b),
    .io_ci(FullAdder_706_io_ci),
    .io_s(FullAdder_706_io_s),
    .io_co(FullAdder_706_io_co)
  );
  FullAdder FullAdder_707 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_707_io_a),
    .io_b(FullAdder_707_io_b),
    .io_ci(FullAdder_707_io_ci),
    .io_s(FullAdder_707_io_s),
    .io_co(FullAdder_707_io_co)
  );
  FullAdder FullAdder_708 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_708_io_a),
    .io_b(FullAdder_708_io_b),
    .io_ci(FullAdder_708_io_ci),
    .io_s(FullAdder_708_io_s),
    .io_co(FullAdder_708_io_co)
  );
  FullAdder FullAdder_709 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_709_io_a),
    .io_b(FullAdder_709_io_b),
    .io_ci(FullAdder_709_io_ci),
    .io_s(FullAdder_709_io_s),
    .io_co(FullAdder_709_io_co)
  );
  FullAdder FullAdder_710 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_710_io_a),
    .io_b(FullAdder_710_io_b),
    .io_ci(FullAdder_710_io_ci),
    .io_s(FullAdder_710_io_s),
    .io_co(FullAdder_710_io_co)
  );
  FullAdder FullAdder_711 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_711_io_a),
    .io_b(FullAdder_711_io_b),
    .io_ci(FullAdder_711_io_ci),
    .io_s(FullAdder_711_io_s),
    .io_co(FullAdder_711_io_co)
  );
  FullAdder FullAdder_712 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_712_io_a),
    .io_b(FullAdder_712_io_b),
    .io_ci(FullAdder_712_io_ci),
    .io_s(FullAdder_712_io_s),
    .io_co(FullAdder_712_io_co)
  );
  FullAdder FullAdder_713 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_713_io_a),
    .io_b(FullAdder_713_io_b),
    .io_ci(FullAdder_713_io_ci),
    .io_s(FullAdder_713_io_s),
    .io_co(FullAdder_713_io_co)
  );
  FullAdder FullAdder_714 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_714_io_a),
    .io_b(FullAdder_714_io_b),
    .io_ci(FullAdder_714_io_ci),
    .io_s(FullAdder_714_io_s),
    .io_co(FullAdder_714_io_co)
  );
  FullAdder FullAdder_715 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_715_io_a),
    .io_b(FullAdder_715_io_b),
    .io_ci(FullAdder_715_io_ci),
    .io_s(FullAdder_715_io_s),
    .io_co(FullAdder_715_io_co)
  );
  FullAdder FullAdder_716 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_716_io_a),
    .io_b(FullAdder_716_io_b),
    .io_ci(FullAdder_716_io_ci),
    .io_s(FullAdder_716_io_s),
    .io_co(FullAdder_716_io_co)
  );
  FullAdder FullAdder_717 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_717_io_a),
    .io_b(FullAdder_717_io_b),
    .io_ci(FullAdder_717_io_ci),
    .io_s(FullAdder_717_io_s),
    .io_co(FullAdder_717_io_co)
  );
  FullAdder FullAdder_718 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_718_io_a),
    .io_b(FullAdder_718_io_b),
    .io_ci(FullAdder_718_io_ci),
    .io_s(FullAdder_718_io_s),
    .io_co(FullAdder_718_io_co)
  );
  FullAdder FullAdder_719 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_719_io_a),
    .io_b(FullAdder_719_io_b),
    .io_ci(FullAdder_719_io_ci),
    .io_s(FullAdder_719_io_s),
    .io_co(FullAdder_719_io_co)
  );
  FullAdder FullAdder_720 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_720_io_a),
    .io_b(FullAdder_720_io_b),
    .io_ci(FullAdder_720_io_ci),
    .io_s(FullAdder_720_io_s),
    .io_co(FullAdder_720_io_co)
  );
  FullAdder FullAdder_721 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_721_io_a),
    .io_b(FullAdder_721_io_b),
    .io_ci(FullAdder_721_io_ci),
    .io_s(FullAdder_721_io_s),
    .io_co(FullAdder_721_io_co)
  );
  FullAdder FullAdder_722 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_722_io_a),
    .io_b(FullAdder_722_io_b),
    .io_ci(FullAdder_722_io_ci),
    .io_s(FullAdder_722_io_s),
    .io_co(FullAdder_722_io_co)
  );
  FullAdder FullAdder_723 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_723_io_a),
    .io_b(FullAdder_723_io_b),
    .io_ci(FullAdder_723_io_ci),
    .io_s(FullAdder_723_io_s),
    .io_co(FullAdder_723_io_co)
  );
  FullAdder FullAdder_724 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_724_io_a),
    .io_b(FullAdder_724_io_b),
    .io_ci(FullAdder_724_io_ci),
    .io_s(FullAdder_724_io_s),
    .io_co(FullAdder_724_io_co)
  );
  FullAdder FullAdder_725 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_725_io_a),
    .io_b(FullAdder_725_io_b),
    .io_ci(FullAdder_725_io_ci),
    .io_s(FullAdder_725_io_s),
    .io_co(FullAdder_725_io_co)
  );
  FullAdder FullAdder_726 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_726_io_a),
    .io_b(FullAdder_726_io_b),
    .io_ci(FullAdder_726_io_ci),
    .io_s(FullAdder_726_io_s),
    .io_co(FullAdder_726_io_co)
  );
  FullAdder FullAdder_727 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_727_io_a),
    .io_b(FullAdder_727_io_b),
    .io_ci(FullAdder_727_io_ci),
    .io_s(FullAdder_727_io_s),
    .io_co(FullAdder_727_io_co)
  );
  FullAdder FullAdder_728 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_728_io_a),
    .io_b(FullAdder_728_io_b),
    .io_ci(FullAdder_728_io_ci),
    .io_s(FullAdder_728_io_s),
    .io_co(FullAdder_728_io_co)
  );
  FullAdder FullAdder_729 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_729_io_a),
    .io_b(FullAdder_729_io_b),
    .io_ci(FullAdder_729_io_ci),
    .io_s(FullAdder_729_io_s),
    .io_co(FullAdder_729_io_co)
  );
  FullAdder FullAdder_730 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_730_io_a),
    .io_b(FullAdder_730_io_b),
    .io_ci(FullAdder_730_io_ci),
    .io_s(FullAdder_730_io_s),
    .io_co(FullAdder_730_io_co)
  );
  FullAdder FullAdder_731 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_731_io_a),
    .io_b(FullAdder_731_io_b),
    .io_ci(FullAdder_731_io_ci),
    .io_s(FullAdder_731_io_s),
    .io_co(FullAdder_731_io_co)
  );
  FullAdder FullAdder_732 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_732_io_a),
    .io_b(FullAdder_732_io_b),
    .io_ci(FullAdder_732_io_ci),
    .io_s(FullAdder_732_io_s),
    .io_co(FullAdder_732_io_co)
  );
  HalfAdder HalfAdder_64 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_64_io_a),
    .io_b(HalfAdder_64_io_b),
    .io_s(HalfAdder_64_io_s),
    .io_co(HalfAdder_64_io_co)
  );
  FullAdder FullAdder_733 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_733_io_a),
    .io_b(FullAdder_733_io_b),
    .io_ci(FullAdder_733_io_ci),
    .io_s(FullAdder_733_io_s),
    .io_co(FullAdder_733_io_co)
  );
  FullAdder FullAdder_734 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_734_io_a),
    .io_b(FullAdder_734_io_b),
    .io_ci(FullAdder_734_io_ci),
    .io_s(FullAdder_734_io_s),
    .io_co(FullAdder_734_io_co)
  );
  HalfAdder HalfAdder_65 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_65_io_a),
    .io_b(HalfAdder_65_io_b),
    .io_s(HalfAdder_65_io_s),
    .io_co(HalfAdder_65_io_co)
  );
  FullAdder FullAdder_735 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_735_io_a),
    .io_b(FullAdder_735_io_b),
    .io_ci(FullAdder_735_io_ci),
    .io_s(FullAdder_735_io_s),
    .io_co(FullAdder_735_io_co)
  );
  FullAdder FullAdder_736 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_736_io_a),
    .io_b(FullAdder_736_io_b),
    .io_ci(FullAdder_736_io_ci),
    .io_s(FullAdder_736_io_s),
    .io_co(FullAdder_736_io_co)
  );
  FullAdder FullAdder_737 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_737_io_a),
    .io_b(FullAdder_737_io_b),
    .io_ci(FullAdder_737_io_ci),
    .io_s(FullAdder_737_io_s),
    .io_co(FullAdder_737_io_co)
  );
  FullAdder FullAdder_738 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_738_io_a),
    .io_b(FullAdder_738_io_b),
    .io_ci(FullAdder_738_io_ci),
    .io_s(FullAdder_738_io_s),
    .io_co(FullAdder_738_io_co)
  );
  FullAdder FullAdder_739 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_739_io_a),
    .io_b(FullAdder_739_io_b),
    .io_ci(FullAdder_739_io_ci),
    .io_s(FullAdder_739_io_s),
    .io_co(FullAdder_739_io_co)
  );
  FullAdder FullAdder_740 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_740_io_a),
    .io_b(FullAdder_740_io_b),
    .io_ci(FullAdder_740_io_ci),
    .io_s(FullAdder_740_io_s),
    .io_co(FullAdder_740_io_co)
  );
  FullAdder FullAdder_741 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_741_io_a),
    .io_b(FullAdder_741_io_b),
    .io_ci(FullAdder_741_io_ci),
    .io_s(FullAdder_741_io_s),
    .io_co(FullAdder_741_io_co)
  );
  FullAdder FullAdder_742 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_742_io_a),
    .io_b(FullAdder_742_io_b),
    .io_ci(FullAdder_742_io_ci),
    .io_s(FullAdder_742_io_s),
    .io_co(FullAdder_742_io_co)
  );
  FullAdder FullAdder_743 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_743_io_a),
    .io_b(FullAdder_743_io_b),
    .io_ci(FullAdder_743_io_ci),
    .io_s(FullAdder_743_io_s),
    .io_co(FullAdder_743_io_co)
  );
  FullAdder FullAdder_744 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_744_io_a),
    .io_b(FullAdder_744_io_b),
    .io_ci(FullAdder_744_io_ci),
    .io_s(FullAdder_744_io_s),
    .io_co(FullAdder_744_io_co)
  );
  FullAdder FullAdder_745 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_745_io_a),
    .io_b(FullAdder_745_io_b),
    .io_ci(FullAdder_745_io_ci),
    .io_s(FullAdder_745_io_s),
    .io_co(FullAdder_745_io_co)
  );
  FullAdder FullAdder_746 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_746_io_a),
    .io_b(FullAdder_746_io_b),
    .io_ci(FullAdder_746_io_ci),
    .io_s(FullAdder_746_io_s),
    .io_co(FullAdder_746_io_co)
  );
  FullAdder FullAdder_747 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_747_io_a),
    .io_b(FullAdder_747_io_b),
    .io_ci(FullAdder_747_io_ci),
    .io_s(FullAdder_747_io_s),
    .io_co(FullAdder_747_io_co)
  );
  FullAdder FullAdder_748 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_748_io_a),
    .io_b(FullAdder_748_io_b),
    .io_ci(FullAdder_748_io_ci),
    .io_s(FullAdder_748_io_s),
    .io_co(FullAdder_748_io_co)
  );
  FullAdder FullAdder_749 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_749_io_a),
    .io_b(FullAdder_749_io_b),
    .io_ci(FullAdder_749_io_ci),
    .io_s(FullAdder_749_io_s),
    .io_co(FullAdder_749_io_co)
  );
  HalfAdder HalfAdder_66 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_66_io_a),
    .io_b(HalfAdder_66_io_b),
    .io_s(HalfAdder_66_io_s),
    .io_co(HalfAdder_66_io_co)
  );
  FullAdder FullAdder_750 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_750_io_a),
    .io_b(FullAdder_750_io_b),
    .io_ci(FullAdder_750_io_ci),
    .io_s(FullAdder_750_io_s),
    .io_co(FullAdder_750_io_co)
  );
  HalfAdder HalfAdder_67 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_67_io_a),
    .io_b(HalfAdder_67_io_b),
    .io_s(HalfAdder_67_io_s),
    .io_co(HalfAdder_67_io_co)
  );
  FullAdder FullAdder_751 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_751_io_a),
    .io_b(FullAdder_751_io_b),
    .io_ci(FullAdder_751_io_ci),
    .io_s(FullAdder_751_io_s),
    .io_co(FullAdder_751_io_co)
  );
  FullAdder FullAdder_752 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_752_io_a),
    .io_b(FullAdder_752_io_b),
    .io_ci(FullAdder_752_io_ci),
    .io_s(FullAdder_752_io_s),
    .io_co(FullAdder_752_io_co)
  );
  FullAdder FullAdder_753 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_753_io_a),
    .io_b(FullAdder_753_io_b),
    .io_ci(FullAdder_753_io_ci),
    .io_s(FullAdder_753_io_s),
    .io_co(FullAdder_753_io_co)
  );
  FullAdder FullAdder_754 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_754_io_a),
    .io_b(FullAdder_754_io_b),
    .io_ci(FullAdder_754_io_ci),
    .io_s(FullAdder_754_io_s),
    .io_co(FullAdder_754_io_co)
  );
  HalfAdder HalfAdder_68 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_68_io_a),
    .io_b(HalfAdder_68_io_b),
    .io_s(HalfAdder_68_io_s),
    .io_co(HalfAdder_68_io_co)
  );
  HalfAdder HalfAdder_69 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_69_io_a),
    .io_b(HalfAdder_69_io_b),
    .io_s(HalfAdder_69_io_s),
    .io_co(HalfAdder_69_io_co)
  );
  FullAdder FullAdder_755 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_755_io_a),
    .io_b(FullAdder_755_io_b),
    .io_ci(FullAdder_755_io_ci),
    .io_s(FullAdder_755_io_s),
    .io_co(FullAdder_755_io_co)
  );
  FullAdder FullAdder_756 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_756_io_a),
    .io_b(FullAdder_756_io_b),
    .io_ci(FullAdder_756_io_ci),
    .io_s(FullAdder_756_io_s),
    .io_co(FullAdder_756_io_co)
  );
  HalfAdder HalfAdder_70 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_70_io_a),
    .io_b(HalfAdder_70_io_b),
    .io_s(HalfAdder_70_io_s),
    .io_co(HalfAdder_70_io_co)
  );
  FullAdder FullAdder_757 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_757_io_a),
    .io_b(FullAdder_757_io_b),
    .io_ci(FullAdder_757_io_ci),
    .io_s(FullAdder_757_io_s),
    .io_co(FullAdder_757_io_co)
  );
  FullAdder FullAdder_758 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_758_io_a),
    .io_b(FullAdder_758_io_b),
    .io_ci(FullAdder_758_io_ci),
    .io_s(FullAdder_758_io_s),
    .io_co(FullAdder_758_io_co)
  );
  HalfAdder HalfAdder_71 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_71_io_a),
    .io_b(HalfAdder_71_io_b),
    .io_s(HalfAdder_71_io_s),
    .io_co(HalfAdder_71_io_co)
  );
  HalfAdder HalfAdder_72 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_72_io_a),
    .io_b(HalfAdder_72_io_b),
    .io_s(HalfAdder_72_io_s),
    .io_co(HalfAdder_72_io_co)
  );
  HalfAdder HalfAdder_73 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_73_io_a),
    .io_b(HalfAdder_73_io_b),
    .io_s(HalfAdder_73_io_s),
    .io_co(HalfAdder_73_io_co)
  );
  HalfAdder HalfAdder_74 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_74_io_a),
    .io_b(HalfAdder_74_io_b),
    .io_s(HalfAdder_74_io_s),
    .io_co(HalfAdder_74_io_co)
  );
  HalfAdder HalfAdder_75 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_75_io_a),
    .io_b(HalfAdder_75_io_b),
    .io_s(HalfAdder_75_io_s),
    .io_co(HalfAdder_75_io_co)
  );
  FullAdder FullAdder_759 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_759_io_a),
    .io_b(FullAdder_759_io_b),
    .io_ci(FullAdder_759_io_ci),
    .io_s(FullAdder_759_io_s),
    .io_co(FullAdder_759_io_co)
  );
  HalfAdder HalfAdder_76 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_76_io_a),
    .io_b(HalfAdder_76_io_b),
    .io_s(HalfAdder_76_io_s),
    .io_co(HalfAdder_76_io_co)
  );
  HalfAdder HalfAdder_77 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_77_io_a),
    .io_b(HalfAdder_77_io_b),
    .io_s(HalfAdder_77_io_s),
    .io_co(HalfAdder_77_io_co)
  );
  FullAdder FullAdder_760 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_760_io_a),
    .io_b(FullAdder_760_io_b),
    .io_ci(FullAdder_760_io_ci),
    .io_s(FullAdder_760_io_s),
    .io_co(FullAdder_760_io_co)
  );
  FullAdder FullAdder_761 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_761_io_a),
    .io_b(FullAdder_761_io_b),
    .io_ci(FullAdder_761_io_ci),
    .io_s(FullAdder_761_io_s),
    .io_co(FullAdder_761_io_co)
  );
  FullAdder FullAdder_762 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_762_io_a),
    .io_b(FullAdder_762_io_b),
    .io_ci(FullAdder_762_io_ci),
    .io_s(FullAdder_762_io_s),
    .io_co(FullAdder_762_io_co)
  );
  FullAdder FullAdder_763 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_763_io_a),
    .io_b(FullAdder_763_io_b),
    .io_ci(FullAdder_763_io_ci),
    .io_s(FullAdder_763_io_s),
    .io_co(FullAdder_763_io_co)
  );
  FullAdder FullAdder_764 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_764_io_a),
    .io_b(FullAdder_764_io_b),
    .io_ci(FullAdder_764_io_ci),
    .io_s(FullAdder_764_io_s),
    .io_co(FullAdder_764_io_co)
  );
  FullAdder FullAdder_765 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_765_io_a),
    .io_b(FullAdder_765_io_b),
    .io_ci(FullAdder_765_io_ci),
    .io_s(FullAdder_765_io_s),
    .io_co(FullAdder_765_io_co)
  );
  HalfAdder HalfAdder_78 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_78_io_a),
    .io_b(HalfAdder_78_io_b),
    .io_s(HalfAdder_78_io_s),
    .io_co(HalfAdder_78_io_co)
  );
  HalfAdder HalfAdder_79 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_79_io_a),
    .io_b(HalfAdder_79_io_b),
    .io_s(HalfAdder_79_io_s),
    .io_co(HalfAdder_79_io_co)
  );
  HalfAdder HalfAdder_80 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_80_io_a),
    .io_b(HalfAdder_80_io_b),
    .io_s(HalfAdder_80_io_s),
    .io_co(HalfAdder_80_io_co)
  );
  FullAdder FullAdder_766 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_766_io_a),
    .io_b(FullAdder_766_io_b),
    .io_ci(FullAdder_766_io_ci),
    .io_s(FullAdder_766_io_s),
    .io_co(FullAdder_766_io_co)
  );
  FullAdder FullAdder_767 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_767_io_a),
    .io_b(FullAdder_767_io_b),
    .io_ci(FullAdder_767_io_ci),
    .io_s(FullAdder_767_io_s),
    .io_co(FullAdder_767_io_co)
  );
  FullAdder FullAdder_768 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_768_io_a),
    .io_b(FullAdder_768_io_b),
    .io_ci(FullAdder_768_io_ci),
    .io_s(FullAdder_768_io_s),
    .io_co(FullAdder_768_io_co)
  );
  FullAdder FullAdder_769 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_769_io_a),
    .io_b(FullAdder_769_io_b),
    .io_ci(FullAdder_769_io_ci),
    .io_s(FullAdder_769_io_s),
    .io_co(FullAdder_769_io_co)
  );
  FullAdder FullAdder_770 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_770_io_a),
    .io_b(FullAdder_770_io_b),
    .io_ci(FullAdder_770_io_ci),
    .io_s(FullAdder_770_io_s),
    .io_co(FullAdder_770_io_co)
  );
  HalfAdder HalfAdder_81 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_81_io_a),
    .io_b(HalfAdder_81_io_b),
    .io_s(HalfAdder_81_io_s),
    .io_co(HalfAdder_81_io_co)
  );
  FullAdder FullAdder_771 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_771_io_a),
    .io_b(FullAdder_771_io_b),
    .io_ci(FullAdder_771_io_ci),
    .io_s(FullAdder_771_io_s),
    .io_co(FullAdder_771_io_co)
  );
  FullAdder FullAdder_772 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_772_io_a),
    .io_b(FullAdder_772_io_b),
    .io_ci(FullAdder_772_io_ci),
    .io_s(FullAdder_772_io_s),
    .io_co(FullAdder_772_io_co)
  );
  FullAdder FullAdder_773 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_773_io_a),
    .io_b(FullAdder_773_io_b),
    .io_ci(FullAdder_773_io_ci),
    .io_s(FullAdder_773_io_s),
    .io_co(FullAdder_773_io_co)
  );
  HalfAdder HalfAdder_82 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_82_io_a),
    .io_b(HalfAdder_82_io_b),
    .io_s(HalfAdder_82_io_s),
    .io_co(HalfAdder_82_io_co)
  );
  HalfAdder HalfAdder_83 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_83_io_a),
    .io_b(HalfAdder_83_io_b),
    .io_s(HalfAdder_83_io_s),
    .io_co(HalfAdder_83_io_co)
  );
  HalfAdder HalfAdder_84 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_84_io_a),
    .io_b(HalfAdder_84_io_b),
    .io_s(HalfAdder_84_io_s),
    .io_co(HalfAdder_84_io_co)
  );
  FullAdder FullAdder_774 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_774_io_a),
    .io_b(FullAdder_774_io_b),
    .io_ci(FullAdder_774_io_ci),
    .io_s(FullAdder_774_io_s),
    .io_co(FullAdder_774_io_co)
  );
  FullAdder FullAdder_775 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_775_io_a),
    .io_b(FullAdder_775_io_b),
    .io_ci(FullAdder_775_io_ci),
    .io_s(FullAdder_775_io_s),
    .io_co(FullAdder_775_io_co)
  );
  FullAdder FullAdder_776 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_776_io_a),
    .io_b(FullAdder_776_io_b),
    .io_ci(FullAdder_776_io_ci),
    .io_s(FullAdder_776_io_s),
    .io_co(FullAdder_776_io_co)
  );
  HalfAdder HalfAdder_85 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_85_io_a),
    .io_b(HalfAdder_85_io_b),
    .io_s(HalfAdder_85_io_s),
    .io_co(HalfAdder_85_io_co)
  );
  FullAdder FullAdder_777 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_777_io_a),
    .io_b(FullAdder_777_io_b),
    .io_ci(FullAdder_777_io_ci),
    .io_s(FullAdder_777_io_s),
    .io_co(FullAdder_777_io_co)
  );
  FullAdder FullAdder_778 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_778_io_a),
    .io_b(FullAdder_778_io_b),
    .io_ci(FullAdder_778_io_ci),
    .io_s(FullAdder_778_io_s),
    .io_co(FullAdder_778_io_co)
  );
  FullAdder FullAdder_779 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_779_io_a),
    .io_b(FullAdder_779_io_b),
    .io_ci(FullAdder_779_io_ci),
    .io_s(FullAdder_779_io_s),
    .io_co(FullAdder_779_io_co)
  );
  FullAdder FullAdder_780 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_780_io_a),
    .io_b(FullAdder_780_io_b),
    .io_ci(FullAdder_780_io_ci),
    .io_s(FullAdder_780_io_s),
    .io_co(FullAdder_780_io_co)
  );
  FullAdder FullAdder_781 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_781_io_a),
    .io_b(FullAdder_781_io_b),
    .io_ci(FullAdder_781_io_ci),
    .io_s(FullAdder_781_io_s),
    .io_co(FullAdder_781_io_co)
  );
  FullAdder FullAdder_782 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_782_io_a),
    .io_b(FullAdder_782_io_b),
    .io_ci(FullAdder_782_io_ci),
    .io_s(FullAdder_782_io_s),
    .io_co(FullAdder_782_io_co)
  );
  FullAdder FullAdder_783 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_783_io_a),
    .io_b(FullAdder_783_io_b),
    .io_ci(FullAdder_783_io_ci),
    .io_s(FullAdder_783_io_s),
    .io_co(FullAdder_783_io_co)
  );
  FullAdder FullAdder_784 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_784_io_a),
    .io_b(FullAdder_784_io_b),
    .io_ci(FullAdder_784_io_ci),
    .io_s(FullAdder_784_io_s),
    .io_co(FullAdder_784_io_co)
  );
  FullAdder FullAdder_785 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_785_io_a),
    .io_b(FullAdder_785_io_b),
    .io_ci(FullAdder_785_io_ci),
    .io_s(FullAdder_785_io_s),
    .io_co(FullAdder_785_io_co)
  );
  FullAdder FullAdder_786 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_786_io_a),
    .io_b(FullAdder_786_io_b),
    .io_ci(FullAdder_786_io_ci),
    .io_s(FullAdder_786_io_s),
    .io_co(FullAdder_786_io_co)
  );
  FullAdder FullAdder_787 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_787_io_a),
    .io_b(FullAdder_787_io_b),
    .io_ci(FullAdder_787_io_ci),
    .io_s(FullAdder_787_io_s),
    .io_co(FullAdder_787_io_co)
  );
  FullAdder FullAdder_788 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_788_io_a),
    .io_b(FullAdder_788_io_b),
    .io_ci(FullAdder_788_io_ci),
    .io_s(FullAdder_788_io_s),
    .io_co(FullAdder_788_io_co)
  );
  FullAdder FullAdder_789 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_789_io_a),
    .io_b(FullAdder_789_io_b),
    .io_ci(FullAdder_789_io_ci),
    .io_s(FullAdder_789_io_s),
    .io_co(FullAdder_789_io_co)
  );
  FullAdder FullAdder_790 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_790_io_a),
    .io_b(FullAdder_790_io_b),
    .io_ci(FullAdder_790_io_ci),
    .io_s(FullAdder_790_io_s),
    .io_co(FullAdder_790_io_co)
  );
  FullAdder FullAdder_791 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_791_io_a),
    .io_b(FullAdder_791_io_b),
    .io_ci(FullAdder_791_io_ci),
    .io_s(FullAdder_791_io_s),
    .io_co(FullAdder_791_io_co)
  );
  FullAdder FullAdder_792 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_792_io_a),
    .io_b(FullAdder_792_io_b),
    .io_ci(FullAdder_792_io_ci),
    .io_s(FullAdder_792_io_s),
    .io_co(FullAdder_792_io_co)
  );
  FullAdder FullAdder_793 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_793_io_a),
    .io_b(FullAdder_793_io_b),
    .io_ci(FullAdder_793_io_ci),
    .io_s(FullAdder_793_io_s),
    .io_co(FullAdder_793_io_co)
  );
  FullAdder FullAdder_794 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_794_io_a),
    .io_b(FullAdder_794_io_b),
    .io_ci(FullAdder_794_io_ci),
    .io_s(FullAdder_794_io_s),
    .io_co(FullAdder_794_io_co)
  );
  FullAdder FullAdder_795 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_795_io_a),
    .io_b(FullAdder_795_io_b),
    .io_ci(FullAdder_795_io_ci),
    .io_s(FullAdder_795_io_s),
    .io_co(FullAdder_795_io_co)
  );
  FullAdder FullAdder_796 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_796_io_a),
    .io_b(FullAdder_796_io_b),
    .io_ci(FullAdder_796_io_ci),
    .io_s(FullAdder_796_io_s),
    .io_co(FullAdder_796_io_co)
  );
  FullAdder FullAdder_797 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_797_io_a),
    .io_b(FullAdder_797_io_b),
    .io_ci(FullAdder_797_io_ci),
    .io_s(FullAdder_797_io_s),
    .io_co(FullAdder_797_io_co)
  );
  FullAdder FullAdder_798 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_798_io_a),
    .io_b(FullAdder_798_io_b),
    .io_ci(FullAdder_798_io_ci),
    .io_s(FullAdder_798_io_s),
    .io_co(FullAdder_798_io_co)
  );
  FullAdder FullAdder_799 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_799_io_a),
    .io_b(FullAdder_799_io_b),
    .io_ci(FullAdder_799_io_ci),
    .io_s(FullAdder_799_io_s),
    .io_co(FullAdder_799_io_co)
  );
  FullAdder FullAdder_800 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_800_io_a),
    .io_b(FullAdder_800_io_b),
    .io_ci(FullAdder_800_io_ci),
    .io_s(FullAdder_800_io_s),
    .io_co(FullAdder_800_io_co)
  );
  FullAdder FullAdder_801 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_801_io_a),
    .io_b(FullAdder_801_io_b),
    .io_ci(FullAdder_801_io_ci),
    .io_s(FullAdder_801_io_s),
    .io_co(FullAdder_801_io_co)
  );
  FullAdder FullAdder_802 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_802_io_a),
    .io_b(FullAdder_802_io_b),
    .io_ci(FullAdder_802_io_ci),
    .io_s(FullAdder_802_io_s),
    .io_co(FullAdder_802_io_co)
  );
  FullAdder FullAdder_803 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_803_io_a),
    .io_b(FullAdder_803_io_b),
    .io_ci(FullAdder_803_io_ci),
    .io_s(FullAdder_803_io_s),
    .io_co(FullAdder_803_io_co)
  );
  HalfAdder HalfAdder_86 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_86_io_a),
    .io_b(HalfAdder_86_io_b),
    .io_s(HalfAdder_86_io_s),
    .io_co(HalfAdder_86_io_co)
  );
  HalfAdder HalfAdder_87 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_87_io_a),
    .io_b(HalfAdder_87_io_b),
    .io_s(HalfAdder_87_io_s),
    .io_co(HalfAdder_87_io_co)
  );
  HalfAdder HalfAdder_88 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_88_io_a),
    .io_b(HalfAdder_88_io_b),
    .io_s(HalfAdder_88_io_s),
    .io_co(HalfAdder_88_io_co)
  );
  FullAdder FullAdder_804 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_804_io_a),
    .io_b(FullAdder_804_io_b),
    .io_ci(FullAdder_804_io_ci),
    .io_s(FullAdder_804_io_s),
    .io_co(FullAdder_804_io_co)
  );
  HalfAdder HalfAdder_89 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_89_io_a),
    .io_b(HalfAdder_89_io_b),
    .io_s(HalfAdder_89_io_s),
    .io_co(HalfAdder_89_io_co)
  );
  FullAdder FullAdder_805 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_805_io_a),
    .io_b(FullAdder_805_io_b),
    .io_ci(FullAdder_805_io_ci),
    .io_s(FullAdder_805_io_s),
    .io_co(FullAdder_805_io_co)
  );
  FullAdder FullAdder_806 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_806_io_a),
    .io_b(FullAdder_806_io_b),
    .io_ci(FullAdder_806_io_ci),
    .io_s(FullAdder_806_io_s),
    .io_co(FullAdder_806_io_co)
  );
  FullAdder FullAdder_807 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_807_io_a),
    .io_b(FullAdder_807_io_b),
    .io_ci(FullAdder_807_io_ci),
    .io_s(FullAdder_807_io_s),
    .io_co(FullAdder_807_io_co)
  );
  FullAdder FullAdder_808 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_808_io_a),
    .io_b(FullAdder_808_io_b),
    .io_ci(FullAdder_808_io_ci),
    .io_s(FullAdder_808_io_s),
    .io_co(FullAdder_808_io_co)
  );
  FullAdder FullAdder_809 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_809_io_a),
    .io_b(FullAdder_809_io_b),
    .io_ci(FullAdder_809_io_ci),
    .io_s(FullAdder_809_io_s),
    .io_co(FullAdder_809_io_co)
  );
  FullAdder FullAdder_810 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_810_io_a),
    .io_b(FullAdder_810_io_b),
    .io_ci(FullAdder_810_io_ci),
    .io_s(FullAdder_810_io_s),
    .io_co(FullAdder_810_io_co)
  );
  FullAdder FullAdder_811 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_811_io_a),
    .io_b(FullAdder_811_io_b),
    .io_ci(FullAdder_811_io_ci),
    .io_s(FullAdder_811_io_s),
    .io_co(FullAdder_811_io_co)
  );
  HalfAdder HalfAdder_90 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_90_io_a),
    .io_b(HalfAdder_90_io_b),
    .io_s(HalfAdder_90_io_s),
    .io_co(HalfAdder_90_io_co)
  );
  HalfAdder HalfAdder_91 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_91_io_a),
    .io_b(HalfAdder_91_io_b),
    .io_s(HalfAdder_91_io_s),
    .io_co(HalfAdder_91_io_co)
  );
  FullAdder FullAdder_812 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_812_io_a),
    .io_b(FullAdder_812_io_b),
    .io_ci(FullAdder_812_io_ci),
    .io_s(FullAdder_812_io_s),
    .io_co(FullAdder_812_io_co)
  );
  FullAdder FullAdder_813 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_813_io_a),
    .io_b(FullAdder_813_io_b),
    .io_ci(FullAdder_813_io_ci),
    .io_s(FullAdder_813_io_s),
    .io_co(FullAdder_813_io_co)
  );
  FullAdder FullAdder_814 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_814_io_a),
    .io_b(FullAdder_814_io_b),
    .io_ci(FullAdder_814_io_ci),
    .io_s(FullAdder_814_io_s),
    .io_co(FullAdder_814_io_co)
  );
  HalfAdder HalfAdder_92 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_92_io_a),
    .io_b(HalfAdder_92_io_b),
    .io_s(HalfAdder_92_io_s),
    .io_co(HalfAdder_92_io_co)
  );
  FullAdder FullAdder_815 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_815_io_a),
    .io_b(FullAdder_815_io_b),
    .io_ci(FullAdder_815_io_ci),
    .io_s(FullAdder_815_io_s),
    .io_co(FullAdder_815_io_co)
  );
  FullAdder FullAdder_816 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_816_io_a),
    .io_b(FullAdder_816_io_b),
    .io_ci(FullAdder_816_io_ci),
    .io_s(FullAdder_816_io_s),
    .io_co(FullAdder_816_io_co)
  );
  HalfAdder HalfAdder_93 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_93_io_a),
    .io_b(HalfAdder_93_io_b),
    .io_s(HalfAdder_93_io_s),
    .io_co(HalfAdder_93_io_co)
  );
  HalfAdder HalfAdder_94 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_94_io_a),
    .io_b(HalfAdder_94_io_b),
    .io_s(HalfAdder_94_io_s),
    .io_co(HalfAdder_94_io_co)
  );
  HalfAdder HalfAdder_95 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_95_io_a),
    .io_b(HalfAdder_95_io_b),
    .io_s(HalfAdder_95_io_s),
    .io_co(HalfAdder_95_io_co)
  );
  HalfAdder HalfAdder_96 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_96_io_a),
    .io_b(HalfAdder_96_io_b),
    .io_s(HalfAdder_96_io_s),
    .io_co(HalfAdder_96_io_co)
  );
  HalfAdder HalfAdder_97 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_97_io_a),
    .io_b(HalfAdder_97_io_b),
    .io_s(HalfAdder_97_io_s),
    .io_co(HalfAdder_97_io_co)
  );
  HalfAdder HalfAdder_98 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_98_io_a),
    .io_b(HalfAdder_98_io_b),
    .io_s(HalfAdder_98_io_s),
    .io_co(HalfAdder_98_io_co)
  );
  HalfAdder HalfAdder_99 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_99_io_a),
    .io_b(HalfAdder_99_io_b),
    .io_s(HalfAdder_99_io_s),
    .io_co(HalfAdder_99_io_co)
  );
  HalfAdder HalfAdder_100 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_100_io_a),
    .io_b(HalfAdder_100_io_b),
    .io_s(HalfAdder_100_io_s),
    .io_co(HalfAdder_100_io_co)
  );
  HalfAdder HalfAdder_101 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_101_io_a),
    .io_b(HalfAdder_101_io_b),
    .io_s(HalfAdder_101_io_s),
    .io_co(HalfAdder_101_io_co)
  );
  FullAdder FullAdder_817 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_817_io_a),
    .io_b(FullAdder_817_io_b),
    .io_ci(FullAdder_817_io_ci),
    .io_s(FullAdder_817_io_s),
    .io_co(FullAdder_817_io_co)
  );
  HalfAdder HalfAdder_102 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_102_io_a),
    .io_b(HalfAdder_102_io_b),
    .io_s(HalfAdder_102_io_s),
    .io_co(HalfAdder_102_io_co)
  );
  HalfAdder HalfAdder_103 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_103_io_a),
    .io_b(HalfAdder_103_io_b),
    .io_s(HalfAdder_103_io_s),
    .io_co(HalfAdder_103_io_co)
  );
  FullAdder FullAdder_818 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_818_io_a),
    .io_b(FullAdder_818_io_b),
    .io_ci(FullAdder_818_io_ci),
    .io_s(FullAdder_818_io_s),
    .io_co(FullAdder_818_io_co)
  );
  FullAdder FullAdder_819 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_819_io_a),
    .io_b(FullAdder_819_io_b),
    .io_ci(FullAdder_819_io_ci),
    .io_s(FullAdder_819_io_s),
    .io_co(FullAdder_819_io_co)
  );
  HalfAdder HalfAdder_104 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_104_io_a),
    .io_b(HalfAdder_104_io_b),
    .io_s(HalfAdder_104_io_s),
    .io_co(HalfAdder_104_io_co)
  );
  HalfAdder HalfAdder_105 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_105_io_a),
    .io_b(HalfAdder_105_io_b),
    .io_s(HalfAdder_105_io_s),
    .io_co(HalfAdder_105_io_co)
  );
  FullAdder FullAdder_820 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_820_io_a),
    .io_b(FullAdder_820_io_b),
    .io_ci(FullAdder_820_io_ci),
    .io_s(FullAdder_820_io_s),
    .io_co(FullAdder_820_io_co)
  );
  FullAdder FullAdder_821 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_821_io_a),
    .io_b(FullAdder_821_io_b),
    .io_ci(FullAdder_821_io_ci),
    .io_s(FullAdder_821_io_s),
    .io_co(FullAdder_821_io_co)
  );
  FullAdder FullAdder_822 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_822_io_a),
    .io_b(FullAdder_822_io_b),
    .io_ci(FullAdder_822_io_ci),
    .io_s(FullAdder_822_io_s),
    .io_co(FullAdder_822_io_co)
  );
  FullAdder FullAdder_823 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_823_io_a),
    .io_b(FullAdder_823_io_b),
    .io_ci(FullAdder_823_io_ci),
    .io_s(FullAdder_823_io_s),
    .io_co(FullAdder_823_io_co)
  );
  FullAdder FullAdder_824 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_824_io_a),
    .io_b(FullAdder_824_io_b),
    .io_ci(FullAdder_824_io_ci),
    .io_s(FullAdder_824_io_s),
    .io_co(FullAdder_824_io_co)
  );
  FullAdder FullAdder_825 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_825_io_a),
    .io_b(FullAdder_825_io_b),
    .io_ci(FullAdder_825_io_ci),
    .io_s(FullAdder_825_io_s),
    .io_co(FullAdder_825_io_co)
  );
  FullAdder FullAdder_826 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_826_io_a),
    .io_b(FullAdder_826_io_b),
    .io_ci(FullAdder_826_io_ci),
    .io_s(FullAdder_826_io_s),
    .io_co(FullAdder_826_io_co)
  );
  FullAdder FullAdder_827 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_827_io_a),
    .io_b(FullAdder_827_io_b),
    .io_ci(FullAdder_827_io_ci),
    .io_s(FullAdder_827_io_s),
    .io_co(FullAdder_827_io_co)
  );
  HalfAdder HalfAdder_106 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_106_io_a),
    .io_b(HalfAdder_106_io_b),
    .io_s(HalfAdder_106_io_s),
    .io_co(HalfAdder_106_io_co)
  );
  HalfAdder HalfAdder_107 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_107_io_a),
    .io_b(HalfAdder_107_io_b),
    .io_s(HalfAdder_107_io_s),
    .io_co(HalfAdder_107_io_co)
  );
  FullAdder FullAdder_828 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_828_io_a),
    .io_b(FullAdder_828_io_b),
    .io_ci(FullAdder_828_io_ci),
    .io_s(FullAdder_828_io_s),
    .io_co(FullAdder_828_io_co)
  );
  HalfAdder HalfAdder_108 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_108_io_a),
    .io_b(HalfAdder_108_io_b),
    .io_s(HalfAdder_108_io_s),
    .io_co(HalfAdder_108_io_co)
  );
  HalfAdder HalfAdder_109 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_109_io_a),
    .io_b(HalfAdder_109_io_b),
    .io_s(HalfAdder_109_io_s),
    .io_co(HalfAdder_109_io_co)
  );
  FullAdder FullAdder_829 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_829_io_a),
    .io_b(FullAdder_829_io_b),
    .io_ci(FullAdder_829_io_ci),
    .io_s(FullAdder_829_io_s),
    .io_co(FullAdder_829_io_co)
  );
  FullAdder FullAdder_830 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_830_io_a),
    .io_b(FullAdder_830_io_b),
    .io_ci(FullAdder_830_io_ci),
    .io_s(FullAdder_830_io_s),
    .io_co(FullAdder_830_io_co)
  );
  FullAdder FullAdder_831 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_831_io_a),
    .io_b(FullAdder_831_io_b),
    .io_ci(FullAdder_831_io_ci),
    .io_s(FullAdder_831_io_s),
    .io_co(FullAdder_831_io_co)
  );
  HalfAdder HalfAdder_110 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_110_io_a),
    .io_b(HalfAdder_110_io_b),
    .io_s(HalfAdder_110_io_s),
    .io_co(HalfAdder_110_io_co)
  );
  FullAdder FullAdder_832 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_832_io_a),
    .io_b(FullAdder_832_io_b),
    .io_ci(FullAdder_832_io_ci),
    .io_s(FullAdder_832_io_s),
    .io_co(FullAdder_832_io_co)
  );
  FullAdder FullAdder_833 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_833_io_a),
    .io_b(FullAdder_833_io_b),
    .io_ci(FullAdder_833_io_ci),
    .io_s(FullAdder_833_io_s),
    .io_co(FullAdder_833_io_co)
  );
  HalfAdder HalfAdder_111 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_111_io_a),
    .io_b(HalfAdder_111_io_b),
    .io_s(HalfAdder_111_io_s),
    .io_co(HalfAdder_111_io_co)
  );
  FullAdder FullAdder_834 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_834_io_a),
    .io_b(FullAdder_834_io_b),
    .io_ci(FullAdder_834_io_ci),
    .io_s(FullAdder_834_io_s),
    .io_co(FullAdder_834_io_co)
  );
  FullAdder FullAdder_835 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_835_io_a),
    .io_b(FullAdder_835_io_b),
    .io_ci(FullAdder_835_io_ci),
    .io_s(FullAdder_835_io_s),
    .io_co(FullAdder_835_io_co)
  );
  FullAdder FullAdder_836 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_836_io_a),
    .io_b(FullAdder_836_io_b),
    .io_ci(FullAdder_836_io_ci),
    .io_s(FullAdder_836_io_s),
    .io_co(FullAdder_836_io_co)
  );
  FullAdder FullAdder_837 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_837_io_a),
    .io_b(FullAdder_837_io_b),
    .io_ci(FullAdder_837_io_ci),
    .io_s(FullAdder_837_io_s),
    .io_co(FullAdder_837_io_co)
  );
  FullAdder FullAdder_838 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_838_io_a),
    .io_b(FullAdder_838_io_b),
    .io_ci(FullAdder_838_io_ci),
    .io_s(FullAdder_838_io_s),
    .io_co(FullAdder_838_io_co)
  );
  FullAdder FullAdder_839 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_839_io_a),
    .io_b(FullAdder_839_io_b),
    .io_ci(FullAdder_839_io_ci),
    .io_s(FullAdder_839_io_s),
    .io_co(FullAdder_839_io_co)
  );
  FullAdder FullAdder_840 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_840_io_a),
    .io_b(FullAdder_840_io_b),
    .io_ci(FullAdder_840_io_ci),
    .io_s(FullAdder_840_io_s),
    .io_co(FullAdder_840_io_co)
  );
  FullAdder FullAdder_841 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_841_io_a),
    .io_b(FullAdder_841_io_b),
    .io_ci(FullAdder_841_io_ci),
    .io_s(FullAdder_841_io_s),
    .io_co(FullAdder_841_io_co)
  );
  FullAdder FullAdder_842 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_842_io_a),
    .io_b(FullAdder_842_io_b),
    .io_ci(FullAdder_842_io_ci),
    .io_s(FullAdder_842_io_s),
    .io_co(FullAdder_842_io_co)
  );
  HalfAdder HalfAdder_112 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_112_io_a),
    .io_b(HalfAdder_112_io_b),
    .io_s(HalfAdder_112_io_s),
    .io_co(HalfAdder_112_io_co)
  );
  HalfAdder HalfAdder_113 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_113_io_a),
    .io_b(HalfAdder_113_io_b),
    .io_s(HalfAdder_113_io_s),
    .io_co(HalfAdder_113_io_co)
  );
  FullAdder FullAdder_843 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_843_io_a),
    .io_b(FullAdder_843_io_b),
    .io_ci(FullAdder_843_io_ci),
    .io_s(FullAdder_843_io_s),
    .io_co(FullAdder_843_io_co)
  );
  FullAdder FullAdder_844 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_844_io_a),
    .io_b(FullAdder_844_io_b),
    .io_ci(FullAdder_844_io_ci),
    .io_s(FullAdder_844_io_s),
    .io_co(FullAdder_844_io_co)
  );
  FullAdder FullAdder_845 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_845_io_a),
    .io_b(FullAdder_845_io_b),
    .io_ci(FullAdder_845_io_ci),
    .io_s(FullAdder_845_io_s),
    .io_co(FullAdder_845_io_co)
  );
  FullAdder FullAdder_846 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_846_io_a),
    .io_b(FullAdder_846_io_b),
    .io_ci(FullAdder_846_io_ci),
    .io_s(FullAdder_846_io_s),
    .io_co(FullAdder_846_io_co)
  );
  FullAdder FullAdder_847 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_847_io_a),
    .io_b(FullAdder_847_io_b),
    .io_ci(FullAdder_847_io_ci),
    .io_s(FullAdder_847_io_s),
    .io_co(FullAdder_847_io_co)
  );
  FullAdder FullAdder_848 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_848_io_a),
    .io_b(FullAdder_848_io_b),
    .io_ci(FullAdder_848_io_ci),
    .io_s(FullAdder_848_io_s),
    .io_co(FullAdder_848_io_co)
  );
  FullAdder FullAdder_849 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_849_io_a),
    .io_b(FullAdder_849_io_b),
    .io_ci(FullAdder_849_io_ci),
    .io_s(FullAdder_849_io_s),
    .io_co(FullAdder_849_io_co)
  );
  HalfAdder HalfAdder_114 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_114_io_a),
    .io_b(HalfAdder_114_io_b),
    .io_s(HalfAdder_114_io_s),
    .io_co(HalfAdder_114_io_co)
  );
  FullAdder FullAdder_850 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_850_io_a),
    .io_b(FullAdder_850_io_b),
    .io_ci(FullAdder_850_io_ci),
    .io_s(FullAdder_850_io_s),
    .io_co(FullAdder_850_io_co)
  );
  HalfAdder HalfAdder_115 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_115_io_a),
    .io_b(HalfAdder_115_io_b),
    .io_s(HalfAdder_115_io_s),
    .io_co(HalfAdder_115_io_co)
  );
  HalfAdder HalfAdder_116 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_116_io_a),
    .io_b(HalfAdder_116_io_b),
    .io_s(HalfAdder_116_io_s),
    .io_co(HalfAdder_116_io_co)
  );
  HalfAdder HalfAdder_117 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_117_io_a),
    .io_b(HalfAdder_117_io_b),
    .io_s(HalfAdder_117_io_s),
    .io_co(HalfAdder_117_io_co)
  );
  FullAdder FullAdder_851 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_851_io_a),
    .io_b(FullAdder_851_io_b),
    .io_ci(FullAdder_851_io_ci),
    .io_s(FullAdder_851_io_s),
    .io_co(FullAdder_851_io_co)
  );
  HalfAdder HalfAdder_118 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_118_io_a),
    .io_b(HalfAdder_118_io_b),
    .io_s(HalfAdder_118_io_s),
    .io_co(HalfAdder_118_io_co)
  );
  FullAdder FullAdder_852 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_852_io_a),
    .io_b(FullAdder_852_io_b),
    .io_ci(FullAdder_852_io_ci),
    .io_s(FullAdder_852_io_s),
    .io_co(FullAdder_852_io_co)
  );
  HalfAdder HalfAdder_119 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_119_io_a),
    .io_b(HalfAdder_119_io_b),
    .io_s(HalfAdder_119_io_s),
    .io_co(HalfAdder_119_io_co)
  );
  FullAdder FullAdder_853 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_853_io_a),
    .io_b(FullAdder_853_io_b),
    .io_ci(FullAdder_853_io_ci),
    .io_s(FullAdder_853_io_s),
    .io_co(FullAdder_853_io_co)
  );
  HalfAdder HalfAdder_120 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_120_io_a),
    .io_b(HalfAdder_120_io_b),
    .io_s(HalfAdder_120_io_s),
    .io_co(HalfAdder_120_io_co)
  );
  HalfAdder HalfAdder_121 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_121_io_a),
    .io_b(HalfAdder_121_io_b),
    .io_s(HalfAdder_121_io_s),
    .io_co(HalfAdder_121_io_co)
  );
  HalfAdder HalfAdder_122 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_122_io_a),
    .io_b(HalfAdder_122_io_b),
    .io_s(HalfAdder_122_io_s),
    .io_co(HalfAdder_122_io_co)
  );
  FullAdder FullAdder_854 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_854_io_a),
    .io_b(FullAdder_854_io_b),
    .io_ci(FullAdder_854_io_ci),
    .io_s(FullAdder_854_io_s),
    .io_co(FullAdder_854_io_co)
  );
  FullAdder FullAdder_855 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_855_io_a),
    .io_b(FullAdder_855_io_b),
    .io_ci(FullAdder_855_io_ci),
    .io_s(FullAdder_855_io_s),
    .io_co(FullAdder_855_io_co)
  );
  FullAdder FullAdder_856 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_856_io_a),
    .io_b(FullAdder_856_io_b),
    .io_ci(FullAdder_856_io_ci),
    .io_s(FullAdder_856_io_s),
    .io_co(FullAdder_856_io_co)
  );
  HalfAdder HalfAdder_123 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_123_io_a),
    .io_b(HalfAdder_123_io_b),
    .io_s(HalfAdder_123_io_s),
    .io_co(HalfAdder_123_io_co)
  );
  HalfAdder HalfAdder_124 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_124_io_a),
    .io_b(HalfAdder_124_io_b),
    .io_s(HalfAdder_124_io_s),
    .io_co(HalfAdder_124_io_co)
  );
  HalfAdder HalfAdder_125 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_125_io_a),
    .io_b(HalfAdder_125_io_b),
    .io_s(HalfAdder_125_io_s),
    .io_co(HalfAdder_125_io_co)
  );
  HalfAdder HalfAdder_126 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_126_io_a),
    .io_b(HalfAdder_126_io_b),
    .io_s(HalfAdder_126_io_s),
    .io_co(HalfAdder_126_io_co)
  );
  FullAdder FullAdder_857 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_857_io_a),
    .io_b(FullAdder_857_io_b),
    .io_ci(FullAdder_857_io_ci),
    .io_s(FullAdder_857_io_s),
    .io_co(FullAdder_857_io_co)
  );
  FullAdder FullAdder_858 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_858_io_a),
    .io_b(FullAdder_858_io_b),
    .io_ci(FullAdder_858_io_ci),
    .io_s(FullAdder_858_io_s),
    .io_co(FullAdder_858_io_co)
  );
  HalfAdder HalfAdder_127 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_127_io_a),
    .io_b(HalfAdder_127_io_b),
    .io_s(HalfAdder_127_io_s),
    .io_co(HalfAdder_127_io_co)
  );
  HalfAdder HalfAdder_128 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_128_io_a),
    .io_b(HalfAdder_128_io_b),
    .io_s(HalfAdder_128_io_s),
    .io_co(HalfAdder_128_io_co)
  );
  FullAdder FullAdder_859 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_859_io_a),
    .io_b(FullAdder_859_io_b),
    .io_ci(FullAdder_859_io_ci),
    .io_s(FullAdder_859_io_s),
    .io_co(FullAdder_859_io_co)
  );
  HalfAdder HalfAdder_129 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_129_io_a),
    .io_b(HalfAdder_129_io_b),
    .io_s(HalfAdder_129_io_s),
    .io_co(HalfAdder_129_io_co)
  );
  FullAdder FullAdder_860 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_860_io_a),
    .io_b(FullAdder_860_io_b),
    .io_ci(FullAdder_860_io_ci),
    .io_s(FullAdder_860_io_s),
    .io_co(FullAdder_860_io_co)
  );
  FullAdder FullAdder_861 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_861_io_a),
    .io_b(FullAdder_861_io_b),
    .io_ci(FullAdder_861_io_ci),
    .io_s(FullAdder_861_io_s),
    .io_co(FullAdder_861_io_co)
  );
  FullAdder FullAdder_862 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_862_io_a),
    .io_b(FullAdder_862_io_b),
    .io_ci(FullAdder_862_io_ci),
    .io_s(FullAdder_862_io_s),
    .io_co(FullAdder_862_io_co)
  );
  FullAdder FullAdder_863 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_863_io_a),
    .io_b(FullAdder_863_io_b),
    .io_ci(FullAdder_863_io_ci),
    .io_s(FullAdder_863_io_s),
    .io_co(FullAdder_863_io_co)
  );
  FullAdder FullAdder_864 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_864_io_a),
    .io_b(FullAdder_864_io_b),
    .io_ci(FullAdder_864_io_ci),
    .io_s(FullAdder_864_io_s),
    .io_co(FullAdder_864_io_co)
  );
  FullAdder FullAdder_865 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_865_io_a),
    .io_b(FullAdder_865_io_b),
    .io_ci(FullAdder_865_io_ci),
    .io_s(FullAdder_865_io_s),
    .io_co(FullAdder_865_io_co)
  );
  FullAdder FullAdder_866 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_866_io_a),
    .io_b(FullAdder_866_io_b),
    .io_ci(FullAdder_866_io_ci),
    .io_s(FullAdder_866_io_s),
    .io_co(FullAdder_866_io_co)
  );
  FullAdder FullAdder_867 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_867_io_a),
    .io_b(FullAdder_867_io_b),
    .io_ci(FullAdder_867_io_ci),
    .io_s(FullAdder_867_io_s),
    .io_co(FullAdder_867_io_co)
  );
  FullAdder FullAdder_868 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_868_io_a),
    .io_b(FullAdder_868_io_b),
    .io_ci(FullAdder_868_io_ci),
    .io_s(FullAdder_868_io_s),
    .io_co(FullAdder_868_io_co)
  );
  FullAdder FullAdder_869 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_869_io_a),
    .io_b(FullAdder_869_io_b),
    .io_ci(FullAdder_869_io_ci),
    .io_s(FullAdder_869_io_s),
    .io_co(FullAdder_869_io_co)
  );
  FullAdder FullAdder_870 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_870_io_a),
    .io_b(FullAdder_870_io_b),
    .io_ci(FullAdder_870_io_ci),
    .io_s(FullAdder_870_io_s),
    .io_co(FullAdder_870_io_co)
  );
  HalfAdder HalfAdder_130 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_130_io_a),
    .io_b(HalfAdder_130_io_b),
    .io_s(HalfAdder_130_io_s),
    .io_co(HalfAdder_130_io_co)
  );
  FullAdder FullAdder_871 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_871_io_a),
    .io_b(FullAdder_871_io_b),
    .io_ci(FullAdder_871_io_ci),
    .io_s(FullAdder_871_io_s),
    .io_co(FullAdder_871_io_co)
  );
  FullAdder FullAdder_872 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_872_io_a),
    .io_b(FullAdder_872_io_b),
    .io_ci(FullAdder_872_io_ci),
    .io_s(FullAdder_872_io_s),
    .io_co(FullAdder_872_io_co)
  );
  HalfAdder HalfAdder_131 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_131_io_a),
    .io_b(HalfAdder_131_io_b),
    .io_s(HalfAdder_131_io_s),
    .io_co(HalfAdder_131_io_co)
  );
  HalfAdder HalfAdder_132 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_132_io_a),
    .io_b(HalfAdder_132_io_b),
    .io_s(HalfAdder_132_io_s),
    .io_co(HalfAdder_132_io_co)
  );
  FullAdder FullAdder_873 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_873_io_a),
    .io_b(FullAdder_873_io_b),
    .io_ci(FullAdder_873_io_ci),
    .io_s(FullAdder_873_io_s),
    .io_co(FullAdder_873_io_co)
  );
  FullAdder FullAdder_874 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_874_io_a),
    .io_b(FullAdder_874_io_b),
    .io_ci(FullAdder_874_io_ci),
    .io_s(FullAdder_874_io_s),
    .io_co(FullAdder_874_io_co)
  );
  FullAdder FullAdder_875 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_875_io_a),
    .io_b(FullAdder_875_io_b),
    .io_ci(FullAdder_875_io_ci),
    .io_s(FullAdder_875_io_s),
    .io_co(FullAdder_875_io_co)
  );
  HalfAdder HalfAdder_133 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_133_io_a),
    .io_b(HalfAdder_133_io_b),
    .io_s(HalfAdder_133_io_s),
    .io_co(HalfAdder_133_io_co)
  );
  FullAdder FullAdder_876 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_876_io_a),
    .io_b(FullAdder_876_io_b),
    .io_ci(FullAdder_876_io_ci),
    .io_s(FullAdder_876_io_s),
    .io_co(FullAdder_876_io_co)
  );
  FullAdder FullAdder_877 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_877_io_a),
    .io_b(FullAdder_877_io_b),
    .io_ci(FullAdder_877_io_ci),
    .io_s(FullAdder_877_io_s),
    .io_co(FullAdder_877_io_co)
  );
  HalfAdder HalfAdder_134 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_134_io_a),
    .io_b(HalfAdder_134_io_b),
    .io_s(HalfAdder_134_io_s),
    .io_co(HalfAdder_134_io_co)
  );
  FullAdder FullAdder_878 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_878_io_a),
    .io_b(FullAdder_878_io_b),
    .io_ci(FullAdder_878_io_ci),
    .io_s(FullAdder_878_io_s),
    .io_co(FullAdder_878_io_co)
  );
  HalfAdder HalfAdder_135 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_135_io_a),
    .io_b(HalfAdder_135_io_b),
    .io_s(HalfAdder_135_io_s),
    .io_co(HalfAdder_135_io_co)
  );
  HalfAdder HalfAdder_136 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_136_io_a),
    .io_b(HalfAdder_136_io_b),
    .io_s(HalfAdder_136_io_s),
    .io_co(HalfAdder_136_io_co)
  );
  HalfAdder HalfAdder_137 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_137_io_a),
    .io_b(HalfAdder_137_io_b),
    .io_s(HalfAdder_137_io_s),
    .io_co(HalfAdder_137_io_co)
  );
  HalfAdder HalfAdder_138 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_138_io_a),
    .io_b(HalfAdder_138_io_b),
    .io_s(HalfAdder_138_io_s),
    .io_co(HalfAdder_138_io_co)
  );
  HalfAdder HalfAdder_139 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_139_io_a),
    .io_b(HalfAdder_139_io_b),
    .io_s(HalfAdder_139_io_s),
    .io_co(HalfAdder_139_io_co)
  );
  HalfAdder HalfAdder_140 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_140_io_a),
    .io_b(HalfAdder_140_io_b),
    .io_s(HalfAdder_140_io_s),
    .io_co(HalfAdder_140_io_co)
  );
  FullAdder FullAdder_879 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_879_io_a),
    .io_b(FullAdder_879_io_b),
    .io_ci(FullAdder_879_io_ci),
    .io_s(FullAdder_879_io_s),
    .io_co(FullAdder_879_io_co)
  );
  HalfAdder HalfAdder_141 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_141_io_a),
    .io_b(HalfAdder_141_io_b),
    .io_s(HalfAdder_141_io_s),
    .io_co(HalfAdder_141_io_co)
  );
  HalfAdder HalfAdder_142 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_142_io_a),
    .io_b(HalfAdder_142_io_b),
    .io_s(HalfAdder_142_io_s),
    .io_co(HalfAdder_142_io_co)
  );
  FullAdder FullAdder_880 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_880_io_a),
    .io_b(FullAdder_880_io_b),
    .io_ci(FullAdder_880_io_ci),
    .io_s(FullAdder_880_io_s),
    .io_co(FullAdder_880_io_co)
  );
  HalfAdder HalfAdder_143 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_143_io_a),
    .io_b(HalfAdder_143_io_b),
    .io_s(HalfAdder_143_io_s),
    .io_co(HalfAdder_143_io_co)
  );
  FullAdder FullAdder_881 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_881_io_a),
    .io_b(FullAdder_881_io_b),
    .io_ci(FullAdder_881_io_ci),
    .io_s(FullAdder_881_io_s),
    .io_co(FullAdder_881_io_co)
  );
  HalfAdder HalfAdder_144 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_144_io_a),
    .io_b(HalfAdder_144_io_b),
    .io_s(HalfAdder_144_io_s),
    .io_co(HalfAdder_144_io_co)
  );
  HalfAdder HalfAdder_145 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_145_io_a),
    .io_b(HalfAdder_145_io_b),
    .io_s(HalfAdder_145_io_s),
    .io_co(HalfAdder_145_io_co)
  );
  FullAdder FullAdder_882 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_882_io_a),
    .io_b(FullAdder_882_io_b),
    .io_ci(FullAdder_882_io_ci),
    .io_s(FullAdder_882_io_s),
    .io_co(FullAdder_882_io_co)
  );
  FullAdder FullAdder_883 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_883_io_a),
    .io_b(FullAdder_883_io_b),
    .io_ci(FullAdder_883_io_ci),
    .io_s(FullAdder_883_io_s),
    .io_co(FullAdder_883_io_co)
  );
  HalfAdder HalfAdder_146 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_146_io_a),
    .io_b(HalfAdder_146_io_b),
    .io_s(HalfAdder_146_io_s),
    .io_co(HalfAdder_146_io_co)
  );
  FullAdder FullAdder_884 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_884_io_a),
    .io_b(FullAdder_884_io_b),
    .io_ci(FullAdder_884_io_ci),
    .io_s(FullAdder_884_io_s),
    .io_co(FullAdder_884_io_co)
  );
  HalfAdder HalfAdder_147 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_147_io_a),
    .io_b(HalfAdder_147_io_b),
    .io_s(HalfAdder_147_io_s),
    .io_co(HalfAdder_147_io_co)
  );
  FullAdder FullAdder_885 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_885_io_a),
    .io_b(FullAdder_885_io_b),
    .io_ci(FullAdder_885_io_ci),
    .io_s(FullAdder_885_io_s),
    .io_co(FullAdder_885_io_co)
  );
  FullAdder FullAdder_886 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_886_io_a),
    .io_b(FullAdder_886_io_b),
    .io_ci(FullAdder_886_io_ci),
    .io_s(FullAdder_886_io_s),
    .io_co(FullAdder_886_io_co)
  );
  HalfAdder HalfAdder_148 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_148_io_a),
    .io_b(HalfAdder_148_io_b),
    .io_s(HalfAdder_148_io_s),
    .io_co(HalfAdder_148_io_co)
  );
  HalfAdder HalfAdder_149 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_149_io_a),
    .io_b(HalfAdder_149_io_b),
    .io_s(HalfAdder_149_io_s),
    .io_co(HalfAdder_149_io_co)
  );
  FullAdder FullAdder_887 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_887_io_a),
    .io_b(FullAdder_887_io_b),
    .io_ci(FullAdder_887_io_ci),
    .io_s(FullAdder_887_io_s),
    .io_co(FullAdder_887_io_co)
  );
  FullAdder FullAdder_888 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_888_io_a),
    .io_b(FullAdder_888_io_b),
    .io_ci(FullAdder_888_io_ci),
    .io_s(FullAdder_888_io_s),
    .io_co(FullAdder_888_io_co)
  );
  FullAdder FullAdder_889 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_889_io_a),
    .io_b(FullAdder_889_io_b),
    .io_ci(FullAdder_889_io_ci),
    .io_s(FullAdder_889_io_s),
    .io_co(FullAdder_889_io_co)
  );
  HalfAdder HalfAdder_150 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_150_io_a),
    .io_b(HalfAdder_150_io_b),
    .io_s(HalfAdder_150_io_s),
    .io_co(HalfAdder_150_io_co)
  );
  HalfAdder HalfAdder_151 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_151_io_a),
    .io_b(HalfAdder_151_io_b),
    .io_s(HalfAdder_151_io_s),
    .io_co(HalfAdder_151_io_co)
  );
  HalfAdder HalfAdder_152 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_152_io_a),
    .io_b(HalfAdder_152_io_b),
    .io_s(HalfAdder_152_io_s),
    .io_co(HalfAdder_152_io_co)
  );
  FullAdder FullAdder_890 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_890_io_a),
    .io_b(FullAdder_890_io_b),
    .io_ci(FullAdder_890_io_ci),
    .io_s(FullAdder_890_io_s),
    .io_co(FullAdder_890_io_co)
  );
  HalfAdder HalfAdder_153 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_153_io_a),
    .io_b(HalfAdder_153_io_b),
    .io_s(HalfAdder_153_io_s),
    .io_co(HalfAdder_153_io_co)
  );
  FullAdder FullAdder_891 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_891_io_a),
    .io_b(FullAdder_891_io_b),
    .io_ci(FullAdder_891_io_ci),
    .io_s(FullAdder_891_io_s),
    .io_co(FullAdder_891_io_co)
  );
  FullAdder FullAdder_892 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_892_io_a),
    .io_b(FullAdder_892_io_b),
    .io_ci(FullAdder_892_io_ci),
    .io_s(FullAdder_892_io_s),
    .io_co(FullAdder_892_io_co)
  );
  HalfAdder HalfAdder_154 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_154_io_a),
    .io_b(HalfAdder_154_io_b),
    .io_s(HalfAdder_154_io_s),
    .io_co(HalfAdder_154_io_co)
  );
  FullAdder FullAdder_893 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_893_io_a),
    .io_b(FullAdder_893_io_b),
    .io_ci(FullAdder_893_io_ci),
    .io_s(FullAdder_893_io_s),
    .io_co(FullAdder_893_io_co)
  );
  HalfAdder HalfAdder_155 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_155_io_a),
    .io_b(HalfAdder_155_io_b),
    .io_s(HalfAdder_155_io_s),
    .io_co(HalfAdder_155_io_co)
  );
  HalfAdder HalfAdder_156 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_156_io_a),
    .io_b(HalfAdder_156_io_b),
    .io_s(HalfAdder_156_io_s),
    .io_co(HalfAdder_156_io_co)
  );
  HalfAdder HalfAdder_157 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_157_io_a),
    .io_b(HalfAdder_157_io_b),
    .io_s(HalfAdder_157_io_s),
    .io_co(HalfAdder_157_io_co)
  );
  FullAdder FullAdder_894 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_894_io_a),
    .io_b(FullAdder_894_io_b),
    .io_ci(FullAdder_894_io_ci),
    .io_s(FullAdder_894_io_s),
    .io_co(FullAdder_894_io_co)
  );
  HalfAdder HalfAdder_158 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_158_io_a),
    .io_b(HalfAdder_158_io_b),
    .io_s(HalfAdder_158_io_s),
    .io_co(HalfAdder_158_io_co)
  );
  HalfAdder HalfAdder_159 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_159_io_a),
    .io_b(HalfAdder_159_io_b),
    .io_s(HalfAdder_159_io_s),
    .io_co(HalfAdder_159_io_co)
  );
  HalfAdder HalfAdder_160 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_160_io_a),
    .io_b(HalfAdder_160_io_b),
    .io_s(HalfAdder_160_io_s),
    .io_co(HalfAdder_160_io_co)
  );
  FullAdder FullAdder_895 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_895_io_a),
    .io_b(FullAdder_895_io_b),
    .io_ci(FullAdder_895_io_ci),
    .io_s(FullAdder_895_io_s),
    .io_co(FullAdder_895_io_co)
  );
  HalfAdder HalfAdder_161 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_161_io_a),
    .io_b(HalfAdder_161_io_b),
    .io_s(HalfAdder_161_io_s),
    .io_co(HalfAdder_161_io_co)
  );
  HalfAdder HalfAdder_162 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_162_io_a),
    .io_b(HalfAdder_162_io_b),
    .io_s(HalfAdder_162_io_s),
    .io_co(HalfAdder_162_io_co)
  );
  FullAdder FullAdder_896 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_896_io_a),
    .io_b(FullAdder_896_io_b),
    .io_ci(FullAdder_896_io_ci),
    .io_s(FullAdder_896_io_s),
    .io_co(FullAdder_896_io_co)
  );
  HalfAdder HalfAdder_163 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_163_io_a),
    .io_b(HalfAdder_163_io_b),
    .io_s(HalfAdder_163_io_s),
    .io_co(HalfAdder_163_io_co)
  );
  HalfAdder HalfAdder_164 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_164_io_a),
    .io_b(HalfAdder_164_io_b),
    .io_s(HalfAdder_164_io_s),
    .io_co(HalfAdder_164_io_co)
  );
  FullAdder FullAdder_897 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_897_io_a),
    .io_b(FullAdder_897_io_b),
    .io_ci(FullAdder_897_io_ci),
    .io_s(FullAdder_897_io_s),
    .io_co(FullAdder_897_io_co)
  );
  FullAdder FullAdder_898 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_898_io_a),
    .io_b(FullAdder_898_io_b),
    .io_ci(FullAdder_898_io_ci),
    .io_s(FullAdder_898_io_s),
    .io_co(FullAdder_898_io_co)
  );
  HalfAdder HalfAdder_165 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_165_io_a),
    .io_b(HalfAdder_165_io_b),
    .io_s(HalfAdder_165_io_s),
    .io_co(HalfAdder_165_io_co)
  );
  FullAdder FullAdder_899 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_899_io_a),
    .io_b(FullAdder_899_io_b),
    .io_ci(FullAdder_899_io_ci),
    .io_s(FullAdder_899_io_s),
    .io_co(FullAdder_899_io_co)
  );
  HalfAdder HalfAdder_166 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_166_io_a),
    .io_b(HalfAdder_166_io_b),
    .io_s(HalfAdder_166_io_s),
    .io_co(HalfAdder_166_io_co)
  );
  HalfAdder HalfAdder_167 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_167_io_a),
    .io_b(HalfAdder_167_io_b),
    .io_s(HalfAdder_167_io_s),
    .io_co(HalfAdder_167_io_co)
  );
  FullAdder FullAdder_900 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_900_io_a),
    .io_b(FullAdder_900_io_b),
    .io_ci(FullAdder_900_io_ci),
    .io_s(FullAdder_900_io_s),
    .io_co(FullAdder_900_io_co)
  );
  FullAdder FullAdder_901 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_901_io_a),
    .io_b(FullAdder_901_io_b),
    .io_ci(FullAdder_901_io_ci),
    .io_s(FullAdder_901_io_s),
    .io_co(FullAdder_901_io_co)
  );
  HalfAdder HalfAdder_168 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_168_io_a),
    .io_b(HalfAdder_168_io_b),
    .io_s(HalfAdder_168_io_s),
    .io_co(HalfAdder_168_io_co)
  );
  HalfAdder HalfAdder_169 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_169_io_a),
    .io_b(HalfAdder_169_io_b),
    .io_s(HalfAdder_169_io_s),
    .io_co(HalfAdder_169_io_co)
  );
  FullAdder FullAdder_902 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_902_io_a),
    .io_b(FullAdder_902_io_b),
    .io_ci(FullAdder_902_io_ci),
    .io_s(FullAdder_902_io_s),
    .io_co(FullAdder_902_io_co)
  );
  HalfAdder HalfAdder_170 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_170_io_a),
    .io_b(HalfAdder_170_io_b),
    .io_s(HalfAdder_170_io_s),
    .io_co(HalfAdder_170_io_co)
  );
  FullAdder FullAdder_903 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_903_io_a),
    .io_b(FullAdder_903_io_b),
    .io_ci(FullAdder_903_io_ci),
    .io_s(FullAdder_903_io_s),
    .io_co(FullAdder_903_io_co)
  );
  FullAdder FullAdder_904 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_904_io_a),
    .io_b(FullAdder_904_io_b),
    .io_ci(FullAdder_904_io_ci),
    .io_s(FullAdder_904_io_s),
    .io_co(FullAdder_904_io_co)
  );
  FullAdder FullAdder_905 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_905_io_a),
    .io_b(FullAdder_905_io_b),
    .io_ci(FullAdder_905_io_ci),
    .io_s(FullAdder_905_io_s),
    .io_co(FullAdder_905_io_co)
  );
  HalfAdder HalfAdder_171 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_171_io_a),
    .io_b(HalfAdder_171_io_b),
    .io_s(HalfAdder_171_io_s),
    .io_co(HalfAdder_171_io_co)
  );
  FullAdder FullAdder_906 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_906_io_a),
    .io_b(FullAdder_906_io_b),
    .io_ci(FullAdder_906_io_ci),
    .io_s(FullAdder_906_io_s),
    .io_co(FullAdder_906_io_co)
  );
  FullAdder FullAdder_907 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_907_io_a),
    .io_b(FullAdder_907_io_b),
    .io_ci(FullAdder_907_io_ci),
    .io_s(FullAdder_907_io_s),
    .io_co(FullAdder_907_io_co)
  );
  FullAdder FullAdder_908 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_908_io_a),
    .io_b(FullAdder_908_io_b),
    .io_ci(FullAdder_908_io_ci),
    .io_s(FullAdder_908_io_s),
    .io_co(FullAdder_908_io_co)
  );
  HalfAdder HalfAdder_172 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_172_io_a),
    .io_b(HalfAdder_172_io_b),
    .io_s(HalfAdder_172_io_s),
    .io_co(HalfAdder_172_io_co)
  );
  HalfAdder HalfAdder_173 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_173_io_a),
    .io_b(HalfAdder_173_io_b),
    .io_s(HalfAdder_173_io_s),
    .io_co(HalfAdder_173_io_co)
  );
  FullAdder FullAdder_909 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_909_io_a),
    .io_b(FullAdder_909_io_b),
    .io_ci(FullAdder_909_io_ci),
    .io_s(FullAdder_909_io_s),
    .io_co(FullAdder_909_io_co)
  );
  HalfAdder HalfAdder_174 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_174_io_a),
    .io_b(HalfAdder_174_io_b),
    .io_s(HalfAdder_174_io_s),
    .io_co(HalfAdder_174_io_co)
  );
  HalfAdder HalfAdder_175 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_175_io_a),
    .io_b(HalfAdder_175_io_b),
    .io_s(HalfAdder_175_io_s),
    .io_co(HalfAdder_175_io_co)
  );
  HalfAdder HalfAdder_176 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_176_io_a),
    .io_b(HalfAdder_176_io_b),
    .io_s(HalfAdder_176_io_s),
    .io_co(HalfAdder_176_io_co)
  );
  FullAdder FullAdder_910 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_910_io_a),
    .io_b(FullAdder_910_io_b),
    .io_ci(FullAdder_910_io_ci),
    .io_s(FullAdder_910_io_s),
    .io_co(FullAdder_910_io_co)
  );
  HalfAdder HalfAdder_177 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_177_io_a),
    .io_b(HalfAdder_177_io_b),
    .io_s(HalfAdder_177_io_s),
    .io_co(HalfAdder_177_io_co)
  );
  FullAdder FullAdder_911 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_911_io_a),
    .io_b(FullAdder_911_io_b),
    .io_ci(FullAdder_911_io_ci),
    .io_s(FullAdder_911_io_s),
    .io_co(FullAdder_911_io_co)
  );
  FullAdder FullAdder_912 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_912_io_a),
    .io_b(FullAdder_912_io_b),
    .io_ci(FullAdder_912_io_ci),
    .io_s(FullAdder_912_io_s),
    .io_co(FullAdder_912_io_co)
  );
  HalfAdder HalfAdder_178 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_178_io_a),
    .io_b(HalfAdder_178_io_b),
    .io_s(HalfAdder_178_io_s),
    .io_co(HalfAdder_178_io_co)
  );
  FullAdder FullAdder_913 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_913_io_a),
    .io_b(FullAdder_913_io_b),
    .io_ci(FullAdder_913_io_ci),
    .io_s(FullAdder_913_io_s),
    .io_co(FullAdder_913_io_co)
  );
  FullAdder FullAdder_914 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_914_io_a),
    .io_b(FullAdder_914_io_b),
    .io_ci(FullAdder_914_io_ci),
    .io_s(FullAdder_914_io_s),
    .io_co(FullAdder_914_io_co)
  );
  HalfAdder HalfAdder_179 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_179_io_a),
    .io_b(HalfAdder_179_io_b),
    .io_s(HalfAdder_179_io_s),
    .io_co(HalfAdder_179_io_co)
  );
  HalfAdder HalfAdder_180 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_180_io_a),
    .io_b(HalfAdder_180_io_b),
    .io_s(HalfAdder_180_io_s),
    .io_co(HalfAdder_180_io_co)
  );
  FullAdder FullAdder_915 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_915_io_a),
    .io_b(FullAdder_915_io_b),
    .io_ci(FullAdder_915_io_ci),
    .io_s(FullAdder_915_io_s),
    .io_co(FullAdder_915_io_co)
  );
  HalfAdder HalfAdder_181 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_181_io_a),
    .io_b(HalfAdder_181_io_b),
    .io_s(HalfAdder_181_io_s),
    .io_co(HalfAdder_181_io_co)
  );
  HalfAdder HalfAdder_182 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_182_io_a),
    .io_b(HalfAdder_182_io_b),
    .io_s(HalfAdder_182_io_s),
    .io_co(HalfAdder_182_io_co)
  );
  FullAdder FullAdder_916 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_916_io_a),
    .io_b(FullAdder_916_io_b),
    .io_ci(FullAdder_916_io_ci),
    .io_s(FullAdder_916_io_s),
    .io_co(FullAdder_916_io_co)
  );
  HalfAdder HalfAdder_183 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_183_io_a),
    .io_b(HalfAdder_183_io_b),
    .io_s(HalfAdder_183_io_s),
    .io_co(HalfAdder_183_io_co)
  );
  FullAdder FullAdder_917 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_917_io_a),
    .io_b(FullAdder_917_io_b),
    .io_ci(FullAdder_917_io_ci),
    .io_s(FullAdder_917_io_s),
    .io_co(FullAdder_917_io_co)
  );
  FullAdder FullAdder_918 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_918_io_a),
    .io_b(FullAdder_918_io_b),
    .io_ci(FullAdder_918_io_ci),
    .io_s(FullAdder_918_io_s),
    .io_co(FullAdder_918_io_co)
  );
  FullAdder FullAdder_919 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_919_io_a),
    .io_b(FullAdder_919_io_b),
    .io_ci(FullAdder_919_io_ci),
    .io_s(FullAdder_919_io_s),
    .io_co(FullAdder_919_io_co)
  );
  HalfAdder HalfAdder_184 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_184_io_a),
    .io_b(HalfAdder_184_io_b),
    .io_s(HalfAdder_184_io_s),
    .io_co(HalfAdder_184_io_co)
  );
  HalfAdder HalfAdder_185 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_185_io_a),
    .io_b(HalfAdder_185_io_b),
    .io_s(HalfAdder_185_io_s),
    .io_co(HalfAdder_185_io_co)
  );
  FullAdder FullAdder_920 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_920_io_a),
    .io_b(FullAdder_920_io_b),
    .io_ci(FullAdder_920_io_ci),
    .io_s(FullAdder_920_io_s),
    .io_co(FullAdder_920_io_co)
  );
  HalfAdder HalfAdder_186 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_186_io_a),
    .io_b(HalfAdder_186_io_b),
    .io_s(HalfAdder_186_io_s),
    .io_co(HalfAdder_186_io_co)
  );
  FullAdder FullAdder_921 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_921_io_a),
    .io_b(FullAdder_921_io_b),
    .io_ci(FullAdder_921_io_ci),
    .io_s(FullAdder_921_io_s),
    .io_co(FullAdder_921_io_co)
  );
  FullAdder FullAdder_922 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_922_io_a),
    .io_b(FullAdder_922_io_b),
    .io_ci(FullAdder_922_io_ci),
    .io_s(FullAdder_922_io_s),
    .io_co(FullAdder_922_io_co)
  );
  HalfAdder HalfAdder_187 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_187_io_a),
    .io_b(HalfAdder_187_io_b),
    .io_s(HalfAdder_187_io_s),
    .io_co(HalfAdder_187_io_co)
  );
  FullAdder FullAdder_923 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_923_io_a),
    .io_b(FullAdder_923_io_b),
    .io_ci(FullAdder_923_io_ci),
    .io_s(FullAdder_923_io_s),
    .io_co(FullAdder_923_io_co)
  );
  FullAdder FullAdder_924 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_924_io_a),
    .io_b(FullAdder_924_io_b),
    .io_ci(FullAdder_924_io_ci),
    .io_s(FullAdder_924_io_s),
    .io_co(FullAdder_924_io_co)
  );
  FullAdder FullAdder_925 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_925_io_a),
    .io_b(FullAdder_925_io_b),
    .io_ci(FullAdder_925_io_ci),
    .io_s(FullAdder_925_io_s),
    .io_co(FullAdder_925_io_co)
  );
  FullAdder FullAdder_926 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_926_io_a),
    .io_b(FullAdder_926_io_b),
    .io_ci(FullAdder_926_io_ci),
    .io_s(FullAdder_926_io_s),
    .io_co(FullAdder_926_io_co)
  );
  FullAdder FullAdder_927 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_927_io_a),
    .io_b(FullAdder_927_io_b),
    .io_ci(FullAdder_927_io_ci),
    .io_s(FullAdder_927_io_s),
    .io_co(FullAdder_927_io_co)
  );
  FullAdder FullAdder_928 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_928_io_a),
    .io_b(FullAdder_928_io_b),
    .io_ci(FullAdder_928_io_ci),
    .io_s(FullAdder_928_io_s),
    .io_co(FullAdder_928_io_co)
  );
  FullAdder FullAdder_929 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_929_io_a),
    .io_b(FullAdder_929_io_b),
    .io_ci(FullAdder_929_io_ci),
    .io_s(FullAdder_929_io_s),
    .io_co(FullAdder_929_io_co)
  );
  HalfAdder HalfAdder_188 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_188_io_a),
    .io_b(HalfAdder_188_io_b),
    .io_s(HalfAdder_188_io_s),
    .io_co(HalfAdder_188_io_co)
  );
  FullAdder FullAdder_930 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_930_io_a),
    .io_b(FullAdder_930_io_b),
    .io_ci(FullAdder_930_io_ci),
    .io_s(FullAdder_930_io_s),
    .io_co(FullAdder_930_io_co)
  );
  HalfAdder HalfAdder_189 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_189_io_a),
    .io_b(HalfAdder_189_io_b),
    .io_s(HalfAdder_189_io_s),
    .io_co(HalfAdder_189_io_co)
  );
  HalfAdder HalfAdder_190 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_190_io_a),
    .io_b(HalfAdder_190_io_b),
    .io_s(HalfAdder_190_io_s),
    .io_co(HalfAdder_190_io_co)
  );
  assign io_augend = {{1'd0}, _T_1085}; // @[wallace.scala 90:13]
  assign io_addend = {{1'd0}, _T_1147}; // @[wallace.scala 91:13]
  assign HalfAdder_io_a = io_pp_30[31]; // @[wallace.scala 59:18]
  assign HalfAdder_io_b = io_pp_31[30]; // @[wallace.scala 60:18]
  assign HalfAdder_1_io_a = io_pp_29[31]; // @[wallace.scala 59:18]
  assign HalfAdder_1_io_b = io_pp_30[30]; // @[wallace.scala 60:18]
  assign FullAdder_io_a = io_pp_28[31]; // @[wallace.scala 69:18]
  assign FullAdder_io_b = io_pp_29[30]; // @[wallace.scala 70:18]
  assign FullAdder_io_ci = io_pp_30[29]; // @[wallace.scala 71:19]
  assign FullAdder_1_io_a = io_pp_27[31]; // @[wallace.scala 69:18]
  assign FullAdder_1_io_b = io_pp_28[30]; // @[wallace.scala 70:18]
  assign FullAdder_1_io_ci = io_pp_29[29]; // @[wallace.scala 71:19]
  assign HalfAdder_2_io_a = io_pp_30[28]; // @[wallace.scala 59:18]
  assign HalfAdder_2_io_b = io_pp_31[27]; // @[wallace.scala 60:18]
  assign FullAdder_2_io_a = io_pp_26[31]; // @[wallace.scala 69:18]
  assign FullAdder_2_io_b = io_pp_27[30]; // @[wallace.scala 70:18]
  assign FullAdder_2_io_ci = io_pp_28[29]; // @[wallace.scala 71:19]
  assign FullAdder_3_io_a = io_pp_29[28]; // @[wallace.scala 69:18]
  assign FullAdder_3_io_b = io_pp_30[27]; // @[wallace.scala 70:18]
  assign FullAdder_3_io_ci = io_pp_31[26]; // @[wallace.scala 71:19]
  assign FullAdder_4_io_a = io_pp_25[31]; // @[wallace.scala 69:18]
  assign FullAdder_4_io_b = io_pp_26[30]; // @[wallace.scala 70:18]
  assign FullAdder_4_io_ci = io_pp_27[29]; // @[wallace.scala 71:19]
  assign FullAdder_5_io_a = io_pp_28[28]; // @[wallace.scala 69:18]
  assign FullAdder_5_io_b = io_pp_29[27]; // @[wallace.scala 70:18]
  assign FullAdder_5_io_ci = io_pp_30[26]; // @[wallace.scala 71:19]
  assign FullAdder_6_io_a = io_pp_24[31]; // @[wallace.scala 69:18]
  assign FullAdder_6_io_b = io_pp_25[30]; // @[wallace.scala 70:18]
  assign FullAdder_6_io_ci = io_pp_26[29]; // @[wallace.scala 71:19]
  assign FullAdder_7_io_a = io_pp_27[28]; // @[wallace.scala 69:18]
  assign FullAdder_7_io_b = io_pp_28[27]; // @[wallace.scala 70:18]
  assign FullAdder_7_io_ci = io_pp_29[26]; // @[wallace.scala 71:19]
  assign FullAdder_8_io_a = io_pp_23[31]; // @[wallace.scala 69:18]
  assign FullAdder_8_io_b = io_pp_24[30]; // @[wallace.scala 70:18]
  assign FullAdder_8_io_ci = io_pp_25[29]; // @[wallace.scala 71:19]
  assign FullAdder_9_io_a = io_pp_26[28]; // @[wallace.scala 69:18]
  assign FullAdder_9_io_b = io_pp_27[27]; // @[wallace.scala 70:18]
  assign FullAdder_9_io_ci = io_pp_28[26]; // @[wallace.scala 71:19]
  assign FullAdder_10_io_a = io_pp_29[25]; // @[wallace.scala 69:18]
  assign FullAdder_10_io_b = io_pp_30[24]; // @[wallace.scala 70:18]
  assign FullAdder_10_io_ci = io_pp_31[23]; // @[wallace.scala 71:19]
  assign FullAdder_11_io_a = io_pp_22[31]; // @[wallace.scala 69:18]
  assign FullAdder_11_io_b = io_pp_23[30]; // @[wallace.scala 70:18]
  assign FullAdder_11_io_ci = io_pp_24[29]; // @[wallace.scala 71:19]
  assign FullAdder_12_io_a = io_pp_25[28]; // @[wallace.scala 69:18]
  assign FullAdder_12_io_b = io_pp_26[27]; // @[wallace.scala 70:18]
  assign FullAdder_12_io_ci = io_pp_27[26]; // @[wallace.scala 71:19]
  assign FullAdder_13_io_a = io_pp_28[25]; // @[wallace.scala 69:18]
  assign FullAdder_13_io_b = io_pp_29[24]; // @[wallace.scala 70:18]
  assign FullAdder_13_io_ci = io_pp_30[23]; // @[wallace.scala 71:19]
  assign FullAdder_14_io_a = io_pp_21[31]; // @[wallace.scala 69:18]
  assign FullAdder_14_io_b = io_pp_22[30]; // @[wallace.scala 70:18]
  assign FullAdder_14_io_ci = io_pp_23[29]; // @[wallace.scala 71:19]
  assign FullAdder_15_io_a = io_pp_24[28]; // @[wallace.scala 69:18]
  assign FullAdder_15_io_b = io_pp_25[27]; // @[wallace.scala 70:18]
  assign FullAdder_15_io_ci = io_pp_26[26]; // @[wallace.scala 71:19]
  assign FullAdder_16_io_a = io_pp_27[25]; // @[wallace.scala 69:18]
  assign FullAdder_16_io_b = io_pp_28[24]; // @[wallace.scala 70:18]
  assign FullAdder_16_io_ci = io_pp_29[23]; // @[wallace.scala 71:19]
  assign HalfAdder_3_io_a = io_pp_30[22]; // @[wallace.scala 59:18]
  assign HalfAdder_3_io_b = io_pp_31[21]; // @[wallace.scala 60:18]
  assign FullAdder_17_io_a = io_pp_20[31]; // @[wallace.scala 69:18]
  assign FullAdder_17_io_b = io_pp_21[30]; // @[wallace.scala 70:18]
  assign FullAdder_17_io_ci = io_pp_22[29]; // @[wallace.scala 71:19]
  assign FullAdder_18_io_a = io_pp_23[28]; // @[wallace.scala 69:18]
  assign FullAdder_18_io_b = io_pp_24[27]; // @[wallace.scala 70:18]
  assign FullAdder_18_io_ci = io_pp_25[26]; // @[wallace.scala 71:19]
  assign FullAdder_19_io_a = io_pp_26[25]; // @[wallace.scala 69:18]
  assign FullAdder_19_io_b = io_pp_27[24]; // @[wallace.scala 70:18]
  assign FullAdder_19_io_ci = io_pp_28[23]; // @[wallace.scala 71:19]
  assign FullAdder_20_io_a = io_pp_29[22]; // @[wallace.scala 69:18]
  assign FullAdder_20_io_b = io_pp_30[21]; // @[wallace.scala 70:18]
  assign FullAdder_20_io_ci = io_pp_31[20]; // @[wallace.scala 71:19]
  assign FullAdder_21_io_a = io_pp_19[31]; // @[wallace.scala 69:18]
  assign FullAdder_21_io_b = io_pp_20[30]; // @[wallace.scala 70:18]
  assign FullAdder_21_io_ci = io_pp_21[29]; // @[wallace.scala 71:19]
  assign FullAdder_22_io_a = io_pp_22[28]; // @[wallace.scala 69:18]
  assign FullAdder_22_io_b = io_pp_23[27]; // @[wallace.scala 70:18]
  assign FullAdder_22_io_ci = io_pp_24[26]; // @[wallace.scala 71:19]
  assign FullAdder_23_io_a = io_pp_25[25]; // @[wallace.scala 69:18]
  assign FullAdder_23_io_b = io_pp_26[24]; // @[wallace.scala 70:18]
  assign FullAdder_23_io_ci = io_pp_27[23]; // @[wallace.scala 71:19]
  assign FullAdder_24_io_a = io_pp_28[22]; // @[wallace.scala 69:18]
  assign FullAdder_24_io_b = io_pp_29[21]; // @[wallace.scala 70:18]
  assign FullAdder_24_io_ci = io_pp_30[20]; // @[wallace.scala 71:19]
  assign FullAdder_25_io_a = io_pp_18[31]; // @[wallace.scala 69:18]
  assign FullAdder_25_io_b = io_pp_19[30]; // @[wallace.scala 70:18]
  assign FullAdder_25_io_ci = io_pp_20[29]; // @[wallace.scala 71:19]
  assign FullAdder_26_io_a = io_pp_21[28]; // @[wallace.scala 69:18]
  assign FullAdder_26_io_b = io_pp_22[27]; // @[wallace.scala 70:18]
  assign FullAdder_26_io_ci = io_pp_23[26]; // @[wallace.scala 71:19]
  assign FullAdder_27_io_a = io_pp_24[25]; // @[wallace.scala 69:18]
  assign FullAdder_27_io_b = io_pp_25[24]; // @[wallace.scala 70:18]
  assign FullAdder_27_io_ci = io_pp_26[23]; // @[wallace.scala 71:19]
  assign FullAdder_28_io_a = io_pp_27[22]; // @[wallace.scala 69:18]
  assign FullAdder_28_io_b = io_pp_28[21]; // @[wallace.scala 70:18]
  assign FullAdder_28_io_ci = io_pp_29[20]; // @[wallace.scala 71:19]
  assign HalfAdder_4_io_a = io_pp_30[19]; // @[wallace.scala 59:18]
  assign HalfAdder_4_io_b = io_pp_31[18]; // @[wallace.scala 60:18]
  assign FullAdder_29_io_a = io_pp_17[31]; // @[wallace.scala 69:18]
  assign FullAdder_29_io_b = io_pp_18[30]; // @[wallace.scala 70:18]
  assign FullAdder_29_io_ci = io_pp_19[29]; // @[wallace.scala 71:19]
  assign FullAdder_30_io_a = io_pp_20[28]; // @[wallace.scala 69:18]
  assign FullAdder_30_io_b = io_pp_21[27]; // @[wallace.scala 70:18]
  assign FullAdder_30_io_ci = io_pp_22[26]; // @[wallace.scala 71:19]
  assign FullAdder_31_io_a = io_pp_23[25]; // @[wallace.scala 69:18]
  assign FullAdder_31_io_b = io_pp_24[24]; // @[wallace.scala 70:18]
  assign FullAdder_31_io_ci = io_pp_25[23]; // @[wallace.scala 71:19]
  assign FullAdder_32_io_a = io_pp_26[22]; // @[wallace.scala 69:18]
  assign FullAdder_32_io_b = io_pp_27[21]; // @[wallace.scala 70:18]
  assign FullAdder_32_io_ci = io_pp_28[20]; // @[wallace.scala 71:19]
  assign FullAdder_33_io_a = io_pp_29[19]; // @[wallace.scala 69:18]
  assign FullAdder_33_io_b = io_pp_30[18]; // @[wallace.scala 70:18]
  assign FullAdder_33_io_ci = io_pp_31[17]; // @[wallace.scala 71:19]
  assign FullAdder_34_io_a = io_pp_16[31]; // @[wallace.scala 69:18]
  assign FullAdder_34_io_b = io_pp_17[30]; // @[wallace.scala 70:18]
  assign FullAdder_34_io_ci = io_pp_18[29]; // @[wallace.scala 71:19]
  assign FullAdder_35_io_a = io_pp_19[28]; // @[wallace.scala 69:18]
  assign FullAdder_35_io_b = io_pp_20[27]; // @[wallace.scala 70:18]
  assign FullAdder_35_io_ci = io_pp_21[26]; // @[wallace.scala 71:19]
  assign FullAdder_36_io_a = io_pp_22[25]; // @[wallace.scala 69:18]
  assign FullAdder_36_io_b = io_pp_23[24]; // @[wallace.scala 70:18]
  assign FullAdder_36_io_ci = io_pp_24[23]; // @[wallace.scala 71:19]
  assign FullAdder_37_io_a = io_pp_25[22]; // @[wallace.scala 69:18]
  assign FullAdder_37_io_b = io_pp_26[21]; // @[wallace.scala 70:18]
  assign FullAdder_37_io_ci = io_pp_27[20]; // @[wallace.scala 71:19]
  assign FullAdder_38_io_a = io_pp_28[19]; // @[wallace.scala 69:18]
  assign FullAdder_38_io_b = io_pp_29[18]; // @[wallace.scala 70:18]
  assign FullAdder_38_io_ci = io_pp_30[17]; // @[wallace.scala 71:19]
  assign FullAdder_39_io_a = io_pp_15[31]; // @[wallace.scala 69:18]
  assign FullAdder_39_io_b = io_pp_16[30]; // @[wallace.scala 70:18]
  assign FullAdder_39_io_ci = io_pp_17[29]; // @[wallace.scala 71:19]
  assign FullAdder_40_io_a = io_pp_18[28]; // @[wallace.scala 69:18]
  assign FullAdder_40_io_b = io_pp_19[27]; // @[wallace.scala 70:18]
  assign FullAdder_40_io_ci = io_pp_20[26]; // @[wallace.scala 71:19]
  assign FullAdder_41_io_a = io_pp_21[25]; // @[wallace.scala 69:18]
  assign FullAdder_41_io_b = io_pp_22[24]; // @[wallace.scala 70:18]
  assign FullAdder_41_io_ci = io_pp_23[23]; // @[wallace.scala 71:19]
  assign FullAdder_42_io_a = io_pp_24[22]; // @[wallace.scala 69:18]
  assign FullAdder_42_io_b = io_pp_25[21]; // @[wallace.scala 70:18]
  assign FullAdder_42_io_ci = io_pp_26[20]; // @[wallace.scala 71:19]
  assign FullAdder_43_io_a = io_pp_27[19]; // @[wallace.scala 69:18]
  assign FullAdder_43_io_b = io_pp_28[18]; // @[wallace.scala 70:18]
  assign FullAdder_43_io_ci = io_pp_29[17]; // @[wallace.scala 71:19]
  assign HalfAdder_5_io_a = io_pp_30[16]; // @[wallace.scala 59:18]
  assign HalfAdder_5_io_b = io_pp_31[15]; // @[wallace.scala 60:18]
  assign FullAdder_44_io_a = io_pp_14[31]; // @[wallace.scala 69:18]
  assign FullAdder_44_io_b = io_pp_15[30]; // @[wallace.scala 70:18]
  assign FullAdder_44_io_ci = io_pp_16[29]; // @[wallace.scala 71:19]
  assign FullAdder_45_io_a = io_pp_17[28]; // @[wallace.scala 69:18]
  assign FullAdder_45_io_b = io_pp_18[27]; // @[wallace.scala 70:18]
  assign FullAdder_45_io_ci = io_pp_19[26]; // @[wallace.scala 71:19]
  assign FullAdder_46_io_a = io_pp_20[25]; // @[wallace.scala 69:18]
  assign FullAdder_46_io_b = io_pp_21[24]; // @[wallace.scala 70:18]
  assign FullAdder_46_io_ci = io_pp_22[23]; // @[wallace.scala 71:19]
  assign FullAdder_47_io_a = io_pp_23[22]; // @[wallace.scala 69:18]
  assign FullAdder_47_io_b = io_pp_24[21]; // @[wallace.scala 70:18]
  assign FullAdder_47_io_ci = io_pp_25[20]; // @[wallace.scala 71:19]
  assign FullAdder_48_io_a = io_pp_26[19]; // @[wallace.scala 69:18]
  assign FullAdder_48_io_b = io_pp_27[18]; // @[wallace.scala 70:18]
  assign FullAdder_48_io_ci = io_pp_28[17]; // @[wallace.scala 71:19]
  assign FullAdder_49_io_a = io_pp_29[16]; // @[wallace.scala 69:18]
  assign FullAdder_49_io_b = io_pp_30[15]; // @[wallace.scala 70:18]
  assign FullAdder_49_io_ci = io_pp_31[14]; // @[wallace.scala 71:19]
  assign FullAdder_50_io_a = io_pp_13[31]; // @[wallace.scala 69:18]
  assign FullAdder_50_io_b = io_pp_14[30]; // @[wallace.scala 70:18]
  assign FullAdder_50_io_ci = io_pp_15[29]; // @[wallace.scala 71:19]
  assign FullAdder_51_io_a = io_pp_16[28]; // @[wallace.scala 69:18]
  assign FullAdder_51_io_b = io_pp_17[27]; // @[wallace.scala 70:18]
  assign FullAdder_51_io_ci = io_pp_18[26]; // @[wallace.scala 71:19]
  assign FullAdder_52_io_a = io_pp_19[25]; // @[wallace.scala 69:18]
  assign FullAdder_52_io_b = io_pp_20[24]; // @[wallace.scala 70:18]
  assign FullAdder_52_io_ci = io_pp_21[23]; // @[wallace.scala 71:19]
  assign FullAdder_53_io_a = io_pp_22[22]; // @[wallace.scala 69:18]
  assign FullAdder_53_io_b = io_pp_23[21]; // @[wallace.scala 70:18]
  assign FullAdder_53_io_ci = io_pp_24[20]; // @[wallace.scala 71:19]
  assign FullAdder_54_io_a = io_pp_25[19]; // @[wallace.scala 69:18]
  assign FullAdder_54_io_b = io_pp_26[18]; // @[wallace.scala 70:18]
  assign FullAdder_54_io_ci = io_pp_27[17]; // @[wallace.scala 71:19]
  assign FullAdder_55_io_a = io_pp_28[16]; // @[wallace.scala 69:18]
  assign FullAdder_55_io_b = io_pp_29[15]; // @[wallace.scala 70:18]
  assign FullAdder_55_io_ci = io_pp_30[14]; // @[wallace.scala 71:19]
  assign FullAdder_56_io_a = io_pp_12[31]; // @[wallace.scala 69:18]
  assign FullAdder_56_io_b = io_pp_13[30]; // @[wallace.scala 70:18]
  assign FullAdder_56_io_ci = io_pp_14[29]; // @[wallace.scala 71:19]
  assign FullAdder_57_io_a = io_pp_15[28]; // @[wallace.scala 69:18]
  assign FullAdder_57_io_b = io_pp_16[27]; // @[wallace.scala 70:18]
  assign FullAdder_57_io_ci = io_pp_17[26]; // @[wallace.scala 71:19]
  assign FullAdder_58_io_a = io_pp_18[25]; // @[wallace.scala 69:18]
  assign FullAdder_58_io_b = io_pp_19[24]; // @[wallace.scala 70:18]
  assign FullAdder_58_io_ci = io_pp_20[23]; // @[wallace.scala 71:19]
  assign FullAdder_59_io_a = io_pp_21[22]; // @[wallace.scala 69:18]
  assign FullAdder_59_io_b = io_pp_22[21]; // @[wallace.scala 70:18]
  assign FullAdder_59_io_ci = io_pp_23[20]; // @[wallace.scala 71:19]
  assign FullAdder_60_io_a = io_pp_24[19]; // @[wallace.scala 69:18]
  assign FullAdder_60_io_b = io_pp_25[18]; // @[wallace.scala 70:18]
  assign FullAdder_60_io_ci = io_pp_26[17]; // @[wallace.scala 71:19]
  assign FullAdder_61_io_a = io_pp_27[16]; // @[wallace.scala 69:18]
  assign FullAdder_61_io_b = io_pp_28[15]; // @[wallace.scala 70:18]
  assign FullAdder_61_io_ci = io_pp_29[14]; // @[wallace.scala 71:19]
  assign FullAdder_62_io_a = io_pp_11[31]; // @[wallace.scala 69:18]
  assign FullAdder_62_io_b = io_pp_12[30]; // @[wallace.scala 70:18]
  assign FullAdder_62_io_ci = io_pp_13[29]; // @[wallace.scala 71:19]
  assign FullAdder_63_io_a = io_pp_14[28]; // @[wallace.scala 69:18]
  assign FullAdder_63_io_b = io_pp_15[27]; // @[wallace.scala 70:18]
  assign FullAdder_63_io_ci = io_pp_16[26]; // @[wallace.scala 71:19]
  assign FullAdder_64_io_a = io_pp_17[25]; // @[wallace.scala 69:18]
  assign FullAdder_64_io_b = io_pp_18[24]; // @[wallace.scala 70:18]
  assign FullAdder_64_io_ci = io_pp_19[23]; // @[wallace.scala 71:19]
  assign FullAdder_65_io_a = io_pp_20[22]; // @[wallace.scala 69:18]
  assign FullAdder_65_io_b = io_pp_21[21]; // @[wallace.scala 70:18]
  assign FullAdder_65_io_ci = io_pp_22[20]; // @[wallace.scala 71:19]
  assign FullAdder_66_io_a = io_pp_23[19]; // @[wallace.scala 69:18]
  assign FullAdder_66_io_b = io_pp_24[18]; // @[wallace.scala 70:18]
  assign FullAdder_66_io_ci = io_pp_25[17]; // @[wallace.scala 71:19]
  assign FullAdder_67_io_a = io_pp_26[16]; // @[wallace.scala 69:18]
  assign FullAdder_67_io_b = io_pp_27[15]; // @[wallace.scala 70:18]
  assign FullAdder_67_io_ci = io_pp_28[14]; // @[wallace.scala 71:19]
  assign FullAdder_68_io_a = io_pp_29[13]; // @[wallace.scala 69:18]
  assign FullAdder_68_io_b = io_pp_30[12]; // @[wallace.scala 70:18]
  assign FullAdder_68_io_ci = io_pp_31[11]; // @[wallace.scala 71:19]
  assign FullAdder_69_io_a = io_pp_10[31]; // @[wallace.scala 69:18]
  assign FullAdder_69_io_b = io_pp_11[30]; // @[wallace.scala 70:18]
  assign FullAdder_69_io_ci = io_pp_12[29]; // @[wallace.scala 71:19]
  assign FullAdder_70_io_a = io_pp_13[28]; // @[wallace.scala 69:18]
  assign FullAdder_70_io_b = io_pp_14[27]; // @[wallace.scala 70:18]
  assign FullAdder_70_io_ci = io_pp_15[26]; // @[wallace.scala 71:19]
  assign FullAdder_71_io_a = io_pp_16[25]; // @[wallace.scala 69:18]
  assign FullAdder_71_io_b = io_pp_17[24]; // @[wallace.scala 70:18]
  assign FullAdder_71_io_ci = io_pp_18[23]; // @[wallace.scala 71:19]
  assign FullAdder_72_io_a = io_pp_19[22]; // @[wallace.scala 69:18]
  assign FullAdder_72_io_b = io_pp_20[21]; // @[wallace.scala 70:18]
  assign FullAdder_72_io_ci = io_pp_21[20]; // @[wallace.scala 71:19]
  assign FullAdder_73_io_a = io_pp_22[19]; // @[wallace.scala 69:18]
  assign FullAdder_73_io_b = io_pp_23[18]; // @[wallace.scala 70:18]
  assign FullAdder_73_io_ci = io_pp_24[17]; // @[wallace.scala 71:19]
  assign FullAdder_74_io_a = io_pp_25[16]; // @[wallace.scala 69:18]
  assign FullAdder_74_io_b = io_pp_26[15]; // @[wallace.scala 70:18]
  assign FullAdder_74_io_ci = io_pp_27[14]; // @[wallace.scala 71:19]
  assign FullAdder_75_io_a = io_pp_28[13]; // @[wallace.scala 69:18]
  assign FullAdder_75_io_b = io_pp_29[12]; // @[wallace.scala 70:18]
  assign FullAdder_75_io_ci = io_pp_30[11]; // @[wallace.scala 71:19]
  assign FullAdder_76_io_a = io_pp_9[31]; // @[wallace.scala 69:18]
  assign FullAdder_76_io_b = io_pp_10[30]; // @[wallace.scala 70:18]
  assign FullAdder_76_io_ci = io_pp_11[29]; // @[wallace.scala 71:19]
  assign FullAdder_77_io_a = io_pp_12[28]; // @[wallace.scala 69:18]
  assign FullAdder_77_io_b = io_pp_13[27]; // @[wallace.scala 70:18]
  assign FullAdder_77_io_ci = io_pp_14[26]; // @[wallace.scala 71:19]
  assign FullAdder_78_io_a = io_pp_15[25]; // @[wallace.scala 69:18]
  assign FullAdder_78_io_b = io_pp_16[24]; // @[wallace.scala 70:18]
  assign FullAdder_78_io_ci = io_pp_17[23]; // @[wallace.scala 71:19]
  assign FullAdder_79_io_a = io_pp_18[22]; // @[wallace.scala 69:18]
  assign FullAdder_79_io_b = io_pp_19[21]; // @[wallace.scala 70:18]
  assign FullAdder_79_io_ci = io_pp_20[20]; // @[wallace.scala 71:19]
  assign FullAdder_80_io_a = io_pp_21[19]; // @[wallace.scala 69:18]
  assign FullAdder_80_io_b = io_pp_22[18]; // @[wallace.scala 70:18]
  assign FullAdder_80_io_ci = io_pp_23[17]; // @[wallace.scala 71:19]
  assign FullAdder_81_io_a = io_pp_24[16]; // @[wallace.scala 69:18]
  assign FullAdder_81_io_b = io_pp_25[15]; // @[wallace.scala 70:18]
  assign FullAdder_81_io_ci = io_pp_26[14]; // @[wallace.scala 71:19]
  assign FullAdder_82_io_a = io_pp_27[13]; // @[wallace.scala 69:18]
  assign FullAdder_82_io_b = io_pp_28[12]; // @[wallace.scala 70:18]
  assign FullAdder_82_io_ci = io_pp_29[11]; // @[wallace.scala 71:19]
  assign HalfAdder_6_io_a = io_pp_30[10]; // @[wallace.scala 59:18]
  assign HalfAdder_6_io_b = io_pp_31[9]; // @[wallace.scala 60:18]
  assign FullAdder_83_io_a = io_pp_8[31]; // @[wallace.scala 69:18]
  assign FullAdder_83_io_b = io_pp_9[30]; // @[wallace.scala 70:18]
  assign FullAdder_83_io_ci = io_pp_10[29]; // @[wallace.scala 71:19]
  assign FullAdder_84_io_a = io_pp_11[28]; // @[wallace.scala 69:18]
  assign FullAdder_84_io_b = io_pp_12[27]; // @[wallace.scala 70:18]
  assign FullAdder_84_io_ci = io_pp_13[26]; // @[wallace.scala 71:19]
  assign FullAdder_85_io_a = io_pp_14[25]; // @[wallace.scala 69:18]
  assign FullAdder_85_io_b = io_pp_15[24]; // @[wallace.scala 70:18]
  assign FullAdder_85_io_ci = io_pp_16[23]; // @[wallace.scala 71:19]
  assign FullAdder_86_io_a = io_pp_17[22]; // @[wallace.scala 69:18]
  assign FullAdder_86_io_b = io_pp_18[21]; // @[wallace.scala 70:18]
  assign FullAdder_86_io_ci = io_pp_19[20]; // @[wallace.scala 71:19]
  assign FullAdder_87_io_a = io_pp_20[19]; // @[wallace.scala 69:18]
  assign FullAdder_87_io_b = io_pp_21[18]; // @[wallace.scala 70:18]
  assign FullAdder_87_io_ci = io_pp_22[17]; // @[wallace.scala 71:19]
  assign FullAdder_88_io_a = io_pp_23[16]; // @[wallace.scala 69:18]
  assign FullAdder_88_io_b = io_pp_24[15]; // @[wallace.scala 70:18]
  assign FullAdder_88_io_ci = io_pp_25[14]; // @[wallace.scala 71:19]
  assign FullAdder_89_io_a = io_pp_26[13]; // @[wallace.scala 69:18]
  assign FullAdder_89_io_b = io_pp_27[12]; // @[wallace.scala 70:18]
  assign FullAdder_89_io_ci = io_pp_28[11]; // @[wallace.scala 71:19]
  assign FullAdder_90_io_a = io_pp_29[10]; // @[wallace.scala 69:18]
  assign FullAdder_90_io_b = io_pp_30[9]; // @[wallace.scala 70:18]
  assign FullAdder_90_io_ci = io_pp_31[8]; // @[wallace.scala 71:19]
  assign FullAdder_91_io_a = io_pp_7[31]; // @[wallace.scala 69:18]
  assign FullAdder_91_io_b = io_pp_8[30]; // @[wallace.scala 70:18]
  assign FullAdder_91_io_ci = io_pp_9[29]; // @[wallace.scala 71:19]
  assign FullAdder_92_io_a = io_pp_10[28]; // @[wallace.scala 69:18]
  assign FullAdder_92_io_b = io_pp_11[27]; // @[wallace.scala 70:18]
  assign FullAdder_92_io_ci = io_pp_12[26]; // @[wallace.scala 71:19]
  assign FullAdder_93_io_a = io_pp_13[25]; // @[wallace.scala 69:18]
  assign FullAdder_93_io_b = io_pp_14[24]; // @[wallace.scala 70:18]
  assign FullAdder_93_io_ci = io_pp_15[23]; // @[wallace.scala 71:19]
  assign FullAdder_94_io_a = io_pp_16[22]; // @[wallace.scala 69:18]
  assign FullAdder_94_io_b = io_pp_17[21]; // @[wallace.scala 70:18]
  assign FullAdder_94_io_ci = io_pp_18[20]; // @[wallace.scala 71:19]
  assign FullAdder_95_io_a = io_pp_19[19]; // @[wallace.scala 69:18]
  assign FullAdder_95_io_b = io_pp_20[18]; // @[wallace.scala 70:18]
  assign FullAdder_95_io_ci = io_pp_21[17]; // @[wallace.scala 71:19]
  assign FullAdder_96_io_a = io_pp_22[16]; // @[wallace.scala 69:18]
  assign FullAdder_96_io_b = io_pp_23[15]; // @[wallace.scala 70:18]
  assign FullAdder_96_io_ci = io_pp_24[14]; // @[wallace.scala 71:19]
  assign FullAdder_97_io_a = io_pp_25[13]; // @[wallace.scala 69:18]
  assign FullAdder_97_io_b = io_pp_26[12]; // @[wallace.scala 70:18]
  assign FullAdder_97_io_ci = io_pp_27[11]; // @[wallace.scala 71:19]
  assign FullAdder_98_io_a = io_pp_28[10]; // @[wallace.scala 69:18]
  assign FullAdder_98_io_b = io_pp_29[9]; // @[wallace.scala 70:18]
  assign FullAdder_98_io_ci = io_pp_30[8]; // @[wallace.scala 71:19]
  assign FullAdder_99_io_a = io_pp_6[31]; // @[wallace.scala 69:18]
  assign FullAdder_99_io_b = io_pp_7[30]; // @[wallace.scala 70:18]
  assign FullAdder_99_io_ci = io_pp_8[29]; // @[wallace.scala 71:19]
  assign FullAdder_100_io_a = io_pp_9[28]; // @[wallace.scala 69:18]
  assign FullAdder_100_io_b = io_pp_10[27]; // @[wallace.scala 70:18]
  assign FullAdder_100_io_ci = io_pp_11[26]; // @[wallace.scala 71:19]
  assign FullAdder_101_io_a = io_pp_12[25]; // @[wallace.scala 69:18]
  assign FullAdder_101_io_b = io_pp_13[24]; // @[wallace.scala 70:18]
  assign FullAdder_101_io_ci = io_pp_14[23]; // @[wallace.scala 71:19]
  assign FullAdder_102_io_a = io_pp_15[22]; // @[wallace.scala 69:18]
  assign FullAdder_102_io_b = io_pp_16[21]; // @[wallace.scala 70:18]
  assign FullAdder_102_io_ci = io_pp_17[20]; // @[wallace.scala 71:19]
  assign FullAdder_103_io_a = io_pp_18[19]; // @[wallace.scala 69:18]
  assign FullAdder_103_io_b = io_pp_19[18]; // @[wallace.scala 70:18]
  assign FullAdder_103_io_ci = io_pp_20[17]; // @[wallace.scala 71:19]
  assign FullAdder_104_io_a = io_pp_21[16]; // @[wallace.scala 69:18]
  assign FullAdder_104_io_b = io_pp_22[15]; // @[wallace.scala 70:18]
  assign FullAdder_104_io_ci = io_pp_23[14]; // @[wallace.scala 71:19]
  assign FullAdder_105_io_a = io_pp_24[13]; // @[wallace.scala 69:18]
  assign FullAdder_105_io_b = io_pp_25[12]; // @[wallace.scala 70:18]
  assign FullAdder_105_io_ci = io_pp_26[11]; // @[wallace.scala 71:19]
  assign FullAdder_106_io_a = io_pp_27[10]; // @[wallace.scala 69:18]
  assign FullAdder_106_io_b = io_pp_28[9]; // @[wallace.scala 70:18]
  assign FullAdder_106_io_ci = io_pp_29[8]; // @[wallace.scala 71:19]
  assign FullAdder_107_io_a = io_pp_5[31]; // @[wallace.scala 69:18]
  assign FullAdder_107_io_b = io_pp_6[30]; // @[wallace.scala 70:18]
  assign FullAdder_107_io_ci = io_pp_7[29]; // @[wallace.scala 71:19]
  assign FullAdder_108_io_a = io_pp_8[28]; // @[wallace.scala 69:18]
  assign FullAdder_108_io_b = io_pp_9[27]; // @[wallace.scala 70:18]
  assign FullAdder_108_io_ci = io_pp_10[26]; // @[wallace.scala 71:19]
  assign FullAdder_109_io_a = io_pp_11[25]; // @[wallace.scala 69:18]
  assign FullAdder_109_io_b = io_pp_12[24]; // @[wallace.scala 70:18]
  assign FullAdder_109_io_ci = io_pp_13[23]; // @[wallace.scala 71:19]
  assign FullAdder_110_io_a = io_pp_14[22]; // @[wallace.scala 69:18]
  assign FullAdder_110_io_b = io_pp_15[21]; // @[wallace.scala 70:18]
  assign FullAdder_110_io_ci = io_pp_16[20]; // @[wallace.scala 71:19]
  assign FullAdder_111_io_a = io_pp_17[19]; // @[wallace.scala 69:18]
  assign FullAdder_111_io_b = io_pp_18[18]; // @[wallace.scala 70:18]
  assign FullAdder_111_io_ci = io_pp_19[17]; // @[wallace.scala 71:19]
  assign FullAdder_112_io_a = io_pp_20[16]; // @[wallace.scala 69:18]
  assign FullAdder_112_io_b = io_pp_21[15]; // @[wallace.scala 70:18]
  assign FullAdder_112_io_ci = io_pp_22[14]; // @[wallace.scala 71:19]
  assign FullAdder_113_io_a = io_pp_23[13]; // @[wallace.scala 69:18]
  assign FullAdder_113_io_b = io_pp_24[12]; // @[wallace.scala 70:18]
  assign FullAdder_113_io_ci = io_pp_25[11]; // @[wallace.scala 71:19]
  assign FullAdder_114_io_a = io_pp_26[10]; // @[wallace.scala 69:18]
  assign FullAdder_114_io_b = io_pp_27[9]; // @[wallace.scala 70:18]
  assign FullAdder_114_io_ci = io_pp_28[8]; // @[wallace.scala 71:19]
  assign FullAdder_115_io_a = io_pp_29[7]; // @[wallace.scala 69:18]
  assign FullAdder_115_io_b = io_pp_30[6]; // @[wallace.scala 70:18]
  assign FullAdder_115_io_ci = io_pp_31[5]; // @[wallace.scala 71:19]
  assign FullAdder_116_io_a = io_pp_4[31]; // @[wallace.scala 69:18]
  assign FullAdder_116_io_b = io_pp_5[30]; // @[wallace.scala 70:18]
  assign FullAdder_116_io_ci = io_pp_6[29]; // @[wallace.scala 71:19]
  assign FullAdder_117_io_a = io_pp_7[28]; // @[wallace.scala 69:18]
  assign FullAdder_117_io_b = io_pp_8[27]; // @[wallace.scala 70:18]
  assign FullAdder_117_io_ci = io_pp_9[26]; // @[wallace.scala 71:19]
  assign FullAdder_118_io_a = io_pp_10[25]; // @[wallace.scala 69:18]
  assign FullAdder_118_io_b = io_pp_11[24]; // @[wallace.scala 70:18]
  assign FullAdder_118_io_ci = io_pp_12[23]; // @[wallace.scala 71:19]
  assign FullAdder_119_io_a = io_pp_13[22]; // @[wallace.scala 69:18]
  assign FullAdder_119_io_b = io_pp_14[21]; // @[wallace.scala 70:18]
  assign FullAdder_119_io_ci = io_pp_15[20]; // @[wallace.scala 71:19]
  assign FullAdder_120_io_a = io_pp_16[19]; // @[wallace.scala 69:18]
  assign FullAdder_120_io_b = io_pp_17[18]; // @[wallace.scala 70:18]
  assign FullAdder_120_io_ci = io_pp_18[17]; // @[wallace.scala 71:19]
  assign FullAdder_121_io_a = io_pp_19[16]; // @[wallace.scala 69:18]
  assign FullAdder_121_io_b = io_pp_20[15]; // @[wallace.scala 70:18]
  assign FullAdder_121_io_ci = io_pp_21[14]; // @[wallace.scala 71:19]
  assign FullAdder_122_io_a = io_pp_22[13]; // @[wallace.scala 69:18]
  assign FullAdder_122_io_b = io_pp_23[12]; // @[wallace.scala 70:18]
  assign FullAdder_122_io_ci = io_pp_24[11]; // @[wallace.scala 71:19]
  assign FullAdder_123_io_a = io_pp_25[10]; // @[wallace.scala 69:18]
  assign FullAdder_123_io_b = io_pp_26[9]; // @[wallace.scala 70:18]
  assign FullAdder_123_io_ci = io_pp_27[8]; // @[wallace.scala 71:19]
  assign FullAdder_124_io_a = io_pp_28[7]; // @[wallace.scala 69:18]
  assign FullAdder_124_io_b = io_pp_29[6]; // @[wallace.scala 70:18]
  assign FullAdder_124_io_ci = io_pp_30[5]; // @[wallace.scala 71:19]
  assign FullAdder_125_io_a = io_pp_3[31]; // @[wallace.scala 69:18]
  assign FullAdder_125_io_b = io_pp_4[30]; // @[wallace.scala 70:18]
  assign FullAdder_125_io_ci = io_pp_5[29]; // @[wallace.scala 71:19]
  assign FullAdder_126_io_a = io_pp_6[28]; // @[wallace.scala 69:18]
  assign FullAdder_126_io_b = io_pp_7[27]; // @[wallace.scala 70:18]
  assign FullAdder_126_io_ci = io_pp_8[26]; // @[wallace.scala 71:19]
  assign FullAdder_127_io_a = io_pp_9[25]; // @[wallace.scala 69:18]
  assign FullAdder_127_io_b = io_pp_10[24]; // @[wallace.scala 70:18]
  assign FullAdder_127_io_ci = io_pp_11[23]; // @[wallace.scala 71:19]
  assign FullAdder_128_io_a = io_pp_12[22]; // @[wallace.scala 69:18]
  assign FullAdder_128_io_b = io_pp_13[21]; // @[wallace.scala 70:18]
  assign FullAdder_128_io_ci = io_pp_14[20]; // @[wallace.scala 71:19]
  assign FullAdder_129_io_a = io_pp_15[19]; // @[wallace.scala 69:18]
  assign FullAdder_129_io_b = io_pp_16[18]; // @[wallace.scala 70:18]
  assign FullAdder_129_io_ci = io_pp_17[17]; // @[wallace.scala 71:19]
  assign FullAdder_130_io_a = io_pp_18[16]; // @[wallace.scala 69:18]
  assign FullAdder_130_io_b = io_pp_19[15]; // @[wallace.scala 70:18]
  assign FullAdder_130_io_ci = io_pp_20[14]; // @[wallace.scala 71:19]
  assign FullAdder_131_io_a = io_pp_21[13]; // @[wallace.scala 69:18]
  assign FullAdder_131_io_b = io_pp_22[12]; // @[wallace.scala 70:18]
  assign FullAdder_131_io_ci = io_pp_23[11]; // @[wallace.scala 71:19]
  assign FullAdder_132_io_a = io_pp_24[10]; // @[wallace.scala 69:18]
  assign FullAdder_132_io_b = io_pp_25[9]; // @[wallace.scala 70:18]
  assign FullAdder_132_io_ci = io_pp_26[8]; // @[wallace.scala 71:19]
  assign FullAdder_133_io_a = io_pp_27[7]; // @[wallace.scala 69:18]
  assign FullAdder_133_io_b = io_pp_28[6]; // @[wallace.scala 70:18]
  assign FullAdder_133_io_ci = io_pp_29[5]; // @[wallace.scala 71:19]
  assign HalfAdder_7_io_a = io_pp_30[4]; // @[wallace.scala 59:18]
  assign HalfAdder_7_io_b = io_pp_31[3]; // @[wallace.scala 60:18]
  assign FullAdder_134_io_a = io_pp_2[31]; // @[wallace.scala 69:18]
  assign FullAdder_134_io_b = io_pp_3[30]; // @[wallace.scala 70:18]
  assign FullAdder_134_io_ci = io_pp_4[29]; // @[wallace.scala 71:19]
  assign FullAdder_135_io_a = io_pp_5[28]; // @[wallace.scala 69:18]
  assign FullAdder_135_io_b = io_pp_6[27]; // @[wallace.scala 70:18]
  assign FullAdder_135_io_ci = io_pp_7[26]; // @[wallace.scala 71:19]
  assign FullAdder_136_io_a = io_pp_8[25]; // @[wallace.scala 69:18]
  assign FullAdder_136_io_b = io_pp_9[24]; // @[wallace.scala 70:18]
  assign FullAdder_136_io_ci = io_pp_10[23]; // @[wallace.scala 71:19]
  assign FullAdder_137_io_a = io_pp_11[22]; // @[wallace.scala 69:18]
  assign FullAdder_137_io_b = io_pp_12[21]; // @[wallace.scala 70:18]
  assign FullAdder_137_io_ci = io_pp_13[20]; // @[wallace.scala 71:19]
  assign FullAdder_138_io_a = io_pp_14[19]; // @[wallace.scala 69:18]
  assign FullAdder_138_io_b = io_pp_15[18]; // @[wallace.scala 70:18]
  assign FullAdder_138_io_ci = io_pp_16[17]; // @[wallace.scala 71:19]
  assign FullAdder_139_io_a = io_pp_17[16]; // @[wallace.scala 69:18]
  assign FullAdder_139_io_b = io_pp_18[15]; // @[wallace.scala 70:18]
  assign FullAdder_139_io_ci = io_pp_19[14]; // @[wallace.scala 71:19]
  assign FullAdder_140_io_a = io_pp_20[13]; // @[wallace.scala 69:18]
  assign FullAdder_140_io_b = io_pp_21[12]; // @[wallace.scala 70:18]
  assign FullAdder_140_io_ci = io_pp_22[11]; // @[wallace.scala 71:19]
  assign FullAdder_141_io_a = io_pp_23[10]; // @[wallace.scala 69:18]
  assign FullAdder_141_io_b = io_pp_24[9]; // @[wallace.scala 70:18]
  assign FullAdder_141_io_ci = io_pp_25[8]; // @[wallace.scala 71:19]
  assign FullAdder_142_io_a = io_pp_26[7]; // @[wallace.scala 69:18]
  assign FullAdder_142_io_b = io_pp_27[6]; // @[wallace.scala 70:18]
  assign FullAdder_142_io_ci = io_pp_28[5]; // @[wallace.scala 71:19]
  assign FullAdder_143_io_a = io_pp_29[4]; // @[wallace.scala 69:18]
  assign FullAdder_143_io_b = io_pp_30[3]; // @[wallace.scala 70:18]
  assign FullAdder_143_io_ci = io_pp_31[2]; // @[wallace.scala 71:19]
  assign FullAdder_144_io_a = io_pp_1[31]; // @[wallace.scala 69:18]
  assign FullAdder_144_io_b = io_pp_2[30]; // @[wallace.scala 70:18]
  assign FullAdder_144_io_ci = io_pp_3[29]; // @[wallace.scala 71:19]
  assign FullAdder_145_io_a = io_pp_4[28]; // @[wallace.scala 69:18]
  assign FullAdder_145_io_b = io_pp_5[27]; // @[wallace.scala 70:18]
  assign FullAdder_145_io_ci = io_pp_6[26]; // @[wallace.scala 71:19]
  assign FullAdder_146_io_a = io_pp_7[25]; // @[wallace.scala 69:18]
  assign FullAdder_146_io_b = io_pp_8[24]; // @[wallace.scala 70:18]
  assign FullAdder_146_io_ci = io_pp_9[23]; // @[wallace.scala 71:19]
  assign FullAdder_147_io_a = io_pp_10[22]; // @[wallace.scala 69:18]
  assign FullAdder_147_io_b = io_pp_11[21]; // @[wallace.scala 70:18]
  assign FullAdder_147_io_ci = io_pp_12[20]; // @[wallace.scala 71:19]
  assign FullAdder_148_io_a = io_pp_13[19]; // @[wallace.scala 69:18]
  assign FullAdder_148_io_b = io_pp_14[18]; // @[wallace.scala 70:18]
  assign FullAdder_148_io_ci = io_pp_15[17]; // @[wallace.scala 71:19]
  assign FullAdder_149_io_a = io_pp_16[16]; // @[wallace.scala 69:18]
  assign FullAdder_149_io_b = io_pp_17[15]; // @[wallace.scala 70:18]
  assign FullAdder_149_io_ci = io_pp_18[14]; // @[wallace.scala 71:19]
  assign FullAdder_150_io_a = io_pp_19[13]; // @[wallace.scala 69:18]
  assign FullAdder_150_io_b = io_pp_20[12]; // @[wallace.scala 70:18]
  assign FullAdder_150_io_ci = io_pp_21[11]; // @[wallace.scala 71:19]
  assign FullAdder_151_io_a = io_pp_22[10]; // @[wallace.scala 69:18]
  assign FullAdder_151_io_b = io_pp_23[9]; // @[wallace.scala 70:18]
  assign FullAdder_151_io_ci = io_pp_24[8]; // @[wallace.scala 71:19]
  assign FullAdder_152_io_a = io_pp_25[7]; // @[wallace.scala 69:18]
  assign FullAdder_152_io_b = io_pp_26[6]; // @[wallace.scala 70:18]
  assign FullAdder_152_io_ci = io_pp_27[5]; // @[wallace.scala 71:19]
  assign FullAdder_153_io_a = io_pp_28[4]; // @[wallace.scala 69:18]
  assign FullAdder_153_io_b = io_pp_29[3]; // @[wallace.scala 70:18]
  assign FullAdder_153_io_ci = io_pp_30[2]; // @[wallace.scala 71:19]
  assign FullAdder_154_io_a = io_pp_0[31]; // @[wallace.scala 69:18]
  assign FullAdder_154_io_b = io_pp_1[30]; // @[wallace.scala 70:18]
  assign FullAdder_154_io_ci = io_pp_2[29]; // @[wallace.scala 71:19]
  assign FullAdder_155_io_a = io_pp_3[28]; // @[wallace.scala 69:18]
  assign FullAdder_155_io_b = io_pp_4[27]; // @[wallace.scala 70:18]
  assign FullAdder_155_io_ci = io_pp_5[26]; // @[wallace.scala 71:19]
  assign FullAdder_156_io_a = io_pp_6[25]; // @[wallace.scala 69:18]
  assign FullAdder_156_io_b = io_pp_7[24]; // @[wallace.scala 70:18]
  assign FullAdder_156_io_ci = io_pp_8[23]; // @[wallace.scala 71:19]
  assign FullAdder_157_io_a = io_pp_9[22]; // @[wallace.scala 69:18]
  assign FullAdder_157_io_b = io_pp_10[21]; // @[wallace.scala 70:18]
  assign FullAdder_157_io_ci = io_pp_11[20]; // @[wallace.scala 71:19]
  assign FullAdder_158_io_a = io_pp_12[19]; // @[wallace.scala 69:18]
  assign FullAdder_158_io_b = io_pp_13[18]; // @[wallace.scala 70:18]
  assign FullAdder_158_io_ci = io_pp_14[17]; // @[wallace.scala 71:19]
  assign FullAdder_159_io_a = io_pp_15[16]; // @[wallace.scala 69:18]
  assign FullAdder_159_io_b = io_pp_16[15]; // @[wallace.scala 70:18]
  assign FullAdder_159_io_ci = io_pp_17[14]; // @[wallace.scala 71:19]
  assign FullAdder_160_io_a = io_pp_18[13]; // @[wallace.scala 69:18]
  assign FullAdder_160_io_b = io_pp_19[12]; // @[wallace.scala 70:18]
  assign FullAdder_160_io_ci = io_pp_20[11]; // @[wallace.scala 71:19]
  assign FullAdder_161_io_a = io_pp_21[10]; // @[wallace.scala 69:18]
  assign FullAdder_161_io_b = io_pp_22[9]; // @[wallace.scala 70:18]
  assign FullAdder_161_io_ci = io_pp_23[8]; // @[wallace.scala 71:19]
  assign FullAdder_162_io_a = io_pp_24[7]; // @[wallace.scala 69:18]
  assign FullAdder_162_io_b = io_pp_25[6]; // @[wallace.scala 70:18]
  assign FullAdder_162_io_ci = io_pp_26[5]; // @[wallace.scala 71:19]
  assign FullAdder_163_io_a = io_pp_27[4]; // @[wallace.scala 69:18]
  assign FullAdder_163_io_b = io_pp_28[3]; // @[wallace.scala 70:18]
  assign FullAdder_163_io_ci = io_pp_29[2]; // @[wallace.scala 71:19]
  assign FullAdder_164_io_a = io_pp_0[30]; // @[wallace.scala 69:18]
  assign FullAdder_164_io_b = io_pp_1[29]; // @[wallace.scala 70:18]
  assign FullAdder_164_io_ci = io_pp_2[28]; // @[wallace.scala 71:19]
  assign FullAdder_165_io_a = io_pp_3[27]; // @[wallace.scala 69:18]
  assign FullAdder_165_io_b = io_pp_4[26]; // @[wallace.scala 70:18]
  assign FullAdder_165_io_ci = io_pp_5[25]; // @[wallace.scala 71:19]
  assign FullAdder_166_io_a = io_pp_6[24]; // @[wallace.scala 69:18]
  assign FullAdder_166_io_b = io_pp_7[23]; // @[wallace.scala 70:18]
  assign FullAdder_166_io_ci = io_pp_8[22]; // @[wallace.scala 71:19]
  assign FullAdder_167_io_a = io_pp_9[21]; // @[wallace.scala 69:18]
  assign FullAdder_167_io_b = io_pp_10[20]; // @[wallace.scala 70:18]
  assign FullAdder_167_io_ci = io_pp_11[19]; // @[wallace.scala 71:19]
  assign FullAdder_168_io_a = io_pp_12[18]; // @[wallace.scala 69:18]
  assign FullAdder_168_io_b = io_pp_13[17]; // @[wallace.scala 70:18]
  assign FullAdder_168_io_ci = io_pp_14[16]; // @[wallace.scala 71:19]
  assign FullAdder_169_io_a = io_pp_15[15]; // @[wallace.scala 69:18]
  assign FullAdder_169_io_b = io_pp_16[14]; // @[wallace.scala 70:18]
  assign FullAdder_169_io_ci = io_pp_17[13]; // @[wallace.scala 71:19]
  assign FullAdder_170_io_a = io_pp_18[12]; // @[wallace.scala 69:18]
  assign FullAdder_170_io_b = io_pp_19[11]; // @[wallace.scala 70:18]
  assign FullAdder_170_io_ci = io_pp_20[10]; // @[wallace.scala 71:19]
  assign FullAdder_171_io_a = io_pp_21[9]; // @[wallace.scala 69:18]
  assign FullAdder_171_io_b = io_pp_22[8]; // @[wallace.scala 70:18]
  assign FullAdder_171_io_ci = io_pp_23[7]; // @[wallace.scala 71:19]
  assign FullAdder_172_io_a = io_pp_24[6]; // @[wallace.scala 69:18]
  assign FullAdder_172_io_b = io_pp_25[5]; // @[wallace.scala 70:18]
  assign FullAdder_172_io_ci = io_pp_26[4]; // @[wallace.scala 71:19]
  assign FullAdder_173_io_a = io_pp_27[3]; // @[wallace.scala 69:18]
  assign FullAdder_173_io_b = io_pp_28[2]; // @[wallace.scala 70:18]
  assign FullAdder_173_io_ci = io_pp_29[1]; // @[wallace.scala 71:19]
  assign FullAdder_174_io_a = io_pp_0[29]; // @[wallace.scala 69:18]
  assign FullAdder_174_io_b = io_pp_1[28]; // @[wallace.scala 70:18]
  assign FullAdder_174_io_ci = io_pp_2[27]; // @[wallace.scala 71:19]
  assign FullAdder_175_io_a = io_pp_3[26]; // @[wallace.scala 69:18]
  assign FullAdder_175_io_b = io_pp_4[25]; // @[wallace.scala 70:18]
  assign FullAdder_175_io_ci = io_pp_5[24]; // @[wallace.scala 71:19]
  assign FullAdder_176_io_a = io_pp_6[23]; // @[wallace.scala 69:18]
  assign FullAdder_176_io_b = io_pp_7[22]; // @[wallace.scala 70:18]
  assign FullAdder_176_io_ci = io_pp_8[21]; // @[wallace.scala 71:19]
  assign FullAdder_177_io_a = io_pp_9[20]; // @[wallace.scala 69:18]
  assign FullAdder_177_io_b = io_pp_10[19]; // @[wallace.scala 70:18]
  assign FullAdder_177_io_ci = io_pp_11[18]; // @[wallace.scala 71:19]
  assign FullAdder_178_io_a = io_pp_12[17]; // @[wallace.scala 69:18]
  assign FullAdder_178_io_b = io_pp_13[16]; // @[wallace.scala 70:18]
  assign FullAdder_178_io_ci = io_pp_14[15]; // @[wallace.scala 71:19]
  assign FullAdder_179_io_a = io_pp_15[14]; // @[wallace.scala 69:18]
  assign FullAdder_179_io_b = io_pp_16[13]; // @[wallace.scala 70:18]
  assign FullAdder_179_io_ci = io_pp_17[12]; // @[wallace.scala 71:19]
  assign FullAdder_180_io_a = io_pp_18[11]; // @[wallace.scala 69:18]
  assign FullAdder_180_io_b = io_pp_19[10]; // @[wallace.scala 70:18]
  assign FullAdder_180_io_ci = io_pp_20[9]; // @[wallace.scala 71:19]
  assign FullAdder_181_io_a = io_pp_21[8]; // @[wallace.scala 69:18]
  assign FullAdder_181_io_b = io_pp_22[7]; // @[wallace.scala 70:18]
  assign FullAdder_181_io_ci = io_pp_23[6]; // @[wallace.scala 71:19]
  assign FullAdder_182_io_a = io_pp_24[5]; // @[wallace.scala 69:18]
  assign FullAdder_182_io_b = io_pp_25[4]; // @[wallace.scala 70:18]
  assign FullAdder_182_io_ci = io_pp_26[3]; // @[wallace.scala 71:19]
  assign FullAdder_183_io_a = io_pp_27[2]; // @[wallace.scala 69:18]
  assign FullAdder_183_io_b = io_pp_28[1]; // @[wallace.scala 70:18]
  assign FullAdder_183_io_ci = io_pp_29[0]; // @[wallace.scala 71:19]
  assign FullAdder_184_io_a = io_pp_0[28]; // @[wallace.scala 69:18]
  assign FullAdder_184_io_b = io_pp_1[27]; // @[wallace.scala 70:18]
  assign FullAdder_184_io_ci = io_pp_2[26]; // @[wallace.scala 71:19]
  assign FullAdder_185_io_a = io_pp_3[25]; // @[wallace.scala 69:18]
  assign FullAdder_185_io_b = io_pp_4[24]; // @[wallace.scala 70:18]
  assign FullAdder_185_io_ci = io_pp_5[23]; // @[wallace.scala 71:19]
  assign FullAdder_186_io_a = io_pp_6[22]; // @[wallace.scala 69:18]
  assign FullAdder_186_io_b = io_pp_7[21]; // @[wallace.scala 70:18]
  assign FullAdder_186_io_ci = io_pp_8[20]; // @[wallace.scala 71:19]
  assign FullAdder_187_io_a = io_pp_9[19]; // @[wallace.scala 69:18]
  assign FullAdder_187_io_b = io_pp_10[18]; // @[wallace.scala 70:18]
  assign FullAdder_187_io_ci = io_pp_11[17]; // @[wallace.scala 71:19]
  assign FullAdder_188_io_a = io_pp_12[16]; // @[wallace.scala 69:18]
  assign FullAdder_188_io_b = io_pp_13[15]; // @[wallace.scala 70:18]
  assign FullAdder_188_io_ci = io_pp_14[14]; // @[wallace.scala 71:19]
  assign FullAdder_189_io_a = io_pp_15[13]; // @[wallace.scala 69:18]
  assign FullAdder_189_io_b = io_pp_16[12]; // @[wallace.scala 70:18]
  assign FullAdder_189_io_ci = io_pp_17[11]; // @[wallace.scala 71:19]
  assign FullAdder_190_io_a = io_pp_18[10]; // @[wallace.scala 69:18]
  assign FullAdder_190_io_b = io_pp_19[9]; // @[wallace.scala 70:18]
  assign FullAdder_190_io_ci = io_pp_20[8]; // @[wallace.scala 71:19]
  assign FullAdder_191_io_a = io_pp_21[7]; // @[wallace.scala 69:18]
  assign FullAdder_191_io_b = io_pp_22[6]; // @[wallace.scala 70:18]
  assign FullAdder_191_io_ci = io_pp_23[5]; // @[wallace.scala 71:19]
  assign FullAdder_192_io_a = io_pp_24[4]; // @[wallace.scala 69:18]
  assign FullAdder_192_io_b = io_pp_25[3]; // @[wallace.scala 70:18]
  assign FullAdder_192_io_ci = io_pp_26[2]; // @[wallace.scala 71:19]
  assign HalfAdder_8_io_a = io_pp_27[1]; // @[wallace.scala 59:18]
  assign HalfAdder_8_io_b = io_pp_28[0]; // @[wallace.scala 60:18]
  assign FullAdder_193_io_a = io_pp_0[27]; // @[wallace.scala 69:18]
  assign FullAdder_193_io_b = io_pp_1[26]; // @[wallace.scala 70:18]
  assign FullAdder_193_io_ci = io_pp_2[25]; // @[wallace.scala 71:19]
  assign FullAdder_194_io_a = io_pp_3[24]; // @[wallace.scala 69:18]
  assign FullAdder_194_io_b = io_pp_4[23]; // @[wallace.scala 70:18]
  assign FullAdder_194_io_ci = io_pp_5[22]; // @[wallace.scala 71:19]
  assign FullAdder_195_io_a = io_pp_6[21]; // @[wallace.scala 69:18]
  assign FullAdder_195_io_b = io_pp_7[20]; // @[wallace.scala 70:18]
  assign FullAdder_195_io_ci = io_pp_8[19]; // @[wallace.scala 71:19]
  assign FullAdder_196_io_a = io_pp_9[18]; // @[wallace.scala 69:18]
  assign FullAdder_196_io_b = io_pp_10[17]; // @[wallace.scala 70:18]
  assign FullAdder_196_io_ci = io_pp_11[16]; // @[wallace.scala 71:19]
  assign FullAdder_197_io_a = io_pp_12[15]; // @[wallace.scala 69:18]
  assign FullAdder_197_io_b = io_pp_13[14]; // @[wallace.scala 70:18]
  assign FullAdder_197_io_ci = io_pp_14[13]; // @[wallace.scala 71:19]
  assign FullAdder_198_io_a = io_pp_15[12]; // @[wallace.scala 69:18]
  assign FullAdder_198_io_b = io_pp_16[11]; // @[wallace.scala 70:18]
  assign FullAdder_198_io_ci = io_pp_17[10]; // @[wallace.scala 71:19]
  assign FullAdder_199_io_a = io_pp_18[9]; // @[wallace.scala 69:18]
  assign FullAdder_199_io_b = io_pp_19[8]; // @[wallace.scala 70:18]
  assign FullAdder_199_io_ci = io_pp_20[7]; // @[wallace.scala 71:19]
  assign FullAdder_200_io_a = io_pp_21[6]; // @[wallace.scala 69:18]
  assign FullAdder_200_io_b = io_pp_22[5]; // @[wallace.scala 70:18]
  assign FullAdder_200_io_ci = io_pp_23[4]; // @[wallace.scala 71:19]
  assign FullAdder_201_io_a = io_pp_24[3]; // @[wallace.scala 69:18]
  assign FullAdder_201_io_b = io_pp_25[2]; // @[wallace.scala 70:18]
  assign FullAdder_201_io_ci = io_pp_26[1]; // @[wallace.scala 71:19]
  assign FullAdder_202_io_a = io_pp_0[26]; // @[wallace.scala 69:18]
  assign FullAdder_202_io_b = io_pp_1[25]; // @[wallace.scala 70:18]
  assign FullAdder_202_io_ci = io_pp_2[24]; // @[wallace.scala 71:19]
  assign FullAdder_203_io_a = io_pp_3[23]; // @[wallace.scala 69:18]
  assign FullAdder_203_io_b = io_pp_4[22]; // @[wallace.scala 70:18]
  assign FullAdder_203_io_ci = io_pp_5[21]; // @[wallace.scala 71:19]
  assign FullAdder_204_io_a = io_pp_6[20]; // @[wallace.scala 69:18]
  assign FullAdder_204_io_b = io_pp_7[19]; // @[wallace.scala 70:18]
  assign FullAdder_204_io_ci = io_pp_8[18]; // @[wallace.scala 71:19]
  assign FullAdder_205_io_a = io_pp_9[17]; // @[wallace.scala 69:18]
  assign FullAdder_205_io_b = io_pp_10[16]; // @[wallace.scala 70:18]
  assign FullAdder_205_io_ci = io_pp_11[15]; // @[wallace.scala 71:19]
  assign FullAdder_206_io_a = io_pp_12[14]; // @[wallace.scala 69:18]
  assign FullAdder_206_io_b = io_pp_13[13]; // @[wallace.scala 70:18]
  assign FullAdder_206_io_ci = io_pp_14[12]; // @[wallace.scala 71:19]
  assign FullAdder_207_io_a = io_pp_15[11]; // @[wallace.scala 69:18]
  assign FullAdder_207_io_b = io_pp_16[10]; // @[wallace.scala 70:18]
  assign FullAdder_207_io_ci = io_pp_17[9]; // @[wallace.scala 71:19]
  assign FullAdder_208_io_a = io_pp_18[8]; // @[wallace.scala 69:18]
  assign FullAdder_208_io_b = io_pp_19[7]; // @[wallace.scala 70:18]
  assign FullAdder_208_io_ci = io_pp_20[6]; // @[wallace.scala 71:19]
  assign FullAdder_209_io_a = io_pp_21[5]; // @[wallace.scala 69:18]
  assign FullAdder_209_io_b = io_pp_22[4]; // @[wallace.scala 70:18]
  assign FullAdder_209_io_ci = io_pp_23[3]; // @[wallace.scala 71:19]
  assign FullAdder_210_io_a = io_pp_24[2]; // @[wallace.scala 69:18]
  assign FullAdder_210_io_b = io_pp_25[1]; // @[wallace.scala 70:18]
  assign FullAdder_210_io_ci = io_pp_26[0]; // @[wallace.scala 71:19]
  assign FullAdder_211_io_a = io_pp_0[25]; // @[wallace.scala 69:18]
  assign FullAdder_211_io_b = io_pp_1[24]; // @[wallace.scala 70:18]
  assign FullAdder_211_io_ci = io_pp_2[23]; // @[wallace.scala 71:19]
  assign FullAdder_212_io_a = io_pp_3[22]; // @[wallace.scala 69:18]
  assign FullAdder_212_io_b = io_pp_4[21]; // @[wallace.scala 70:18]
  assign FullAdder_212_io_ci = io_pp_5[20]; // @[wallace.scala 71:19]
  assign FullAdder_213_io_a = io_pp_6[19]; // @[wallace.scala 69:18]
  assign FullAdder_213_io_b = io_pp_7[18]; // @[wallace.scala 70:18]
  assign FullAdder_213_io_ci = io_pp_8[17]; // @[wallace.scala 71:19]
  assign FullAdder_214_io_a = io_pp_9[16]; // @[wallace.scala 69:18]
  assign FullAdder_214_io_b = io_pp_10[15]; // @[wallace.scala 70:18]
  assign FullAdder_214_io_ci = io_pp_11[14]; // @[wallace.scala 71:19]
  assign FullAdder_215_io_a = io_pp_12[13]; // @[wallace.scala 69:18]
  assign FullAdder_215_io_b = io_pp_13[12]; // @[wallace.scala 70:18]
  assign FullAdder_215_io_ci = io_pp_14[11]; // @[wallace.scala 71:19]
  assign FullAdder_216_io_a = io_pp_15[10]; // @[wallace.scala 69:18]
  assign FullAdder_216_io_b = io_pp_16[9]; // @[wallace.scala 70:18]
  assign FullAdder_216_io_ci = io_pp_17[8]; // @[wallace.scala 71:19]
  assign FullAdder_217_io_a = io_pp_18[7]; // @[wallace.scala 69:18]
  assign FullAdder_217_io_b = io_pp_19[6]; // @[wallace.scala 70:18]
  assign FullAdder_217_io_ci = io_pp_20[5]; // @[wallace.scala 71:19]
  assign FullAdder_218_io_a = io_pp_21[4]; // @[wallace.scala 69:18]
  assign FullAdder_218_io_b = io_pp_22[3]; // @[wallace.scala 70:18]
  assign FullAdder_218_io_ci = io_pp_23[2]; // @[wallace.scala 71:19]
  assign HalfAdder_9_io_a = io_pp_24[1]; // @[wallace.scala 59:18]
  assign HalfAdder_9_io_b = io_pp_25[0]; // @[wallace.scala 60:18]
  assign FullAdder_219_io_a = io_pp_0[24]; // @[wallace.scala 69:18]
  assign FullAdder_219_io_b = io_pp_1[23]; // @[wallace.scala 70:18]
  assign FullAdder_219_io_ci = io_pp_2[22]; // @[wallace.scala 71:19]
  assign FullAdder_220_io_a = io_pp_3[21]; // @[wallace.scala 69:18]
  assign FullAdder_220_io_b = io_pp_4[20]; // @[wallace.scala 70:18]
  assign FullAdder_220_io_ci = io_pp_5[19]; // @[wallace.scala 71:19]
  assign FullAdder_221_io_a = io_pp_6[18]; // @[wallace.scala 69:18]
  assign FullAdder_221_io_b = io_pp_7[17]; // @[wallace.scala 70:18]
  assign FullAdder_221_io_ci = io_pp_8[16]; // @[wallace.scala 71:19]
  assign FullAdder_222_io_a = io_pp_9[15]; // @[wallace.scala 69:18]
  assign FullAdder_222_io_b = io_pp_10[14]; // @[wallace.scala 70:18]
  assign FullAdder_222_io_ci = io_pp_11[13]; // @[wallace.scala 71:19]
  assign FullAdder_223_io_a = io_pp_12[12]; // @[wallace.scala 69:18]
  assign FullAdder_223_io_b = io_pp_13[11]; // @[wallace.scala 70:18]
  assign FullAdder_223_io_ci = io_pp_14[10]; // @[wallace.scala 71:19]
  assign FullAdder_224_io_a = io_pp_15[9]; // @[wallace.scala 69:18]
  assign FullAdder_224_io_b = io_pp_16[8]; // @[wallace.scala 70:18]
  assign FullAdder_224_io_ci = io_pp_17[7]; // @[wallace.scala 71:19]
  assign FullAdder_225_io_a = io_pp_18[6]; // @[wallace.scala 69:18]
  assign FullAdder_225_io_b = io_pp_19[5]; // @[wallace.scala 70:18]
  assign FullAdder_225_io_ci = io_pp_20[4]; // @[wallace.scala 71:19]
  assign FullAdder_226_io_a = io_pp_21[3]; // @[wallace.scala 69:18]
  assign FullAdder_226_io_b = io_pp_22[2]; // @[wallace.scala 70:18]
  assign FullAdder_226_io_ci = io_pp_23[1]; // @[wallace.scala 71:19]
  assign FullAdder_227_io_a = io_pp_0[23]; // @[wallace.scala 69:18]
  assign FullAdder_227_io_b = io_pp_1[22]; // @[wallace.scala 70:18]
  assign FullAdder_227_io_ci = io_pp_2[21]; // @[wallace.scala 71:19]
  assign FullAdder_228_io_a = io_pp_3[20]; // @[wallace.scala 69:18]
  assign FullAdder_228_io_b = io_pp_4[19]; // @[wallace.scala 70:18]
  assign FullAdder_228_io_ci = io_pp_5[18]; // @[wallace.scala 71:19]
  assign FullAdder_229_io_a = io_pp_6[17]; // @[wallace.scala 69:18]
  assign FullAdder_229_io_b = io_pp_7[16]; // @[wallace.scala 70:18]
  assign FullAdder_229_io_ci = io_pp_8[15]; // @[wallace.scala 71:19]
  assign FullAdder_230_io_a = io_pp_9[14]; // @[wallace.scala 69:18]
  assign FullAdder_230_io_b = io_pp_10[13]; // @[wallace.scala 70:18]
  assign FullAdder_230_io_ci = io_pp_11[12]; // @[wallace.scala 71:19]
  assign FullAdder_231_io_a = io_pp_12[11]; // @[wallace.scala 69:18]
  assign FullAdder_231_io_b = io_pp_13[10]; // @[wallace.scala 70:18]
  assign FullAdder_231_io_ci = io_pp_14[9]; // @[wallace.scala 71:19]
  assign FullAdder_232_io_a = io_pp_15[8]; // @[wallace.scala 69:18]
  assign FullAdder_232_io_b = io_pp_16[7]; // @[wallace.scala 70:18]
  assign FullAdder_232_io_ci = io_pp_17[6]; // @[wallace.scala 71:19]
  assign FullAdder_233_io_a = io_pp_18[5]; // @[wallace.scala 69:18]
  assign FullAdder_233_io_b = io_pp_19[4]; // @[wallace.scala 70:18]
  assign FullAdder_233_io_ci = io_pp_20[3]; // @[wallace.scala 71:19]
  assign FullAdder_234_io_a = io_pp_21[2]; // @[wallace.scala 69:18]
  assign FullAdder_234_io_b = io_pp_22[1]; // @[wallace.scala 70:18]
  assign FullAdder_234_io_ci = io_pp_23[0]; // @[wallace.scala 71:19]
  assign FullAdder_235_io_a = io_pp_0[22]; // @[wallace.scala 69:18]
  assign FullAdder_235_io_b = io_pp_1[21]; // @[wallace.scala 70:18]
  assign FullAdder_235_io_ci = io_pp_2[20]; // @[wallace.scala 71:19]
  assign FullAdder_236_io_a = io_pp_3[19]; // @[wallace.scala 69:18]
  assign FullAdder_236_io_b = io_pp_4[18]; // @[wallace.scala 70:18]
  assign FullAdder_236_io_ci = io_pp_5[17]; // @[wallace.scala 71:19]
  assign FullAdder_237_io_a = io_pp_6[16]; // @[wallace.scala 69:18]
  assign FullAdder_237_io_b = io_pp_7[15]; // @[wallace.scala 70:18]
  assign FullAdder_237_io_ci = io_pp_8[14]; // @[wallace.scala 71:19]
  assign FullAdder_238_io_a = io_pp_9[13]; // @[wallace.scala 69:18]
  assign FullAdder_238_io_b = io_pp_10[12]; // @[wallace.scala 70:18]
  assign FullAdder_238_io_ci = io_pp_11[11]; // @[wallace.scala 71:19]
  assign FullAdder_239_io_a = io_pp_12[10]; // @[wallace.scala 69:18]
  assign FullAdder_239_io_b = io_pp_13[9]; // @[wallace.scala 70:18]
  assign FullAdder_239_io_ci = io_pp_14[8]; // @[wallace.scala 71:19]
  assign FullAdder_240_io_a = io_pp_15[7]; // @[wallace.scala 69:18]
  assign FullAdder_240_io_b = io_pp_16[6]; // @[wallace.scala 70:18]
  assign FullAdder_240_io_ci = io_pp_17[5]; // @[wallace.scala 71:19]
  assign FullAdder_241_io_a = io_pp_18[4]; // @[wallace.scala 69:18]
  assign FullAdder_241_io_b = io_pp_19[3]; // @[wallace.scala 70:18]
  assign FullAdder_241_io_ci = io_pp_20[2]; // @[wallace.scala 71:19]
  assign FullAdder_242_io_a = io_pp_0[21]; // @[wallace.scala 69:18]
  assign FullAdder_242_io_b = io_pp_1[20]; // @[wallace.scala 70:18]
  assign FullAdder_242_io_ci = io_pp_2[19]; // @[wallace.scala 71:19]
  assign FullAdder_243_io_a = io_pp_3[18]; // @[wallace.scala 69:18]
  assign FullAdder_243_io_b = io_pp_4[17]; // @[wallace.scala 70:18]
  assign FullAdder_243_io_ci = io_pp_5[16]; // @[wallace.scala 71:19]
  assign FullAdder_244_io_a = io_pp_6[15]; // @[wallace.scala 69:18]
  assign FullAdder_244_io_b = io_pp_7[14]; // @[wallace.scala 70:18]
  assign FullAdder_244_io_ci = io_pp_8[13]; // @[wallace.scala 71:19]
  assign FullAdder_245_io_a = io_pp_9[12]; // @[wallace.scala 69:18]
  assign FullAdder_245_io_b = io_pp_10[11]; // @[wallace.scala 70:18]
  assign FullAdder_245_io_ci = io_pp_11[10]; // @[wallace.scala 71:19]
  assign FullAdder_246_io_a = io_pp_12[9]; // @[wallace.scala 69:18]
  assign FullAdder_246_io_b = io_pp_13[8]; // @[wallace.scala 70:18]
  assign FullAdder_246_io_ci = io_pp_14[7]; // @[wallace.scala 71:19]
  assign FullAdder_247_io_a = io_pp_15[6]; // @[wallace.scala 69:18]
  assign FullAdder_247_io_b = io_pp_16[5]; // @[wallace.scala 70:18]
  assign FullAdder_247_io_ci = io_pp_17[4]; // @[wallace.scala 71:19]
  assign FullAdder_248_io_a = io_pp_18[3]; // @[wallace.scala 69:18]
  assign FullAdder_248_io_b = io_pp_19[2]; // @[wallace.scala 70:18]
  assign FullAdder_248_io_ci = io_pp_20[1]; // @[wallace.scala 71:19]
  assign FullAdder_249_io_a = io_pp_0[20]; // @[wallace.scala 69:18]
  assign FullAdder_249_io_b = io_pp_1[19]; // @[wallace.scala 70:18]
  assign FullAdder_249_io_ci = io_pp_2[18]; // @[wallace.scala 71:19]
  assign FullAdder_250_io_a = io_pp_3[17]; // @[wallace.scala 69:18]
  assign FullAdder_250_io_b = io_pp_4[16]; // @[wallace.scala 70:18]
  assign FullAdder_250_io_ci = io_pp_5[15]; // @[wallace.scala 71:19]
  assign FullAdder_251_io_a = io_pp_6[14]; // @[wallace.scala 69:18]
  assign FullAdder_251_io_b = io_pp_7[13]; // @[wallace.scala 70:18]
  assign FullAdder_251_io_ci = io_pp_8[12]; // @[wallace.scala 71:19]
  assign FullAdder_252_io_a = io_pp_9[11]; // @[wallace.scala 69:18]
  assign FullAdder_252_io_b = io_pp_10[10]; // @[wallace.scala 70:18]
  assign FullAdder_252_io_ci = io_pp_11[9]; // @[wallace.scala 71:19]
  assign FullAdder_253_io_a = io_pp_12[8]; // @[wallace.scala 69:18]
  assign FullAdder_253_io_b = io_pp_13[7]; // @[wallace.scala 70:18]
  assign FullAdder_253_io_ci = io_pp_14[6]; // @[wallace.scala 71:19]
  assign FullAdder_254_io_a = io_pp_15[5]; // @[wallace.scala 69:18]
  assign FullAdder_254_io_b = io_pp_16[4]; // @[wallace.scala 70:18]
  assign FullAdder_254_io_ci = io_pp_17[3]; // @[wallace.scala 71:19]
  assign FullAdder_255_io_a = io_pp_18[2]; // @[wallace.scala 69:18]
  assign FullAdder_255_io_b = io_pp_19[1]; // @[wallace.scala 70:18]
  assign FullAdder_255_io_ci = io_pp_20[0]; // @[wallace.scala 71:19]
  assign FullAdder_256_io_a = io_pp_0[19]; // @[wallace.scala 69:18]
  assign FullAdder_256_io_b = io_pp_1[18]; // @[wallace.scala 70:18]
  assign FullAdder_256_io_ci = io_pp_2[17]; // @[wallace.scala 71:19]
  assign FullAdder_257_io_a = io_pp_3[16]; // @[wallace.scala 69:18]
  assign FullAdder_257_io_b = io_pp_4[15]; // @[wallace.scala 70:18]
  assign FullAdder_257_io_ci = io_pp_5[14]; // @[wallace.scala 71:19]
  assign FullAdder_258_io_a = io_pp_6[13]; // @[wallace.scala 69:18]
  assign FullAdder_258_io_b = io_pp_7[12]; // @[wallace.scala 70:18]
  assign FullAdder_258_io_ci = io_pp_8[11]; // @[wallace.scala 71:19]
  assign FullAdder_259_io_a = io_pp_9[10]; // @[wallace.scala 69:18]
  assign FullAdder_259_io_b = io_pp_10[9]; // @[wallace.scala 70:18]
  assign FullAdder_259_io_ci = io_pp_11[8]; // @[wallace.scala 71:19]
  assign FullAdder_260_io_a = io_pp_12[7]; // @[wallace.scala 69:18]
  assign FullAdder_260_io_b = io_pp_13[6]; // @[wallace.scala 70:18]
  assign FullAdder_260_io_ci = io_pp_14[5]; // @[wallace.scala 71:19]
  assign FullAdder_261_io_a = io_pp_15[4]; // @[wallace.scala 69:18]
  assign FullAdder_261_io_b = io_pp_16[3]; // @[wallace.scala 70:18]
  assign FullAdder_261_io_ci = io_pp_17[2]; // @[wallace.scala 71:19]
  assign FullAdder_262_io_a = io_pp_0[18]; // @[wallace.scala 69:18]
  assign FullAdder_262_io_b = io_pp_1[17]; // @[wallace.scala 70:18]
  assign FullAdder_262_io_ci = io_pp_2[16]; // @[wallace.scala 71:19]
  assign FullAdder_263_io_a = io_pp_3[15]; // @[wallace.scala 69:18]
  assign FullAdder_263_io_b = io_pp_4[14]; // @[wallace.scala 70:18]
  assign FullAdder_263_io_ci = io_pp_5[13]; // @[wallace.scala 71:19]
  assign FullAdder_264_io_a = io_pp_6[12]; // @[wallace.scala 69:18]
  assign FullAdder_264_io_b = io_pp_7[11]; // @[wallace.scala 70:18]
  assign FullAdder_264_io_ci = io_pp_8[10]; // @[wallace.scala 71:19]
  assign FullAdder_265_io_a = io_pp_9[9]; // @[wallace.scala 69:18]
  assign FullAdder_265_io_b = io_pp_10[8]; // @[wallace.scala 70:18]
  assign FullAdder_265_io_ci = io_pp_11[7]; // @[wallace.scala 71:19]
  assign FullAdder_266_io_a = io_pp_12[6]; // @[wallace.scala 69:18]
  assign FullAdder_266_io_b = io_pp_13[5]; // @[wallace.scala 70:18]
  assign FullAdder_266_io_ci = io_pp_14[4]; // @[wallace.scala 71:19]
  assign FullAdder_267_io_a = io_pp_15[3]; // @[wallace.scala 69:18]
  assign FullAdder_267_io_b = io_pp_16[2]; // @[wallace.scala 70:18]
  assign FullAdder_267_io_ci = io_pp_17[1]; // @[wallace.scala 71:19]
  assign FullAdder_268_io_a = io_pp_0[17]; // @[wallace.scala 69:18]
  assign FullAdder_268_io_b = io_pp_1[16]; // @[wallace.scala 70:18]
  assign FullAdder_268_io_ci = io_pp_2[15]; // @[wallace.scala 71:19]
  assign FullAdder_269_io_a = io_pp_3[14]; // @[wallace.scala 69:18]
  assign FullAdder_269_io_b = io_pp_4[13]; // @[wallace.scala 70:18]
  assign FullAdder_269_io_ci = io_pp_5[12]; // @[wallace.scala 71:19]
  assign FullAdder_270_io_a = io_pp_6[11]; // @[wallace.scala 69:18]
  assign FullAdder_270_io_b = io_pp_7[10]; // @[wallace.scala 70:18]
  assign FullAdder_270_io_ci = io_pp_8[9]; // @[wallace.scala 71:19]
  assign FullAdder_271_io_a = io_pp_9[8]; // @[wallace.scala 69:18]
  assign FullAdder_271_io_b = io_pp_10[7]; // @[wallace.scala 70:18]
  assign FullAdder_271_io_ci = io_pp_11[6]; // @[wallace.scala 71:19]
  assign FullAdder_272_io_a = io_pp_12[5]; // @[wallace.scala 69:18]
  assign FullAdder_272_io_b = io_pp_13[4]; // @[wallace.scala 70:18]
  assign FullAdder_272_io_ci = io_pp_14[3]; // @[wallace.scala 71:19]
  assign FullAdder_273_io_a = io_pp_15[2]; // @[wallace.scala 69:18]
  assign FullAdder_273_io_b = io_pp_16[1]; // @[wallace.scala 70:18]
  assign FullAdder_273_io_ci = io_pp_17[0]; // @[wallace.scala 71:19]
  assign FullAdder_274_io_a = io_pp_0[16]; // @[wallace.scala 69:18]
  assign FullAdder_274_io_b = io_pp_1[15]; // @[wallace.scala 70:18]
  assign FullAdder_274_io_ci = io_pp_2[14]; // @[wallace.scala 71:19]
  assign FullAdder_275_io_a = io_pp_3[13]; // @[wallace.scala 69:18]
  assign FullAdder_275_io_b = io_pp_4[12]; // @[wallace.scala 70:18]
  assign FullAdder_275_io_ci = io_pp_5[11]; // @[wallace.scala 71:19]
  assign FullAdder_276_io_a = io_pp_6[10]; // @[wallace.scala 69:18]
  assign FullAdder_276_io_b = io_pp_7[9]; // @[wallace.scala 70:18]
  assign FullAdder_276_io_ci = io_pp_8[8]; // @[wallace.scala 71:19]
  assign FullAdder_277_io_a = io_pp_9[7]; // @[wallace.scala 69:18]
  assign FullAdder_277_io_b = io_pp_10[6]; // @[wallace.scala 70:18]
  assign FullAdder_277_io_ci = io_pp_11[5]; // @[wallace.scala 71:19]
  assign FullAdder_278_io_a = io_pp_12[4]; // @[wallace.scala 69:18]
  assign FullAdder_278_io_b = io_pp_13[3]; // @[wallace.scala 70:18]
  assign FullAdder_278_io_ci = io_pp_14[2]; // @[wallace.scala 71:19]
  assign HalfAdder_10_io_a = io_pp_15[1]; // @[wallace.scala 59:18]
  assign HalfAdder_10_io_b = io_pp_16[0]; // @[wallace.scala 60:18]
  assign FullAdder_279_io_a = io_pp_0[15]; // @[wallace.scala 69:18]
  assign FullAdder_279_io_b = io_pp_1[14]; // @[wallace.scala 70:18]
  assign FullAdder_279_io_ci = io_pp_2[13]; // @[wallace.scala 71:19]
  assign FullAdder_280_io_a = io_pp_3[12]; // @[wallace.scala 69:18]
  assign FullAdder_280_io_b = io_pp_4[11]; // @[wallace.scala 70:18]
  assign FullAdder_280_io_ci = io_pp_5[10]; // @[wallace.scala 71:19]
  assign FullAdder_281_io_a = io_pp_6[9]; // @[wallace.scala 69:18]
  assign FullAdder_281_io_b = io_pp_7[8]; // @[wallace.scala 70:18]
  assign FullAdder_281_io_ci = io_pp_8[7]; // @[wallace.scala 71:19]
  assign FullAdder_282_io_a = io_pp_9[6]; // @[wallace.scala 69:18]
  assign FullAdder_282_io_b = io_pp_10[5]; // @[wallace.scala 70:18]
  assign FullAdder_282_io_ci = io_pp_11[4]; // @[wallace.scala 71:19]
  assign FullAdder_283_io_a = io_pp_12[3]; // @[wallace.scala 69:18]
  assign FullAdder_283_io_b = io_pp_13[2]; // @[wallace.scala 70:18]
  assign FullAdder_283_io_ci = io_pp_14[1]; // @[wallace.scala 71:19]
  assign FullAdder_284_io_a = io_pp_0[14]; // @[wallace.scala 69:18]
  assign FullAdder_284_io_b = io_pp_1[13]; // @[wallace.scala 70:18]
  assign FullAdder_284_io_ci = io_pp_2[12]; // @[wallace.scala 71:19]
  assign FullAdder_285_io_a = io_pp_3[11]; // @[wallace.scala 69:18]
  assign FullAdder_285_io_b = io_pp_4[10]; // @[wallace.scala 70:18]
  assign FullAdder_285_io_ci = io_pp_5[9]; // @[wallace.scala 71:19]
  assign FullAdder_286_io_a = io_pp_6[8]; // @[wallace.scala 69:18]
  assign FullAdder_286_io_b = io_pp_7[7]; // @[wallace.scala 70:18]
  assign FullAdder_286_io_ci = io_pp_8[6]; // @[wallace.scala 71:19]
  assign FullAdder_287_io_a = io_pp_9[5]; // @[wallace.scala 69:18]
  assign FullAdder_287_io_b = io_pp_10[4]; // @[wallace.scala 70:18]
  assign FullAdder_287_io_ci = io_pp_11[3]; // @[wallace.scala 71:19]
  assign FullAdder_288_io_a = io_pp_12[2]; // @[wallace.scala 69:18]
  assign FullAdder_288_io_b = io_pp_13[1]; // @[wallace.scala 70:18]
  assign FullAdder_288_io_ci = io_pp_14[0]; // @[wallace.scala 71:19]
  assign FullAdder_289_io_a = io_pp_0[13]; // @[wallace.scala 69:18]
  assign FullAdder_289_io_b = io_pp_1[12]; // @[wallace.scala 70:18]
  assign FullAdder_289_io_ci = io_pp_2[11]; // @[wallace.scala 71:19]
  assign FullAdder_290_io_a = io_pp_3[10]; // @[wallace.scala 69:18]
  assign FullAdder_290_io_b = io_pp_4[9]; // @[wallace.scala 70:18]
  assign FullAdder_290_io_ci = io_pp_5[8]; // @[wallace.scala 71:19]
  assign FullAdder_291_io_a = io_pp_6[7]; // @[wallace.scala 69:18]
  assign FullAdder_291_io_b = io_pp_7[6]; // @[wallace.scala 70:18]
  assign FullAdder_291_io_ci = io_pp_8[5]; // @[wallace.scala 71:19]
  assign FullAdder_292_io_a = io_pp_9[4]; // @[wallace.scala 69:18]
  assign FullAdder_292_io_b = io_pp_10[3]; // @[wallace.scala 70:18]
  assign FullAdder_292_io_ci = io_pp_11[2]; // @[wallace.scala 71:19]
  assign FullAdder_293_io_a = io_pp_0[12]; // @[wallace.scala 69:18]
  assign FullAdder_293_io_b = io_pp_1[11]; // @[wallace.scala 70:18]
  assign FullAdder_293_io_ci = io_pp_2[10]; // @[wallace.scala 71:19]
  assign FullAdder_294_io_a = io_pp_3[9]; // @[wallace.scala 69:18]
  assign FullAdder_294_io_b = io_pp_4[8]; // @[wallace.scala 70:18]
  assign FullAdder_294_io_ci = io_pp_5[7]; // @[wallace.scala 71:19]
  assign FullAdder_295_io_a = io_pp_6[6]; // @[wallace.scala 69:18]
  assign FullAdder_295_io_b = io_pp_7[5]; // @[wallace.scala 70:18]
  assign FullAdder_295_io_ci = io_pp_8[4]; // @[wallace.scala 71:19]
  assign FullAdder_296_io_a = io_pp_9[3]; // @[wallace.scala 69:18]
  assign FullAdder_296_io_b = io_pp_10[2]; // @[wallace.scala 70:18]
  assign FullAdder_296_io_ci = io_pp_11[1]; // @[wallace.scala 71:19]
  assign FullAdder_297_io_a = io_pp_0[11]; // @[wallace.scala 69:18]
  assign FullAdder_297_io_b = io_pp_1[10]; // @[wallace.scala 70:18]
  assign FullAdder_297_io_ci = io_pp_2[9]; // @[wallace.scala 71:19]
  assign FullAdder_298_io_a = io_pp_3[8]; // @[wallace.scala 69:18]
  assign FullAdder_298_io_b = io_pp_4[7]; // @[wallace.scala 70:18]
  assign FullAdder_298_io_ci = io_pp_5[6]; // @[wallace.scala 71:19]
  assign FullAdder_299_io_a = io_pp_6[5]; // @[wallace.scala 69:18]
  assign FullAdder_299_io_b = io_pp_7[4]; // @[wallace.scala 70:18]
  assign FullAdder_299_io_ci = io_pp_8[3]; // @[wallace.scala 71:19]
  assign FullAdder_300_io_a = io_pp_9[2]; // @[wallace.scala 69:18]
  assign FullAdder_300_io_b = io_pp_10[1]; // @[wallace.scala 70:18]
  assign FullAdder_300_io_ci = io_pp_11[0]; // @[wallace.scala 71:19]
  assign FullAdder_301_io_a = io_pp_0[10]; // @[wallace.scala 69:18]
  assign FullAdder_301_io_b = io_pp_1[9]; // @[wallace.scala 70:18]
  assign FullAdder_301_io_ci = io_pp_2[8]; // @[wallace.scala 71:19]
  assign FullAdder_302_io_a = io_pp_3[7]; // @[wallace.scala 69:18]
  assign FullAdder_302_io_b = io_pp_4[6]; // @[wallace.scala 70:18]
  assign FullAdder_302_io_ci = io_pp_5[5]; // @[wallace.scala 71:19]
  assign FullAdder_303_io_a = io_pp_6[4]; // @[wallace.scala 69:18]
  assign FullAdder_303_io_b = io_pp_7[3]; // @[wallace.scala 70:18]
  assign FullAdder_303_io_ci = io_pp_8[2]; // @[wallace.scala 71:19]
  assign HalfAdder_11_io_a = io_pp_9[1]; // @[wallace.scala 59:18]
  assign HalfAdder_11_io_b = io_pp_10[0]; // @[wallace.scala 60:18]
  assign FullAdder_304_io_a = io_pp_0[9]; // @[wallace.scala 69:18]
  assign FullAdder_304_io_b = io_pp_1[8]; // @[wallace.scala 70:18]
  assign FullAdder_304_io_ci = io_pp_2[7]; // @[wallace.scala 71:19]
  assign FullAdder_305_io_a = io_pp_3[6]; // @[wallace.scala 69:18]
  assign FullAdder_305_io_b = io_pp_4[5]; // @[wallace.scala 70:18]
  assign FullAdder_305_io_ci = io_pp_5[4]; // @[wallace.scala 71:19]
  assign FullAdder_306_io_a = io_pp_6[3]; // @[wallace.scala 69:18]
  assign FullAdder_306_io_b = io_pp_7[2]; // @[wallace.scala 70:18]
  assign FullAdder_306_io_ci = io_pp_8[1]; // @[wallace.scala 71:19]
  assign FullAdder_307_io_a = io_pp_0[8]; // @[wallace.scala 69:18]
  assign FullAdder_307_io_b = io_pp_1[7]; // @[wallace.scala 70:18]
  assign FullAdder_307_io_ci = io_pp_2[6]; // @[wallace.scala 71:19]
  assign FullAdder_308_io_a = io_pp_3[5]; // @[wallace.scala 69:18]
  assign FullAdder_308_io_b = io_pp_4[4]; // @[wallace.scala 70:18]
  assign FullAdder_308_io_ci = io_pp_5[3]; // @[wallace.scala 71:19]
  assign FullAdder_309_io_a = io_pp_6[2]; // @[wallace.scala 69:18]
  assign FullAdder_309_io_b = io_pp_7[1]; // @[wallace.scala 70:18]
  assign FullAdder_309_io_ci = io_pp_8[0]; // @[wallace.scala 71:19]
  assign FullAdder_310_io_a = io_pp_0[7]; // @[wallace.scala 69:18]
  assign FullAdder_310_io_b = io_pp_1[6]; // @[wallace.scala 70:18]
  assign FullAdder_310_io_ci = io_pp_2[5]; // @[wallace.scala 71:19]
  assign FullAdder_311_io_a = io_pp_3[4]; // @[wallace.scala 69:18]
  assign FullAdder_311_io_b = io_pp_4[3]; // @[wallace.scala 70:18]
  assign FullAdder_311_io_ci = io_pp_5[2]; // @[wallace.scala 71:19]
  assign HalfAdder_12_io_a = io_pp_6[1]; // @[wallace.scala 59:18]
  assign HalfAdder_12_io_b = io_pp_7[0]; // @[wallace.scala 60:18]
  assign FullAdder_312_io_a = io_pp_0[6]; // @[wallace.scala 69:18]
  assign FullAdder_312_io_b = io_pp_1[5]; // @[wallace.scala 70:18]
  assign FullAdder_312_io_ci = io_pp_2[4]; // @[wallace.scala 71:19]
  assign FullAdder_313_io_a = io_pp_3[3]; // @[wallace.scala 69:18]
  assign FullAdder_313_io_b = io_pp_4[2]; // @[wallace.scala 70:18]
  assign FullAdder_313_io_ci = io_pp_5[1]; // @[wallace.scala 71:19]
  assign FullAdder_314_io_a = io_pp_0[5]; // @[wallace.scala 69:18]
  assign FullAdder_314_io_b = io_pp_1[4]; // @[wallace.scala 70:18]
  assign FullAdder_314_io_ci = io_pp_2[3]; // @[wallace.scala 71:19]
  assign FullAdder_315_io_a = io_pp_3[2]; // @[wallace.scala 69:18]
  assign FullAdder_315_io_b = io_pp_4[1]; // @[wallace.scala 70:18]
  assign FullAdder_315_io_ci = io_pp_5[0]; // @[wallace.scala 71:19]
  assign FullAdder_316_io_a = io_pp_0[4]; // @[wallace.scala 69:18]
  assign FullAdder_316_io_b = io_pp_1[3]; // @[wallace.scala 70:18]
  assign FullAdder_316_io_ci = io_pp_2[2]; // @[wallace.scala 71:19]
  assign HalfAdder_13_io_a = io_pp_3[1]; // @[wallace.scala 59:18]
  assign HalfAdder_13_io_b = io_pp_4[0]; // @[wallace.scala 60:18]
  assign FullAdder_317_io_a = io_pp_0[3]; // @[wallace.scala 69:18]
  assign FullAdder_317_io_b = io_pp_1[2]; // @[wallace.scala 70:18]
  assign FullAdder_317_io_ci = io_pp_2[1]; // @[wallace.scala 71:19]
  assign FullAdder_318_io_a = io_pp_0[2]; // @[wallace.scala 69:18]
  assign FullAdder_318_io_b = io_pp_1[1]; // @[wallace.scala 70:18]
  assign FullAdder_318_io_ci = io_pp_2[0]; // @[wallace.scala 71:19]
  assign HalfAdder_14_io_a = io_pp_31[31]; // @[wallace.scala 59:18]
  assign HalfAdder_14_io_b = HalfAdder_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_15_io_a = HalfAdder_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_15_io_b = HalfAdder_1_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_16_io_a = io_pp_31[29]; // @[wallace.scala 59:18]
  assign HalfAdder_16_io_b = HalfAdder_1_io_s; // @[wallace.scala 60:18]
  assign FullAdder_319_io_a = io_pp_31[28]; // @[wallace.scala 69:18]
  assign FullAdder_319_io_b = FullAdder_io_s; // @[wallace.scala 70:18]
  assign FullAdder_319_io_ci = FullAdder_1_io_co; // @[wallace.scala 71:19]
  assign FullAdder_320_io_a = FullAdder_1_io_s; // @[wallace.scala 69:18]
  assign FullAdder_320_io_b = HalfAdder_2_io_s; // @[wallace.scala 70:18]
  assign FullAdder_320_io_ci = FullAdder_2_io_co; // @[wallace.scala 71:19]
  assign FullAdder_321_io_a = FullAdder_2_io_s; // @[wallace.scala 69:18]
  assign FullAdder_321_io_b = FullAdder_3_io_s; // @[wallace.scala 70:18]
  assign FullAdder_321_io_ci = FullAdder_4_io_co; // @[wallace.scala 71:19]
  assign FullAdder_322_io_a = io_pp_31[25]; // @[wallace.scala 69:18]
  assign FullAdder_322_io_b = FullAdder_4_io_s; // @[wallace.scala 70:18]
  assign FullAdder_322_io_ci = FullAdder_5_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_17_io_a = FullAdder_6_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_17_io_b = FullAdder_7_io_co; // @[wallace.scala 60:18]
  assign FullAdder_323_io_a = io_pp_30[25]; // @[wallace.scala 69:18]
  assign FullAdder_323_io_b = io_pp_31[24]; // @[wallace.scala 70:18]
  assign FullAdder_323_io_ci = FullAdder_6_io_s; // @[wallace.scala 71:19]
  assign FullAdder_324_io_a = FullAdder_7_io_s; // @[wallace.scala 69:18]
  assign FullAdder_324_io_b = FullAdder_8_io_co; // @[wallace.scala 70:18]
  assign FullAdder_324_io_ci = FullAdder_9_io_co; // @[wallace.scala 71:19]
  assign FullAdder_325_io_a = FullAdder_8_io_s; // @[wallace.scala 69:18]
  assign FullAdder_325_io_b = FullAdder_9_io_s; // @[wallace.scala 70:18]
  assign FullAdder_325_io_ci = FullAdder_10_io_s; // @[wallace.scala 71:19]
  assign FullAdder_326_io_a = FullAdder_11_io_co; // @[wallace.scala 69:18]
  assign FullAdder_326_io_b = FullAdder_12_io_co; // @[wallace.scala 70:18]
  assign FullAdder_326_io_ci = FullAdder_13_io_co; // @[wallace.scala 71:19]
  assign FullAdder_327_io_a = io_pp_31[22]; // @[wallace.scala 69:18]
  assign FullAdder_327_io_b = FullAdder_11_io_s; // @[wallace.scala 70:18]
  assign FullAdder_327_io_ci = FullAdder_12_io_s; // @[wallace.scala 71:19]
  assign FullAdder_328_io_a = FullAdder_13_io_s; // @[wallace.scala 69:18]
  assign FullAdder_328_io_b = FullAdder_14_io_co; // @[wallace.scala 70:18]
  assign FullAdder_328_io_ci = FullAdder_15_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_18_io_a = FullAdder_16_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_18_io_b = HalfAdder_3_io_co; // @[wallace.scala 60:18]
  assign FullAdder_329_io_a = FullAdder_14_io_s; // @[wallace.scala 69:18]
  assign FullAdder_329_io_b = FullAdder_15_io_s; // @[wallace.scala 70:18]
  assign FullAdder_329_io_ci = FullAdder_16_io_s; // @[wallace.scala 71:19]
  assign FullAdder_330_io_a = HalfAdder_3_io_s; // @[wallace.scala 69:18]
  assign FullAdder_330_io_b = FullAdder_17_io_co; // @[wallace.scala 70:18]
  assign FullAdder_330_io_ci = FullAdder_18_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_19_io_a = FullAdder_19_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_19_io_b = FullAdder_20_io_co; // @[wallace.scala 60:18]
  assign FullAdder_331_io_a = FullAdder_17_io_s; // @[wallace.scala 69:18]
  assign FullAdder_331_io_b = FullAdder_18_io_s; // @[wallace.scala 70:18]
  assign FullAdder_331_io_ci = FullAdder_19_io_s; // @[wallace.scala 71:19]
  assign FullAdder_332_io_a = FullAdder_20_io_s; // @[wallace.scala 69:18]
  assign FullAdder_332_io_b = FullAdder_21_io_co; // @[wallace.scala 70:18]
  assign FullAdder_332_io_ci = FullAdder_22_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_20_io_a = FullAdder_23_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_20_io_b = FullAdder_24_io_co; // @[wallace.scala 60:18]
  assign FullAdder_333_io_a = io_pp_31[19]; // @[wallace.scala 69:18]
  assign FullAdder_333_io_b = FullAdder_21_io_s; // @[wallace.scala 70:18]
  assign FullAdder_333_io_ci = FullAdder_22_io_s; // @[wallace.scala 71:19]
  assign FullAdder_334_io_a = FullAdder_23_io_s; // @[wallace.scala 69:18]
  assign FullAdder_334_io_b = FullAdder_24_io_s; // @[wallace.scala 70:18]
  assign FullAdder_334_io_ci = FullAdder_25_io_co; // @[wallace.scala 71:19]
  assign FullAdder_335_io_a = FullAdder_26_io_co; // @[wallace.scala 69:18]
  assign FullAdder_335_io_b = FullAdder_27_io_co; // @[wallace.scala 70:18]
  assign FullAdder_335_io_ci = FullAdder_28_io_co; // @[wallace.scala 71:19]
  assign FullAdder_336_io_a = FullAdder_25_io_s; // @[wallace.scala 69:18]
  assign FullAdder_336_io_b = FullAdder_26_io_s; // @[wallace.scala 70:18]
  assign FullAdder_336_io_ci = FullAdder_27_io_s; // @[wallace.scala 71:19]
  assign FullAdder_337_io_a = FullAdder_28_io_s; // @[wallace.scala 69:18]
  assign FullAdder_337_io_b = HalfAdder_4_io_s; // @[wallace.scala 70:18]
  assign FullAdder_337_io_ci = FullAdder_29_io_co; // @[wallace.scala 71:19]
  assign FullAdder_338_io_a = FullAdder_30_io_co; // @[wallace.scala 69:18]
  assign FullAdder_338_io_b = FullAdder_31_io_co; // @[wallace.scala 70:18]
  assign FullAdder_338_io_ci = FullAdder_32_io_co; // @[wallace.scala 71:19]
  assign FullAdder_339_io_a = FullAdder_29_io_s; // @[wallace.scala 69:18]
  assign FullAdder_339_io_b = FullAdder_30_io_s; // @[wallace.scala 70:18]
  assign FullAdder_339_io_ci = FullAdder_31_io_s; // @[wallace.scala 71:19]
  assign FullAdder_340_io_a = FullAdder_32_io_s; // @[wallace.scala 69:18]
  assign FullAdder_340_io_b = FullAdder_33_io_s; // @[wallace.scala 70:18]
  assign FullAdder_340_io_ci = FullAdder_34_io_co; // @[wallace.scala 71:19]
  assign FullAdder_341_io_a = FullAdder_35_io_co; // @[wallace.scala 69:18]
  assign FullAdder_341_io_b = FullAdder_36_io_co; // @[wallace.scala 70:18]
  assign FullAdder_341_io_ci = FullAdder_37_io_co; // @[wallace.scala 71:19]
  assign FullAdder_342_io_a = io_pp_31[16]; // @[wallace.scala 69:18]
  assign FullAdder_342_io_b = FullAdder_34_io_s; // @[wallace.scala 70:18]
  assign FullAdder_342_io_ci = FullAdder_35_io_s; // @[wallace.scala 71:19]
  assign FullAdder_343_io_a = FullAdder_36_io_s; // @[wallace.scala 69:18]
  assign FullAdder_343_io_b = FullAdder_37_io_s; // @[wallace.scala 70:18]
  assign FullAdder_343_io_ci = FullAdder_38_io_s; // @[wallace.scala 71:19]
  assign FullAdder_344_io_a = FullAdder_39_io_co; // @[wallace.scala 69:18]
  assign FullAdder_344_io_b = FullAdder_40_io_co; // @[wallace.scala 70:18]
  assign FullAdder_344_io_ci = FullAdder_41_io_co; // @[wallace.scala 71:19]
  assign FullAdder_345_io_a = FullAdder_42_io_co; // @[wallace.scala 69:18]
  assign FullAdder_345_io_b = FullAdder_43_io_co; // @[wallace.scala 70:18]
  assign FullAdder_345_io_ci = HalfAdder_5_io_co; // @[wallace.scala 71:19]
  assign FullAdder_346_io_a = FullAdder_39_io_s; // @[wallace.scala 69:18]
  assign FullAdder_346_io_b = FullAdder_40_io_s; // @[wallace.scala 70:18]
  assign FullAdder_346_io_ci = FullAdder_41_io_s; // @[wallace.scala 71:19]
  assign FullAdder_347_io_a = FullAdder_42_io_s; // @[wallace.scala 69:18]
  assign FullAdder_347_io_b = FullAdder_43_io_s; // @[wallace.scala 70:18]
  assign FullAdder_347_io_ci = HalfAdder_5_io_s; // @[wallace.scala 71:19]
  assign FullAdder_348_io_a = FullAdder_44_io_co; // @[wallace.scala 69:18]
  assign FullAdder_348_io_b = FullAdder_45_io_co; // @[wallace.scala 70:18]
  assign FullAdder_348_io_ci = FullAdder_46_io_co; // @[wallace.scala 71:19]
  assign FullAdder_349_io_a = FullAdder_47_io_co; // @[wallace.scala 69:18]
  assign FullAdder_349_io_b = FullAdder_48_io_co; // @[wallace.scala 70:18]
  assign FullAdder_349_io_ci = FullAdder_49_io_co; // @[wallace.scala 71:19]
  assign FullAdder_350_io_a = FullAdder_44_io_s; // @[wallace.scala 69:18]
  assign FullAdder_350_io_b = FullAdder_45_io_s; // @[wallace.scala 70:18]
  assign FullAdder_350_io_ci = FullAdder_46_io_s; // @[wallace.scala 71:19]
  assign FullAdder_351_io_a = FullAdder_47_io_s; // @[wallace.scala 69:18]
  assign FullAdder_351_io_b = FullAdder_48_io_s; // @[wallace.scala 70:18]
  assign FullAdder_351_io_ci = FullAdder_49_io_s; // @[wallace.scala 71:19]
  assign FullAdder_352_io_a = FullAdder_50_io_co; // @[wallace.scala 69:18]
  assign FullAdder_352_io_b = FullAdder_51_io_co; // @[wallace.scala 70:18]
  assign FullAdder_352_io_ci = FullAdder_52_io_co; // @[wallace.scala 71:19]
  assign FullAdder_353_io_a = FullAdder_53_io_co; // @[wallace.scala 69:18]
  assign FullAdder_353_io_b = FullAdder_54_io_co; // @[wallace.scala 70:18]
  assign FullAdder_353_io_ci = FullAdder_55_io_co; // @[wallace.scala 71:19]
  assign FullAdder_354_io_a = io_pp_31[13]; // @[wallace.scala 69:18]
  assign FullAdder_354_io_b = FullAdder_50_io_s; // @[wallace.scala 70:18]
  assign FullAdder_354_io_ci = FullAdder_51_io_s; // @[wallace.scala 71:19]
  assign FullAdder_355_io_a = FullAdder_52_io_s; // @[wallace.scala 69:18]
  assign FullAdder_355_io_b = FullAdder_53_io_s; // @[wallace.scala 70:18]
  assign FullAdder_355_io_ci = FullAdder_54_io_s; // @[wallace.scala 71:19]
  assign FullAdder_356_io_a = FullAdder_55_io_s; // @[wallace.scala 69:18]
  assign FullAdder_356_io_b = FullAdder_56_io_co; // @[wallace.scala 70:18]
  assign FullAdder_356_io_ci = FullAdder_57_io_co; // @[wallace.scala 71:19]
  assign FullAdder_357_io_a = FullAdder_58_io_co; // @[wallace.scala 69:18]
  assign FullAdder_357_io_b = FullAdder_59_io_co; // @[wallace.scala 70:18]
  assign FullAdder_357_io_ci = FullAdder_60_io_co; // @[wallace.scala 71:19]
  assign FullAdder_358_io_a = io_pp_30[13]; // @[wallace.scala 69:18]
  assign FullAdder_358_io_b = io_pp_31[12]; // @[wallace.scala 70:18]
  assign FullAdder_358_io_ci = FullAdder_56_io_s; // @[wallace.scala 71:19]
  assign FullAdder_359_io_a = FullAdder_57_io_s; // @[wallace.scala 69:18]
  assign FullAdder_359_io_b = FullAdder_58_io_s; // @[wallace.scala 70:18]
  assign FullAdder_359_io_ci = FullAdder_59_io_s; // @[wallace.scala 71:19]
  assign FullAdder_360_io_a = FullAdder_60_io_s; // @[wallace.scala 69:18]
  assign FullAdder_360_io_b = FullAdder_61_io_s; // @[wallace.scala 70:18]
  assign FullAdder_360_io_ci = FullAdder_62_io_co; // @[wallace.scala 71:19]
  assign FullAdder_361_io_a = FullAdder_63_io_co; // @[wallace.scala 69:18]
  assign FullAdder_361_io_b = FullAdder_64_io_co; // @[wallace.scala 70:18]
  assign FullAdder_361_io_ci = FullAdder_65_io_co; // @[wallace.scala 71:19]
  assign FullAdder_362_io_a = FullAdder_66_io_co; // @[wallace.scala 69:18]
  assign FullAdder_362_io_b = FullAdder_67_io_co; // @[wallace.scala 70:18]
  assign FullAdder_362_io_ci = FullAdder_68_io_co; // @[wallace.scala 71:19]
  assign FullAdder_363_io_a = FullAdder_62_io_s; // @[wallace.scala 69:18]
  assign FullAdder_363_io_b = FullAdder_63_io_s; // @[wallace.scala 70:18]
  assign FullAdder_363_io_ci = FullAdder_64_io_s; // @[wallace.scala 71:19]
  assign FullAdder_364_io_a = FullAdder_65_io_s; // @[wallace.scala 69:18]
  assign FullAdder_364_io_b = FullAdder_66_io_s; // @[wallace.scala 70:18]
  assign FullAdder_364_io_ci = FullAdder_67_io_s; // @[wallace.scala 71:19]
  assign FullAdder_365_io_a = FullAdder_68_io_s; // @[wallace.scala 69:18]
  assign FullAdder_365_io_b = FullAdder_69_io_co; // @[wallace.scala 70:18]
  assign FullAdder_365_io_ci = FullAdder_70_io_co; // @[wallace.scala 71:19]
  assign FullAdder_366_io_a = FullAdder_71_io_co; // @[wallace.scala 69:18]
  assign FullAdder_366_io_b = FullAdder_72_io_co; // @[wallace.scala 70:18]
  assign FullAdder_366_io_ci = FullAdder_73_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_21_io_a = FullAdder_74_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_21_io_b = FullAdder_75_io_co; // @[wallace.scala 60:18]
  assign FullAdder_367_io_a = io_pp_31[10]; // @[wallace.scala 69:18]
  assign FullAdder_367_io_b = FullAdder_69_io_s; // @[wallace.scala 70:18]
  assign FullAdder_367_io_ci = FullAdder_70_io_s; // @[wallace.scala 71:19]
  assign FullAdder_368_io_a = FullAdder_71_io_s; // @[wallace.scala 69:18]
  assign FullAdder_368_io_b = FullAdder_72_io_s; // @[wallace.scala 70:18]
  assign FullAdder_368_io_ci = FullAdder_73_io_s; // @[wallace.scala 71:19]
  assign FullAdder_369_io_a = FullAdder_74_io_s; // @[wallace.scala 69:18]
  assign FullAdder_369_io_b = FullAdder_75_io_s; // @[wallace.scala 70:18]
  assign FullAdder_369_io_ci = FullAdder_76_io_co; // @[wallace.scala 71:19]
  assign FullAdder_370_io_a = FullAdder_77_io_co; // @[wallace.scala 69:18]
  assign FullAdder_370_io_b = FullAdder_78_io_co; // @[wallace.scala 70:18]
  assign FullAdder_370_io_ci = FullAdder_79_io_co; // @[wallace.scala 71:19]
  assign FullAdder_371_io_a = FullAdder_80_io_co; // @[wallace.scala 69:18]
  assign FullAdder_371_io_b = FullAdder_81_io_co; // @[wallace.scala 70:18]
  assign FullAdder_371_io_ci = FullAdder_82_io_co; // @[wallace.scala 71:19]
  assign FullAdder_372_io_a = FullAdder_76_io_s; // @[wallace.scala 69:18]
  assign FullAdder_372_io_b = FullAdder_77_io_s; // @[wallace.scala 70:18]
  assign FullAdder_372_io_ci = FullAdder_78_io_s; // @[wallace.scala 71:19]
  assign FullAdder_373_io_a = FullAdder_79_io_s; // @[wallace.scala 69:18]
  assign FullAdder_373_io_b = FullAdder_80_io_s; // @[wallace.scala 70:18]
  assign FullAdder_373_io_ci = FullAdder_81_io_s; // @[wallace.scala 71:19]
  assign FullAdder_374_io_a = FullAdder_82_io_s; // @[wallace.scala 69:18]
  assign FullAdder_374_io_b = HalfAdder_6_io_s; // @[wallace.scala 70:18]
  assign FullAdder_374_io_ci = FullAdder_83_io_co; // @[wallace.scala 71:19]
  assign FullAdder_375_io_a = FullAdder_84_io_co; // @[wallace.scala 69:18]
  assign FullAdder_375_io_b = FullAdder_85_io_co; // @[wallace.scala 70:18]
  assign FullAdder_375_io_ci = FullAdder_86_io_co; // @[wallace.scala 71:19]
  assign FullAdder_376_io_a = FullAdder_87_io_co; // @[wallace.scala 69:18]
  assign FullAdder_376_io_b = FullAdder_88_io_co; // @[wallace.scala 70:18]
  assign FullAdder_376_io_ci = FullAdder_89_io_co; // @[wallace.scala 71:19]
  assign FullAdder_377_io_a = FullAdder_83_io_s; // @[wallace.scala 69:18]
  assign FullAdder_377_io_b = FullAdder_84_io_s; // @[wallace.scala 70:18]
  assign FullAdder_377_io_ci = FullAdder_85_io_s; // @[wallace.scala 71:19]
  assign FullAdder_378_io_a = FullAdder_86_io_s; // @[wallace.scala 69:18]
  assign FullAdder_378_io_b = FullAdder_87_io_s; // @[wallace.scala 70:18]
  assign FullAdder_378_io_ci = FullAdder_88_io_s; // @[wallace.scala 71:19]
  assign FullAdder_379_io_a = FullAdder_89_io_s; // @[wallace.scala 69:18]
  assign FullAdder_379_io_b = FullAdder_90_io_s; // @[wallace.scala 70:18]
  assign FullAdder_379_io_ci = FullAdder_91_io_co; // @[wallace.scala 71:19]
  assign FullAdder_380_io_a = FullAdder_92_io_co; // @[wallace.scala 69:18]
  assign FullAdder_380_io_b = FullAdder_93_io_co; // @[wallace.scala 70:18]
  assign FullAdder_380_io_ci = FullAdder_94_io_co; // @[wallace.scala 71:19]
  assign FullAdder_381_io_a = FullAdder_95_io_co; // @[wallace.scala 69:18]
  assign FullAdder_381_io_b = FullAdder_96_io_co; // @[wallace.scala 70:18]
  assign FullAdder_381_io_ci = FullAdder_97_io_co; // @[wallace.scala 71:19]
  assign FullAdder_382_io_a = io_pp_31[7]; // @[wallace.scala 69:18]
  assign FullAdder_382_io_b = FullAdder_91_io_s; // @[wallace.scala 70:18]
  assign FullAdder_382_io_ci = FullAdder_92_io_s; // @[wallace.scala 71:19]
  assign FullAdder_383_io_a = FullAdder_93_io_s; // @[wallace.scala 69:18]
  assign FullAdder_383_io_b = FullAdder_94_io_s; // @[wallace.scala 70:18]
  assign FullAdder_383_io_ci = FullAdder_95_io_s; // @[wallace.scala 71:19]
  assign FullAdder_384_io_a = FullAdder_96_io_s; // @[wallace.scala 69:18]
  assign FullAdder_384_io_b = FullAdder_97_io_s; // @[wallace.scala 70:18]
  assign FullAdder_384_io_ci = FullAdder_98_io_s; // @[wallace.scala 71:19]
  assign FullAdder_385_io_a = FullAdder_99_io_co; // @[wallace.scala 69:18]
  assign FullAdder_385_io_b = FullAdder_100_io_co; // @[wallace.scala 70:18]
  assign FullAdder_385_io_ci = FullAdder_101_io_co; // @[wallace.scala 71:19]
  assign FullAdder_386_io_a = FullAdder_102_io_co; // @[wallace.scala 69:18]
  assign FullAdder_386_io_b = FullAdder_103_io_co; // @[wallace.scala 70:18]
  assign FullAdder_386_io_ci = FullAdder_104_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_22_io_a = FullAdder_105_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_22_io_b = FullAdder_106_io_co; // @[wallace.scala 60:18]
  assign FullAdder_387_io_a = io_pp_30[7]; // @[wallace.scala 69:18]
  assign FullAdder_387_io_b = io_pp_31[6]; // @[wallace.scala 70:18]
  assign FullAdder_387_io_ci = FullAdder_99_io_s; // @[wallace.scala 71:19]
  assign FullAdder_388_io_a = FullAdder_100_io_s; // @[wallace.scala 69:18]
  assign FullAdder_388_io_b = FullAdder_101_io_s; // @[wallace.scala 70:18]
  assign FullAdder_388_io_ci = FullAdder_102_io_s; // @[wallace.scala 71:19]
  assign FullAdder_389_io_a = FullAdder_103_io_s; // @[wallace.scala 69:18]
  assign FullAdder_389_io_b = FullAdder_104_io_s; // @[wallace.scala 70:18]
  assign FullAdder_389_io_ci = FullAdder_105_io_s; // @[wallace.scala 71:19]
  assign FullAdder_390_io_a = FullAdder_106_io_s; // @[wallace.scala 69:18]
  assign FullAdder_390_io_b = FullAdder_107_io_co; // @[wallace.scala 70:18]
  assign FullAdder_390_io_ci = FullAdder_108_io_co; // @[wallace.scala 71:19]
  assign FullAdder_391_io_a = FullAdder_109_io_co; // @[wallace.scala 69:18]
  assign FullAdder_391_io_b = FullAdder_110_io_co; // @[wallace.scala 70:18]
  assign FullAdder_391_io_ci = FullAdder_111_io_co; // @[wallace.scala 71:19]
  assign FullAdder_392_io_a = FullAdder_112_io_co; // @[wallace.scala 69:18]
  assign FullAdder_392_io_b = FullAdder_113_io_co; // @[wallace.scala 70:18]
  assign FullAdder_392_io_ci = FullAdder_114_io_co; // @[wallace.scala 71:19]
  assign FullAdder_393_io_a = FullAdder_107_io_s; // @[wallace.scala 69:18]
  assign FullAdder_393_io_b = FullAdder_108_io_s; // @[wallace.scala 70:18]
  assign FullAdder_393_io_ci = FullAdder_109_io_s; // @[wallace.scala 71:19]
  assign FullAdder_394_io_a = FullAdder_110_io_s; // @[wallace.scala 69:18]
  assign FullAdder_394_io_b = FullAdder_111_io_s; // @[wallace.scala 70:18]
  assign FullAdder_394_io_ci = FullAdder_112_io_s; // @[wallace.scala 71:19]
  assign FullAdder_395_io_a = FullAdder_113_io_s; // @[wallace.scala 69:18]
  assign FullAdder_395_io_b = FullAdder_114_io_s; // @[wallace.scala 70:18]
  assign FullAdder_395_io_ci = FullAdder_115_io_s; // @[wallace.scala 71:19]
  assign FullAdder_396_io_a = FullAdder_116_io_co; // @[wallace.scala 69:18]
  assign FullAdder_396_io_b = FullAdder_117_io_co; // @[wallace.scala 70:18]
  assign FullAdder_396_io_ci = FullAdder_118_io_co; // @[wallace.scala 71:19]
  assign FullAdder_397_io_a = FullAdder_119_io_co; // @[wallace.scala 69:18]
  assign FullAdder_397_io_b = FullAdder_120_io_co; // @[wallace.scala 70:18]
  assign FullAdder_397_io_ci = FullAdder_121_io_co; // @[wallace.scala 71:19]
  assign FullAdder_398_io_a = FullAdder_122_io_co; // @[wallace.scala 69:18]
  assign FullAdder_398_io_b = FullAdder_123_io_co; // @[wallace.scala 70:18]
  assign FullAdder_398_io_ci = FullAdder_124_io_co; // @[wallace.scala 71:19]
  assign FullAdder_399_io_a = io_pp_31[4]; // @[wallace.scala 69:18]
  assign FullAdder_399_io_b = FullAdder_116_io_s; // @[wallace.scala 70:18]
  assign FullAdder_399_io_ci = FullAdder_117_io_s; // @[wallace.scala 71:19]
  assign FullAdder_400_io_a = FullAdder_118_io_s; // @[wallace.scala 69:18]
  assign FullAdder_400_io_b = FullAdder_119_io_s; // @[wallace.scala 70:18]
  assign FullAdder_400_io_ci = FullAdder_120_io_s; // @[wallace.scala 71:19]
  assign FullAdder_401_io_a = FullAdder_121_io_s; // @[wallace.scala 69:18]
  assign FullAdder_401_io_b = FullAdder_122_io_s; // @[wallace.scala 70:18]
  assign FullAdder_401_io_ci = FullAdder_123_io_s; // @[wallace.scala 71:19]
  assign FullAdder_402_io_a = FullAdder_124_io_s; // @[wallace.scala 69:18]
  assign FullAdder_402_io_b = FullAdder_125_io_co; // @[wallace.scala 70:18]
  assign FullAdder_402_io_ci = FullAdder_126_io_co; // @[wallace.scala 71:19]
  assign FullAdder_403_io_a = FullAdder_127_io_co; // @[wallace.scala 69:18]
  assign FullAdder_403_io_b = FullAdder_128_io_co; // @[wallace.scala 70:18]
  assign FullAdder_403_io_ci = FullAdder_129_io_co; // @[wallace.scala 71:19]
  assign FullAdder_404_io_a = FullAdder_130_io_co; // @[wallace.scala 69:18]
  assign FullAdder_404_io_b = FullAdder_131_io_co; // @[wallace.scala 70:18]
  assign FullAdder_404_io_ci = FullAdder_132_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_23_io_a = FullAdder_133_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_23_io_b = HalfAdder_7_io_co; // @[wallace.scala 60:18]
  assign FullAdder_405_io_a = FullAdder_125_io_s; // @[wallace.scala 69:18]
  assign FullAdder_405_io_b = FullAdder_126_io_s; // @[wallace.scala 70:18]
  assign FullAdder_405_io_ci = FullAdder_127_io_s; // @[wallace.scala 71:19]
  assign FullAdder_406_io_a = FullAdder_128_io_s; // @[wallace.scala 69:18]
  assign FullAdder_406_io_b = FullAdder_129_io_s; // @[wallace.scala 70:18]
  assign FullAdder_406_io_ci = FullAdder_130_io_s; // @[wallace.scala 71:19]
  assign FullAdder_407_io_a = FullAdder_131_io_s; // @[wallace.scala 69:18]
  assign FullAdder_407_io_b = FullAdder_132_io_s; // @[wallace.scala 70:18]
  assign FullAdder_407_io_ci = FullAdder_133_io_s; // @[wallace.scala 71:19]
  assign FullAdder_408_io_a = HalfAdder_7_io_s; // @[wallace.scala 69:18]
  assign FullAdder_408_io_b = FullAdder_134_io_co; // @[wallace.scala 70:18]
  assign FullAdder_408_io_ci = FullAdder_135_io_co; // @[wallace.scala 71:19]
  assign FullAdder_409_io_a = FullAdder_136_io_co; // @[wallace.scala 69:18]
  assign FullAdder_409_io_b = FullAdder_137_io_co; // @[wallace.scala 70:18]
  assign FullAdder_409_io_ci = FullAdder_138_io_co; // @[wallace.scala 71:19]
  assign FullAdder_410_io_a = FullAdder_139_io_co; // @[wallace.scala 69:18]
  assign FullAdder_410_io_b = FullAdder_140_io_co; // @[wallace.scala 70:18]
  assign FullAdder_410_io_ci = FullAdder_141_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_24_io_a = FullAdder_142_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_24_io_b = FullAdder_143_io_co; // @[wallace.scala 60:18]
  assign FullAdder_411_io_a = FullAdder_134_io_s; // @[wallace.scala 69:18]
  assign FullAdder_411_io_b = FullAdder_135_io_s; // @[wallace.scala 70:18]
  assign FullAdder_411_io_ci = FullAdder_136_io_s; // @[wallace.scala 71:19]
  assign FullAdder_412_io_a = FullAdder_137_io_s; // @[wallace.scala 69:18]
  assign FullAdder_412_io_b = FullAdder_138_io_s; // @[wallace.scala 70:18]
  assign FullAdder_412_io_ci = FullAdder_139_io_s; // @[wallace.scala 71:19]
  assign FullAdder_413_io_a = FullAdder_140_io_s; // @[wallace.scala 69:18]
  assign FullAdder_413_io_b = FullAdder_141_io_s; // @[wallace.scala 70:18]
  assign FullAdder_413_io_ci = FullAdder_142_io_s; // @[wallace.scala 71:19]
  assign FullAdder_414_io_a = FullAdder_143_io_s; // @[wallace.scala 69:18]
  assign FullAdder_414_io_b = FullAdder_144_io_co; // @[wallace.scala 70:18]
  assign FullAdder_414_io_ci = FullAdder_145_io_co; // @[wallace.scala 71:19]
  assign FullAdder_415_io_a = FullAdder_146_io_co; // @[wallace.scala 69:18]
  assign FullAdder_415_io_b = FullAdder_147_io_co; // @[wallace.scala 70:18]
  assign FullAdder_415_io_ci = FullAdder_148_io_co; // @[wallace.scala 71:19]
  assign FullAdder_416_io_a = FullAdder_149_io_co; // @[wallace.scala 69:18]
  assign FullAdder_416_io_b = FullAdder_150_io_co; // @[wallace.scala 70:18]
  assign FullAdder_416_io_ci = FullAdder_151_io_co; // @[wallace.scala 71:19]
  assign FullAdder_417_io_a = io_pp_31[1]; // @[wallace.scala 69:18]
  assign FullAdder_417_io_b = FullAdder_144_io_s; // @[wallace.scala 70:18]
  assign FullAdder_417_io_ci = FullAdder_145_io_s; // @[wallace.scala 71:19]
  assign FullAdder_418_io_a = FullAdder_146_io_s; // @[wallace.scala 69:18]
  assign FullAdder_418_io_b = FullAdder_147_io_s; // @[wallace.scala 70:18]
  assign FullAdder_418_io_ci = FullAdder_148_io_s; // @[wallace.scala 71:19]
  assign FullAdder_419_io_a = FullAdder_149_io_s; // @[wallace.scala 69:18]
  assign FullAdder_419_io_b = FullAdder_150_io_s; // @[wallace.scala 70:18]
  assign FullAdder_419_io_ci = FullAdder_151_io_s; // @[wallace.scala 71:19]
  assign FullAdder_420_io_a = FullAdder_152_io_s; // @[wallace.scala 69:18]
  assign FullAdder_420_io_b = FullAdder_153_io_s; // @[wallace.scala 70:18]
  assign FullAdder_420_io_ci = FullAdder_154_io_co; // @[wallace.scala 71:19]
  assign FullAdder_421_io_a = FullAdder_155_io_co; // @[wallace.scala 69:18]
  assign FullAdder_421_io_b = FullAdder_156_io_co; // @[wallace.scala 70:18]
  assign FullAdder_421_io_ci = FullAdder_157_io_co; // @[wallace.scala 71:19]
  assign FullAdder_422_io_a = FullAdder_158_io_co; // @[wallace.scala 69:18]
  assign FullAdder_422_io_b = FullAdder_159_io_co; // @[wallace.scala 70:18]
  assign FullAdder_422_io_ci = FullAdder_160_io_co; // @[wallace.scala 71:19]
  assign FullAdder_423_io_a = FullAdder_161_io_co; // @[wallace.scala 69:18]
  assign FullAdder_423_io_b = FullAdder_162_io_co; // @[wallace.scala 70:18]
  assign FullAdder_423_io_ci = FullAdder_163_io_co; // @[wallace.scala 71:19]
  assign FullAdder_424_io_a = io_pp_30[1]; // @[wallace.scala 69:18]
  assign FullAdder_424_io_b = io_pp_31[0]; // @[wallace.scala 70:18]
  assign FullAdder_424_io_ci = FullAdder_154_io_s; // @[wallace.scala 71:19]
  assign FullAdder_425_io_a = FullAdder_155_io_s; // @[wallace.scala 69:18]
  assign FullAdder_425_io_b = FullAdder_156_io_s; // @[wallace.scala 70:18]
  assign FullAdder_425_io_ci = FullAdder_157_io_s; // @[wallace.scala 71:19]
  assign FullAdder_426_io_a = FullAdder_158_io_s; // @[wallace.scala 69:18]
  assign FullAdder_426_io_b = FullAdder_159_io_s; // @[wallace.scala 70:18]
  assign FullAdder_426_io_ci = FullAdder_160_io_s; // @[wallace.scala 71:19]
  assign FullAdder_427_io_a = FullAdder_161_io_s; // @[wallace.scala 69:18]
  assign FullAdder_427_io_b = FullAdder_162_io_s; // @[wallace.scala 70:18]
  assign FullAdder_427_io_ci = FullAdder_163_io_s; // @[wallace.scala 71:19]
  assign FullAdder_428_io_a = FullAdder_164_io_co; // @[wallace.scala 69:18]
  assign FullAdder_428_io_b = FullAdder_165_io_co; // @[wallace.scala 70:18]
  assign FullAdder_428_io_ci = FullAdder_166_io_co; // @[wallace.scala 71:19]
  assign FullAdder_429_io_a = FullAdder_167_io_co; // @[wallace.scala 69:18]
  assign FullAdder_429_io_b = FullAdder_168_io_co; // @[wallace.scala 70:18]
  assign FullAdder_429_io_ci = FullAdder_169_io_co; // @[wallace.scala 71:19]
  assign FullAdder_430_io_a = FullAdder_170_io_co; // @[wallace.scala 69:18]
  assign FullAdder_430_io_b = FullAdder_171_io_co; // @[wallace.scala 70:18]
  assign FullAdder_430_io_ci = FullAdder_172_io_co; // @[wallace.scala 71:19]
  assign FullAdder_431_io_a = io_pp_30[0]; // @[wallace.scala 69:18]
  assign FullAdder_431_io_b = FullAdder_164_io_s; // @[wallace.scala 70:18]
  assign FullAdder_431_io_ci = FullAdder_165_io_s; // @[wallace.scala 71:19]
  assign FullAdder_432_io_a = FullAdder_166_io_s; // @[wallace.scala 69:18]
  assign FullAdder_432_io_b = FullAdder_167_io_s; // @[wallace.scala 70:18]
  assign FullAdder_432_io_ci = FullAdder_168_io_s; // @[wallace.scala 71:19]
  assign FullAdder_433_io_a = FullAdder_169_io_s; // @[wallace.scala 69:18]
  assign FullAdder_433_io_b = FullAdder_170_io_s; // @[wallace.scala 70:18]
  assign FullAdder_433_io_ci = FullAdder_171_io_s; // @[wallace.scala 71:19]
  assign FullAdder_434_io_a = FullAdder_172_io_s; // @[wallace.scala 69:18]
  assign FullAdder_434_io_b = FullAdder_173_io_s; // @[wallace.scala 70:18]
  assign FullAdder_434_io_ci = FullAdder_174_io_co; // @[wallace.scala 71:19]
  assign FullAdder_435_io_a = FullAdder_175_io_co; // @[wallace.scala 69:18]
  assign FullAdder_435_io_b = FullAdder_176_io_co; // @[wallace.scala 70:18]
  assign FullAdder_435_io_ci = FullAdder_177_io_co; // @[wallace.scala 71:19]
  assign FullAdder_436_io_a = FullAdder_178_io_co; // @[wallace.scala 69:18]
  assign FullAdder_436_io_b = FullAdder_179_io_co; // @[wallace.scala 70:18]
  assign FullAdder_436_io_ci = FullAdder_180_io_co; // @[wallace.scala 71:19]
  assign FullAdder_437_io_a = FullAdder_181_io_co; // @[wallace.scala 69:18]
  assign FullAdder_437_io_b = FullAdder_182_io_co; // @[wallace.scala 70:18]
  assign FullAdder_437_io_ci = FullAdder_183_io_co; // @[wallace.scala 71:19]
  assign FullAdder_438_io_a = FullAdder_174_io_s; // @[wallace.scala 69:18]
  assign FullAdder_438_io_b = FullAdder_175_io_s; // @[wallace.scala 70:18]
  assign FullAdder_438_io_ci = FullAdder_176_io_s; // @[wallace.scala 71:19]
  assign FullAdder_439_io_a = FullAdder_177_io_s; // @[wallace.scala 69:18]
  assign FullAdder_439_io_b = FullAdder_178_io_s; // @[wallace.scala 70:18]
  assign FullAdder_439_io_ci = FullAdder_179_io_s; // @[wallace.scala 71:19]
  assign FullAdder_440_io_a = FullAdder_180_io_s; // @[wallace.scala 69:18]
  assign FullAdder_440_io_b = FullAdder_181_io_s; // @[wallace.scala 70:18]
  assign FullAdder_440_io_ci = FullAdder_182_io_s; // @[wallace.scala 71:19]
  assign FullAdder_441_io_a = FullAdder_183_io_s; // @[wallace.scala 69:18]
  assign FullAdder_441_io_b = FullAdder_184_io_co; // @[wallace.scala 70:18]
  assign FullAdder_441_io_ci = FullAdder_185_io_co; // @[wallace.scala 71:19]
  assign FullAdder_442_io_a = FullAdder_186_io_co; // @[wallace.scala 69:18]
  assign FullAdder_442_io_b = FullAdder_187_io_co; // @[wallace.scala 70:18]
  assign FullAdder_442_io_ci = FullAdder_188_io_co; // @[wallace.scala 71:19]
  assign FullAdder_443_io_a = FullAdder_189_io_co; // @[wallace.scala 69:18]
  assign FullAdder_443_io_b = FullAdder_190_io_co; // @[wallace.scala 70:18]
  assign FullAdder_443_io_ci = FullAdder_191_io_co; // @[wallace.scala 71:19]
  assign FullAdder_444_io_a = FullAdder_184_io_s; // @[wallace.scala 69:18]
  assign FullAdder_444_io_b = FullAdder_185_io_s; // @[wallace.scala 70:18]
  assign FullAdder_444_io_ci = FullAdder_186_io_s; // @[wallace.scala 71:19]
  assign FullAdder_445_io_a = FullAdder_187_io_s; // @[wallace.scala 69:18]
  assign FullAdder_445_io_b = FullAdder_188_io_s; // @[wallace.scala 70:18]
  assign FullAdder_445_io_ci = FullAdder_189_io_s; // @[wallace.scala 71:19]
  assign FullAdder_446_io_a = FullAdder_190_io_s; // @[wallace.scala 69:18]
  assign FullAdder_446_io_b = FullAdder_191_io_s; // @[wallace.scala 70:18]
  assign FullAdder_446_io_ci = FullAdder_192_io_s; // @[wallace.scala 71:19]
  assign FullAdder_447_io_a = HalfAdder_8_io_s; // @[wallace.scala 69:18]
  assign FullAdder_447_io_b = FullAdder_193_io_co; // @[wallace.scala 70:18]
  assign FullAdder_447_io_ci = FullAdder_194_io_co; // @[wallace.scala 71:19]
  assign FullAdder_448_io_a = FullAdder_195_io_co; // @[wallace.scala 69:18]
  assign FullAdder_448_io_b = FullAdder_196_io_co; // @[wallace.scala 70:18]
  assign FullAdder_448_io_ci = FullAdder_197_io_co; // @[wallace.scala 71:19]
  assign FullAdder_449_io_a = FullAdder_198_io_co; // @[wallace.scala 69:18]
  assign FullAdder_449_io_b = FullAdder_199_io_co; // @[wallace.scala 70:18]
  assign FullAdder_449_io_ci = FullAdder_200_io_co; // @[wallace.scala 71:19]
  assign FullAdder_450_io_a = io_pp_27[0]; // @[wallace.scala 69:18]
  assign FullAdder_450_io_b = FullAdder_193_io_s; // @[wallace.scala 70:18]
  assign FullAdder_450_io_ci = FullAdder_194_io_s; // @[wallace.scala 71:19]
  assign FullAdder_451_io_a = FullAdder_195_io_s; // @[wallace.scala 69:18]
  assign FullAdder_451_io_b = FullAdder_196_io_s; // @[wallace.scala 70:18]
  assign FullAdder_451_io_ci = FullAdder_197_io_s; // @[wallace.scala 71:19]
  assign FullAdder_452_io_a = FullAdder_198_io_s; // @[wallace.scala 69:18]
  assign FullAdder_452_io_b = FullAdder_199_io_s; // @[wallace.scala 70:18]
  assign FullAdder_452_io_ci = FullAdder_200_io_s; // @[wallace.scala 71:19]
  assign FullAdder_453_io_a = FullAdder_201_io_s; // @[wallace.scala 69:18]
  assign FullAdder_453_io_b = FullAdder_202_io_co; // @[wallace.scala 70:18]
  assign FullAdder_453_io_ci = FullAdder_203_io_co; // @[wallace.scala 71:19]
  assign FullAdder_454_io_a = FullAdder_204_io_co; // @[wallace.scala 69:18]
  assign FullAdder_454_io_b = FullAdder_205_io_co; // @[wallace.scala 70:18]
  assign FullAdder_454_io_ci = FullAdder_206_io_co; // @[wallace.scala 71:19]
  assign FullAdder_455_io_a = FullAdder_207_io_co; // @[wallace.scala 69:18]
  assign FullAdder_455_io_b = FullAdder_208_io_co; // @[wallace.scala 70:18]
  assign FullAdder_455_io_ci = FullAdder_209_io_co; // @[wallace.scala 71:19]
  assign FullAdder_456_io_a = FullAdder_202_io_s; // @[wallace.scala 69:18]
  assign FullAdder_456_io_b = FullAdder_203_io_s; // @[wallace.scala 70:18]
  assign FullAdder_456_io_ci = FullAdder_204_io_s; // @[wallace.scala 71:19]
  assign FullAdder_457_io_a = FullAdder_205_io_s; // @[wallace.scala 69:18]
  assign FullAdder_457_io_b = FullAdder_206_io_s; // @[wallace.scala 70:18]
  assign FullAdder_457_io_ci = FullAdder_207_io_s; // @[wallace.scala 71:19]
  assign FullAdder_458_io_a = FullAdder_208_io_s; // @[wallace.scala 69:18]
  assign FullAdder_458_io_b = FullAdder_209_io_s; // @[wallace.scala 70:18]
  assign FullAdder_458_io_ci = FullAdder_210_io_s; // @[wallace.scala 71:19]
  assign FullAdder_459_io_a = FullAdder_211_io_co; // @[wallace.scala 69:18]
  assign FullAdder_459_io_b = FullAdder_212_io_co; // @[wallace.scala 70:18]
  assign FullAdder_459_io_ci = FullAdder_213_io_co; // @[wallace.scala 71:19]
  assign FullAdder_460_io_a = FullAdder_214_io_co; // @[wallace.scala 69:18]
  assign FullAdder_460_io_b = FullAdder_215_io_co; // @[wallace.scala 70:18]
  assign FullAdder_460_io_ci = FullAdder_216_io_co; // @[wallace.scala 71:19]
  assign FullAdder_461_io_a = FullAdder_217_io_co; // @[wallace.scala 69:18]
  assign FullAdder_461_io_b = FullAdder_218_io_co; // @[wallace.scala 70:18]
  assign FullAdder_461_io_ci = HalfAdder_9_io_co; // @[wallace.scala 71:19]
  assign FullAdder_462_io_a = FullAdder_211_io_s; // @[wallace.scala 69:18]
  assign FullAdder_462_io_b = FullAdder_212_io_s; // @[wallace.scala 70:18]
  assign FullAdder_462_io_ci = FullAdder_213_io_s; // @[wallace.scala 71:19]
  assign FullAdder_463_io_a = FullAdder_214_io_s; // @[wallace.scala 69:18]
  assign FullAdder_463_io_b = FullAdder_215_io_s; // @[wallace.scala 70:18]
  assign FullAdder_463_io_ci = FullAdder_216_io_s; // @[wallace.scala 71:19]
  assign FullAdder_464_io_a = FullAdder_217_io_s; // @[wallace.scala 69:18]
  assign FullAdder_464_io_b = FullAdder_218_io_s; // @[wallace.scala 70:18]
  assign FullAdder_464_io_ci = HalfAdder_9_io_s; // @[wallace.scala 71:19]
  assign FullAdder_465_io_a = FullAdder_219_io_co; // @[wallace.scala 69:18]
  assign FullAdder_465_io_b = FullAdder_220_io_co; // @[wallace.scala 70:18]
  assign FullAdder_465_io_ci = FullAdder_221_io_co; // @[wallace.scala 71:19]
  assign FullAdder_466_io_a = FullAdder_222_io_co; // @[wallace.scala 69:18]
  assign FullAdder_466_io_b = FullAdder_223_io_co; // @[wallace.scala 70:18]
  assign FullAdder_466_io_ci = FullAdder_224_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_25_io_a = FullAdder_225_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_25_io_b = FullAdder_226_io_co; // @[wallace.scala 60:18]
  assign FullAdder_467_io_a = io_pp_24[0]; // @[wallace.scala 69:18]
  assign FullAdder_467_io_b = FullAdder_219_io_s; // @[wallace.scala 70:18]
  assign FullAdder_467_io_ci = FullAdder_220_io_s; // @[wallace.scala 71:19]
  assign FullAdder_468_io_a = FullAdder_221_io_s; // @[wallace.scala 69:18]
  assign FullAdder_468_io_b = FullAdder_222_io_s; // @[wallace.scala 70:18]
  assign FullAdder_468_io_ci = FullAdder_223_io_s; // @[wallace.scala 71:19]
  assign FullAdder_469_io_a = FullAdder_224_io_s; // @[wallace.scala 69:18]
  assign FullAdder_469_io_b = FullAdder_225_io_s; // @[wallace.scala 70:18]
  assign FullAdder_469_io_ci = FullAdder_226_io_s; // @[wallace.scala 71:19]
  assign FullAdder_470_io_a = FullAdder_227_io_co; // @[wallace.scala 69:18]
  assign FullAdder_470_io_b = FullAdder_228_io_co; // @[wallace.scala 70:18]
  assign FullAdder_470_io_ci = FullAdder_229_io_co; // @[wallace.scala 71:19]
  assign FullAdder_471_io_a = FullAdder_230_io_co; // @[wallace.scala 69:18]
  assign FullAdder_471_io_b = FullAdder_231_io_co; // @[wallace.scala 70:18]
  assign FullAdder_471_io_ci = FullAdder_232_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_26_io_a = FullAdder_233_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_26_io_b = FullAdder_234_io_co; // @[wallace.scala 60:18]
  assign FullAdder_472_io_a = FullAdder_227_io_s; // @[wallace.scala 69:18]
  assign FullAdder_472_io_b = FullAdder_228_io_s; // @[wallace.scala 70:18]
  assign FullAdder_472_io_ci = FullAdder_229_io_s; // @[wallace.scala 71:19]
  assign FullAdder_473_io_a = FullAdder_230_io_s; // @[wallace.scala 69:18]
  assign FullAdder_473_io_b = FullAdder_231_io_s; // @[wallace.scala 70:18]
  assign FullAdder_473_io_ci = FullAdder_232_io_s; // @[wallace.scala 71:19]
  assign FullAdder_474_io_a = FullAdder_233_io_s; // @[wallace.scala 69:18]
  assign FullAdder_474_io_b = FullAdder_234_io_s; // @[wallace.scala 70:18]
  assign FullAdder_474_io_ci = FullAdder_235_io_co; // @[wallace.scala 71:19]
  assign FullAdder_475_io_a = FullAdder_236_io_co; // @[wallace.scala 69:18]
  assign FullAdder_475_io_b = FullAdder_237_io_co; // @[wallace.scala 70:18]
  assign FullAdder_475_io_ci = FullAdder_238_io_co; // @[wallace.scala 71:19]
  assign FullAdder_476_io_a = FullAdder_239_io_co; // @[wallace.scala 69:18]
  assign FullAdder_476_io_b = FullAdder_240_io_co; // @[wallace.scala 70:18]
  assign FullAdder_476_io_ci = FullAdder_241_io_co; // @[wallace.scala 71:19]
  assign FullAdder_477_io_a = io_pp_21[1]; // @[wallace.scala 69:18]
  assign FullAdder_477_io_b = io_pp_22[0]; // @[wallace.scala 70:18]
  assign FullAdder_477_io_ci = FullAdder_235_io_s; // @[wallace.scala 71:19]
  assign FullAdder_478_io_a = FullAdder_236_io_s; // @[wallace.scala 69:18]
  assign FullAdder_478_io_b = FullAdder_237_io_s; // @[wallace.scala 70:18]
  assign FullAdder_478_io_ci = FullAdder_238_io_s; // @[wallace.scala 71:19]
  assign FullAdder_479_io_a = FullAdder_239_io_s; // @[wallace.scala 69:18]
  assign FullAdder_479_io_b = FullAdder_240_io_s; // @[wallace.scala 70:18]
  assign FullAdder_479_io_ci = FullAdder_241_io_s; // @[wallace.scala 71:19]
  assign FullAdder_480_io_a = FullAdder_242_io_co; // @[wallace.scala 69:18]
  assign FullAdder_480_io_b = FullAdder_243_io_co; // @[wallace.scala 70:18]
  assign FullAdder_480_io_ci = FullAdder_244_io_co; // @[wallace.scala 71:19]
  assign FullAdder_481_io_a = FullAdder_245_io_co; // @[wallace.scala 69:18]
  assign FullAdder_481_io_b = FullAdder_246_io_co; // @[wallace.scala 70:18]
  assign FullAdder_481_io_ci = FullAdder_247_io_co; // @[wallace.scala 71:19]
  assign FullAdder_482_io_a = io_pp_21[0]; // @[wallace.scala 69:18]
  assign FullAdder_482_io_b = FullAdder_242_io_s; // @[wallace.scala 70:18]
  assign FullAdder_482_io_ci = FullAdder_243_io_s; // @[wallace.scala 71:19]
  assign FullAdder_483_io_a = FullAdder_244_io_s; // @[wallace.scala 69:18]
  assign FullAdder_483_io_b = FullAdder_245_io_s; // @[wallace.scala 70:18]
  assign FullAdder_483_io_ci = FullAdder_246_io_s; // @[wallace.scala 71:19]
  assign FullAdder_484_io_a = FullAdder_247_io_s; // @[wallace.scala 69:18]
  assign FullAdder_484_io_b = FullAdder_248_io_s; // @[wallace.scala 70:18]
  assign FullAdder_484_io_ci = FullAdder_249_io_co; // @[wallace.scala 71:19]
  assign FullAdder_485_io_a = FullAdder_250_io_co; // @[wallace.scala 69:18]
  assign FullAdder_485_io_b = FullAdder_251_io_co; // @[wallace.scala 70:18]
  assign FullAdder_485_io_ci = FullAdder_252_io_co; // @[wallace.scala 71:19]
  assign FullAdder_486_io_a = FullAdder_253_io_co; // @[wallace.scala 69:18]
  assign FullAdder_486_io_b = FullAdder_254_io_co; // @[wallace.scala 70:18]
  assign FullAdder_486_io_ci = FullAdder_255_io_co; // @[wallace.scala 71:19]
  assign FullAdder_487_io_a = FullAdder_249_io_s; // @[wallace.scala 69:18]
  assign FullAdder_487_io_b = FullAdder_250_io_s; // @[wallace.scala 70:18]
  assign FullAdder_487_io_ci = FullAdder_251_io_s; // @[wallace.scala 71:19]
  assign FullAdder_488_io_a = FullAdder_252_io_s; // @[wallace.scala 69:18]
  assign FullAdder_488_io_b = FullAdder_253_io_s; // @[wallace.scala 70:18]
  assign FullAdder_488_io_ci = FullAdder_254_io_s; // @[wallace.scala 71:19]
  assign FullAdder_489_io_a = FullAdder_255_io_s; // @[wallace.scala 69:18]
  assign FullAdder_489_io_b = FullAdder_256_io_co; // @[wallace.scala 70:18]
  assign FullAdder_489_io_ci = FullAdder_257_io_co; // @[wallace.scala 71:19]
  assign FullAdder_490_io_a = FullAdder_258_io_co; // @[wallace.scala 69:18]
  assign FullAdder_490_io_b = FullAdder_259_io_co; // @[wallace.scala 70:18]
  assign FullAdder_490_io_ci = FullAdder_260_io_co; // @[wallace.scala 71:19]
  assign FullAdder_491_io_a = io_pp_18[1]; // @[wallace.scala 69:18]
  assign FullAdder_491_io_b = io_pp_19[0]; // @[wallace.scala 70:18]
  assign FullAdder_491_io_ci = FullAdder_256_io_s; // @[wallace.scala 71:19]
  assign FullAdder_492_io_a = FullAdder_257_io_s; // @[wallace.scala 69:18]
  assign FullAdder_492_io_b = FullAdder_258_io_s; // @[wallace.scala 70:18]
  assign FullAdder_492_io_ci = FullAdder_259_io_s; // @[wallace.scala 71:19]
  assign FullAdder_493_io_a = FullAdder_260_io_s; // @[wallace.scala 69:18]
  assign FullAdder_493_io_b = FullAdder_261_io_s; // @[wallace.scala 70:18]
  assign FullAdder_493_io_ci = FullAdder_262_io_co; // @[wallace.scala 71:19]
  assign FullAdder_494_io_a = FullAdder_263_io_co; // @[wallace.scala 69:18]
  assign FullAdder_494_io_b = FullAdder_264_io_co; // @[wallace.scala 70:18]
  assign FullAdder_494_io_ci = FullAdder_265_io_co; // @[wallace.scala 71:19]
  assign FullAdder_495_io_a = io_pp_18[0]; // @[wallace.scala 69:18]
  assign FullAdder_495_io_b = FullAdder_262_io_s; // @[wallace.scala 70:18]
  assign FullAdder_495_io_ci = FullAdder_263_io_s; // @[wallace.scala 71:19]
  assign FullAdder_496_io_a = FullAdder_264_io_s; // @[wallace.scala 69:18]
  assign FullAdder_496_io_b = FullAdder_265_io_s; // @[wallace.scala 70:18]
  assign FullAdder_496_io_ci = FullAdder_266_io_s; // @[wallace.scala 71:19]
  assign FullAdder_497_io_a = FullAdder_267_io_s; // @[wallace.scala 69:18]
  assign FullAdder_497_io_b = FullAdder_268_io_co; // @[wallace.scala 70:18]
  assign FullAdder_497_io_ci = FullAdder_269_io_co; // @[wallace.scala 71:19]
  assign FullAdder_498_io_a = FullAdder_270_io_co; // @[wallace.scala 69:18]
  assign FullAdder_498_io_b = FullAdder_271_io_co; // @[wallace.scala 70:18]
  assign FullAdder_498_io_ci = FullAdder_272_io_co; // @[wallace.scala 71:19]
  assign FullAdder_499_io_a = FullAdder_268_io_s; // @[wallace.scala 69:18]
  assign FullAdder_499_io_b = FullAdder_269_io_s; // @[wallace.scala 70:18]
  assign FullAdder_499_io_ci = FullAdder_270_io_s; // @[wallace.scala 71:19]
  assign FullAdder_500_io_a = FullAdder_271_io_s; // @[wallace.scala 69:18]
  assign FullAdder_500_io_b = FullAdder_272_io_s; // @[wallace.scala 70:18]
  assign FullAdder_500_io_ci = FullAdder_273_io_s; // @[wallace.scala 71:19]
  assign FullAdder_501_io_a = FullAdder_274_io_co; // @[wallace.scala 69:18]
  assign FullAdder_501_io_b = FullAdder_275_io_co; // @[wallace.scala 70:18]
  assign FullAdder_501_io_ci = FullAdder_276_io_co; // @[wallace.scala 71:19]
  assign FullAdder_502_io_a = FullAdder_277_io_co; // @[wallace.scala 69:18]
  assign FullAdder_502_io_b = FullAdder_278_io_co; // @[wallace.scala 70:18]
  assign FullAdder_502_io_ci = HalfAdder_10_io_co; // @[wallace.scala 71:19]
  assign FullAdder_503_io_a = FullAdder_274_io_s; // @[wallace.scala 69:18]
  assign FullAdder_503_io_b = FullAdder_275_io_s; // @[wallace.scala 70:18]
  assign FullAdder_503_io_ci = FullAdder_276_io_s; // @[wallace.scala 71:19]
  assign FullAdder_504_io_a = FullAdder_277_io_s; // @[wallace.scala 69:18]
  assign FullAdder_504_io_b = FullAdder_278_io_s; // @[wallace.scala 70:18]
  assign FullAdder_504_io_ci = HalfAdder_10_io_s; // @[wallace.scala 71:19]
  assign FullAdder_505_io_a = FullAdder_279_io_co; // @[wallace.scala 69:18]
  assign FullAdder_505_io_b = FullAdder_280_io_co; // @[wallace.scala 70:18]
  assign FullAdder_505_io_ci = FullAdder_281_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_27_io_a = FullAdder_282_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_27_io_b = FullAdder_283_io_co; // @[wallace.scala 60:18]
  assign FullAdder_506_io_a = io_pp_15[0]; // @[wallace.scala 69:18]
  assign FullAdder_506_io_b = FullAdder_279_io_s; // @[wallace.scala 70:18]
  assign FullAdder_506_io_ci = FullAdder_280_io_s; // @[wallace.scala 71:19]
  assign FullAdder_507_io_a = FullAdder_281_io_s; // @[wallace.scala 69:18]
  assign FullAdder_507_io_b = FullAdder_282_io_s; // @[wallace.scala 70:18]
  assign FullAdder_507_io_ci = FullAdder_283_io_s; // @[wallace.scala 71:19]
  assign FullAdder_508_io_a = FullAdder_284_io_co; // @[wallace.scala 69:18]
  assign FullAdder_508_io_b = FullAdder_285_io_co; // @[wallace.scala 70:18]
  assign FullAdder_508_io_ci = FullAdder_286_io_co; // @[wallace.scala 71:19]
  assign FullAdder_509_io_a = FullAdder_284_io_s; // @[wallace.scala 69:18]
  assign FullAdder_509_io_b = FullAdder_285_io_s; // @[wallace.scala 70:18]
  assign FullAdder_509_io_ci = FullAdder_286_io_s; // @[wallace.scala 71:19]
  assign FullAdder_510_io_a = FullAdder_287_io_s; // @[wallace.scala 69:18]
  assign FullAdder_510_io_b = FullAdder_288_io_s; // @[wallace.scala 70:18]
  assign FullAdder_510_io_ci = FullAdder_289_io_co; // @[wallace.scala 71:19]
  assign FullAdder_511_io_a = FullAdder_290_io_co; // @[wallace.scala 69:18]
  assign FullAdder_511_io_b = FullAdder_291_io_co; // @[wallace.scala 70:18]
  assign FullAdder_511_io_ci = FullAdder_292_io_co; // @[wallace.scala 71:19]
  assign FullAdder_512_io_a = io_pp_12[1]; // @[wallace.scala 69:18]
  assign FullAdder_512_io_b = io_pp_13[0]; // @[wallace.scala 70:18]
  assign FullAdder_512_io_ci = FullAdder_289_io_s; // @[wallace.scala 71:19]
  assign FullAdder_513_io_a = FullAdder_290_io_s; // @[wallace.scala 69:18]
  assign FullAdder_513_io_b = FullAdder_291_io_s; // @[wallace.scala 70:18]
  assign FullAdder_513_io_ci = FullAdder_292_io_s; // @[wallace.scala 71:19]
  assign FullAdder_514_io_a = FullAdder_293_io_co; // @[wallace.scala 69:18]
  assign FullAdder_514_io_b = FullAdder_294_io_co; // @[wallace.scala 70:18]
  assign FullAdder_514_io_ci = FullAdder_295_io_co; // @[wallace.scala 71:19]
  assign FullAdder_515_io_a = io_pp_12[0]; // @[wallace.scala 69:18]
  assign FullAdder_515_io_b = FullAdder_293_io_s; // @[wallace.scala 70:18]
  assign FullAdder_515_io_ci = FullAdder_294_io_s; // @[wallace.scala 71:19]
  assign FullAdder_516_io_a = FullAdder_295_io_s; // @[wallace.scala 69:18]
  assign FullAdder_516_io_b = FullAdder_296_io_s; // @[wallace.scala 70:18]
  assign FullAdder_516_io_ci = FullAdder_297_io_co; // @[wallace.scala 71:19]
  assign FullAdder_517_io_a = FullAdder_298_io_co; // @[wallace.scala 69:18]
  assign FullAdder_517_io_b = FullAdder_299_io_co; // @[wallace.scala 70:18]
  assign FullAdder_517_io_ci = FullAdder_300_io_co; // @[wallace.scala 71:19]
  assign FullAdder_518_io_a = FullAdder_297_io_s; // @[wallace.scala 69:18]
  assign FullAdder_518_io_b = FullAdder_298_io_s; // @[wallace.scala 70:18]
  assign FullAdder_518_io_ci = FullAdder_299_io_s; // @[wallace.scala 71:19]
  assign FullAdder_519_io_a = FullAdder_300_io_s; // @[wallace.scala 69:18]
  assign FullAdder_519_io_b = FullAdder_301_io_co; // @[wallace.scala 70:18]
  assign FullAdder_519_io_ci = FullAdder_302_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_28_io_a = FullAdder_303_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_28_io_b = HalfAdder_11_io_co; // @[wallace.scala 60:18]
  assign FullAdder_520_io_a = FullAdder_301_io_s; // @[wallace.scala 69:18]
  assign FullAdder_520_io_b = FullAdder_302_io_s; // @[wallace.scala 70:18]
  assign FullAdder_520_io_ci = FullAdder_303_io_s; // @[wallace.scala 71:19]
  assign FullAdder_521_io_a = HalfAdder_11_io_s; // @[wallace.scala 69:18]
  assign FullAdder_521_io_b = FullAdder_304_io_co; // @[wallace.scala 70:18]
  assign FullAdder_521_io_ci = FullAdder_305_io_co; // @[wallace.scala 71:19]
  assign FullAdder_522_io_a = io_pp_9[0]; // @[wallace.scala 69:18]
  assign FullAdder_522_io_b = FullAdder_304_io_s; // @[wallace.scala 70:18]
  assign FullAdder_522_io_ci = FullAdder_305_io_s; // @[wallace.scala 71:19]
  assign FullAdder_523_io_a = FullAdder_306_io_s; // @[wallace.scala 69:18]
  assign FullAdder_523_io_b = FullAdder_307_io_co; // @[wallace.scala 70:18]
  assign FullAdder_523_io_ci = FullAdder_308_io_co; // @[wallace.scala 71:19]
  assign FullAdder_524_io_a = FullAdder_307_io_s; // @[wallace.scala 69:18]
  assign FullAdder_524_io_b = FullAdder_308_io_s; // @[wallace.scala 70:18]
  assign FullAdder_524_io_ci = FullAdder_309_io_s; // @[wallace.scala 71:19]
  assign FullAdder_525_io_a = FullAdder_310_io_co; // @[wallace.scala 69:18]
  assign FullAdder_525_io_b = FullAdder_311_io_co; // @[wallace.scala 70:18]
  assign FullAdder_525_io_ci = HalfAdder_12_io_co; // @[wallace.scala 71:19]
  assign FullAdder_526_io_a = FullAdder_310_io_s; // @[wallace.scala 69:18]
  assign FullAdder_526_io_b = FullAdder_311_io_s; // @[wallace.scala 70:18]
  assign FullAdder_526_io_ci = HalfAdder_12_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_29_io_a = FullAdder_312_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_29_io_b = FullAdder_313_io_co; // @[wallace.scala 60:18]
  assign FullAdder_527_io_a = io_pp_6[0]; // @[wallace.scala 69:18]
  assign FullAdder_527_io_b = FullAdder_312_io_s; // @[wallace.scala 70:18]
  assign FullAdder_527_io_ci = FullAdder_313_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_30_io_a = FullAdder_314_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_30_io_b = FullAdder_315_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_31_io_a = FullAdder_314_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_31_io_b = FullAdder_315_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_32_io_a = FullAdder_316_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_32_io_b = HalfAdder_13_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_33_io_a = FullAdder_316_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_33_io_b = HalfAdder_13_io_s; // @[wallace.scala 60:18]
  assign FullAdder_528_io_a = io_pp_3[0]; // @[wallace.scala 69:18]
  assign FullAdder_528_io_b = FullAdder_317_io_s; // @[wallace.scala 70:18]
  assign FullAdder_528_io_ci = FullAdder_318_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_34_io_a = HalfAdder_14_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_34_io_b = HalfAdder_15_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_35_io_a = HalfAdder_15_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_35_io_b = HalfAdder_16_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_36_io_a = FullAdder_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_36_io_b = HalfAdder_16_io_s; // @[wallace.scala 60:18]
  assign FullAdder_529_io_a = HalfAdder_2_io_co; // @[wallace.scala 69:18]
  assign FullAdder_529_io_b = FullAdder_319_io_s; // @[wallace.scala 70:18]
  assign FullAdder_529_io_ci = FullAdder_320_io_co; // @[wallace.scala 71:19]
  assign FullAdder_530_io_a = FullAdder_3_io_co; // @[wallace.scala 69:18]
  assign FullAdder_530_io_b = FullAdder_320_io_s; // @[wallace.scala 70:18]
  assign FullAdder_530_io_ci = FullAdder_321_io_co; // @[wallace.scala 71:19]
  assign FullAdder_531_io_a = FullAdder_5_io_co; // @[wallace.scala 69:18]
  assign FullAdder_531_io_b = FullAdder_321_io_s; // @[wallace.scala 70:18]
  assign FullAdder_531_io_ci = FullAdder_322_io_co; // @[wallace.scala 71:19]
  assign FullAdder_532_io_a = FullAdder_322_io_s; // @[wallace.scala 69:18]
  assign FullAdder_532_io_b = HalfAdder_17_io_s; // @[wallace.scala 70:18]
  assign FullAdder_532_io_ci = FullAdder_323_io_co; // @[wallace.scala 71:19]
  assign FullAdder_533_io_a = FullAdder_10_io_co; // @[wallace.scala 69:18]
  assign FullAdder_533_io_b = FullAdder_323_io_s; // @[wallace.scala 70:18]
  assign FullAdder_533_io_ci = FullAdder_324_io_s; // @[wallace.scala 71:19]
  assign FullAdder_534_io_a = FullAdder_325_io_s; // @[wallace.scala 69:18]
  assign FullAdder_534_io_b = FullAdder_326_io_s; // @[wallace.scala 70:18]
  assign FullAdder_534_io_ci = FullAdder_327_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_37_io_a = FullAdder_328_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_37_io_b = HalfAdder_18_io_co; // @[wallace.scala 60:18]
  assign FullAdder_535_io_a = FullAdder_327_io_s; // @[wallace.scala 69:18]
  assign FullAdder_535_io_b = FullAdder_328_io_s; // @[wallace.scala 70:18]
  assign FullAdder_535_io_ci = HalfAdder_18_io_s; // @[wallace.scala 71:19]
  assign FullAdder_536_io_a = FullAdder_329_io_co; // @[wallace.scala 69:18]
  assign FullAdder_536_io_b = FullAdder_330_io_co; // @[wallace.scala 70:18]
  assign FullAdder_536_io_ci = HalfAdder_19_io_co; // @[wallace.scala 71:19]
  assign FullAdder_537_io_a = FullAdder_329_io_s; // @[wallace.scala 69:18]
  assign FullAdder_537_io_b = FullAdder_330_io_s; // @[wallace.scala 70:18]
  assign FullAdder_537_io_ci = HalfAdder_19_io_s; // @[wallace.scala 71:19]
  assign FullAdder_538_io_a = FullAdder_331_io_co; // @[wallace.scala 69:18]
  assign FullAdder_538_io_b = FullAdder_332_io_co; // @[wallace.scala 70:18]
  assign FullAdder_538_io_ci = HalfAdder_20_io_co; // @[wallace.scala 71:19]
  assign FullAdder_539_io_a = FullAdder_331_io_s; // @[wallace.scala 69:18]
  assign FullAdder_539_io_b = FullAdder_332_io_s; // @[wallace.scala 70:18]
  assign FullAdder_539_io_ci = HalfAdder_20_io_s; // @[wallace.scala 71:19]
  assign FullAdder_540_io_a = FullAdder_333_io_co; // @[wallace.scala 69:18]
  assign FullAdder_540_io_b = FullAdder_334_io_co; // @[wallace.scala 70:18]
  assign FullAdder_540_io_ci = FullAdder_335_io_co; // @[wallace.scala 71:19]
  assign FullAdder_541_io_a = HalfAdder_4_io_co; // @[wallace.scala 69:18]
  assign FullAdder_541_io_b = FullAdder_333_io_s; // @[wallace.scala 70:18]
  assign FullAdder_541_io_ci = FullAdder_334_io_s; // @[wallace.scala 71:19]
  assign FullAdder_542_io_a = FullAdder_335_io_s; // @[wallace.scala 69:18]
  assign FullAdder_542_io_b = FullAdder_336_io_co; // @[wallace.scala 70:18]
  assign FullAdder_542_io_ci = FullAdder_337_io_co; // @[wallace.scala 71:19]
  assign FullAdder_543_io_a = FullAdder_33_io_co; // @[wallace.scala 69:18]
  assign FullAdder_543_io_b = FullAdder_336_io_s; // @[wallace.scala 70:18]
  assign FullAdder_543_io_ci = FullAdder_337_io_s; // @[wallace.scala 71:19]
  assign FullAdder_544_io_a = FullAdder_338_io_s; // @[wallace.scala 69:18]
  assign FullAdder_544_io_b = FullAdder_339_io_co; // @[wallace.scala 70:18]
  assign FullAdder_544_io_ci = FullAdder_340_io_co; // @[wallace.scala 71:19]
  assign FullAdder_545_io_a = FullAdder_38_io_co; // @[wallace.scala 69:18]
  assign FullAdder_545_io_b = FullAdder_339_io_s; // @[wallace.scala 70:18]
  assign FullAdder_545_io_ci = FullAdder_340_io_s; // @[wallace.scala 71:19]
  assign FullAdder_546_io_a = FullAdder_341_io_s; // @[wallace.scala 69:18]
  assign FullAdder_546_io_b = FullAdder_342_io_co; // @[wallace.scala 70:18]
  assign FullAdder_546_io_ci = FullAdder_343_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_38_io_a = FullAdder_344_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_38_io_b = FullAdder_345_io_co; // @[wallace.scala 60:18]
  assign FullAdder_547_io_a = FullAdder_342_io_s; // @[wallace.scala 69:18]
  assign FullAdder_547_io_b = FullAdder_343_io_s; // @[wallace.scala 70:18]
  assign FullAdder_547_io_ci = FullAdder_344_io_s; // @[wallace.scala 71:19]
  assign FullAdder_548_io_a = FullAdder_345_io_s; // @[wallace.scala 69:18]
  assign FullAdder_548_io_b = FullAdder_346_io_co; // @[wallace.scala 70:18]
  assign FullAdder_548_io_ci = FullAdder_347_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_39_io_a = FullAdder_348_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_39_io_b = FullAdder_349_io_co; // @[wallace.scala 60:18]
  assign FullAdder_549_io_a = FullAdder_346_io_s; // @[wallace.scala 69:18]
  assign FullAdder_549_io_b = FullAdder_347_io_s; // @[wallace.scala 70:18]
  assign FullAdder_549_io_ci = FullAdder_348_io_s; // @[wallace.scala 71:19]
  assign FullAdder_550_io_a = FullAdder_349_io_s; // @[wallace.scala 69:18]
  assign FullAdder_550_io_b = FullAdder_350_io_co; // @[wallace.scala 70:18]
  assign FullAdder_550_io_ci = FullAdder_351_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_40_io_a = FullAdder_352_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_40_io_b = FullAdder_353_io_co; // @[wallace.scala 60:18]
  assign FullAdder_551_io_a = FullAdder_350_io_s; // @[wallace.scala 69:18]
  assign FullAdder_551_io_b = FullAdder_351_io_s; // @[wallace.scala 70:18]
  assign FullAdder_551_io_ci = FullAdder_352_io_s; // @[wallace.scala 71:19]
  assign FullAdder_552_io_a = FullAdder_353_io_s; // @[wallace.scala 69:18]
  assign FullAdder_552_io_b = FullAdder_354_io_co; // @[wallace.scala 70:18]
  assign FullAdder_552_io_ci = FullAdder_355_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_41_io_a = FullAdder_356_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_41_io_b = FullAdder_357_io_co; // @[wallace.scala 60:18]
  assign FullAdder_553_io_a = FullAdder_61_io_co; // @[wallace.scala 69:18]
  assign FullAdder_553_io_b = FullAdder_354_io_s; // @[wallace.scala 70:18]
  assign FullAdder_553_io_ci = FullAdder_355_io_s; // @[wallace.scala 71:19]
  assign FullAdder_554_io_a = FullAdder_356_io_s; // @[wallace.scala 69:18]
  assign FullAdder_554_io_b = FullAdder_357_io_s; // @[wallace.scala 70:18]
  assign FullAdder_554_io_ci = FullAdder_358_io_co; // @[wallace.scala 71:19]
  assign FullAdder_555_io_a = FullAdder_359_io_co; // @[wallace.scala 69:18]
  assign FullAdder_555_io_b = FullAdder_360_io_co; // @[wallace.scala 70:18]
  assign FullAdder_555_io_ci = FullAdder_361_io_co; // @[wallace.scala 71:19]
  assign FullAdder_556_io_a = FullAdder_358_io_s; // @[wallace.scala 69:18]
  assign FullAdder_556_io_b = FullAdder_359_io_s; // @[wallace.scala 70:18]
  assign FullAdder_556_io_ci = FullAdder_360_io_s; // @[wallace.scala 71:19]
  assign FullAdder_557_io_a = FullAdder_361_io_s; // @[wallace.scala 69:18]
  assign FullAdder_557_io_b = FullAdder_362_io_s; // @[wallace.scala 70:18]
  assign FullAdder_557_io_ci = FullAdder_363_io_co; // @[wallace.scala 71:19]
  assign FullAdder_558_io_a = FullAdder_364_io_co; // @[wallace.scala 69:18]
  assign FullAdder_558_io_b = FullAdder_365_io_co; // @[wallace.scala 70:18]
  assign FullAdder_558_io_ci = FullAdder_366_io_co; // @[wallace.scala 71:19]
  assign FullAdder_559_io_a = FullAdder_363_io_s; // @[wallace.scala 69:18]
  assign FullAdder_559_io_b = FullAdder_364_io_s; // @[wallace.scala 70:18]
  assign FullAdder_559_io_ci = FullAdder_365_io_s; // @[wallace.scala 71:19]
  assign FullAdder_560_io_a = FullAdder_366_io_s; // @[wallace.scala 69:18]
  assign FullAdder_560_io_b = HalfAdder_21_io_s; // @[wallace.scala 70:18]
  assign FullAdder_560_io_ci = FullAdder_367_io_co; // @[wallace.scala 71:19]
  assign FullAdder_561_io_a = FullAdder_368_io_co; // @[wallace.scala 69:18]
  assign FullAdder_561_io_b = FullAdder_369_io_co; // @[wallace.scala 70:18]
  assign FullAdder_561_io_ci = FullAdder_370_io_co; // @[wallace.scala 71:19]
  assign FullAdder_562_io_a = HalfAdder_6_io_co; // @[wallace.scala 69:18]
  assign FullAdder_562_io_b = FullAdder_367_io_s; // @[wallace.scala 70:18]
  assign FullAdder_562_io_ci = FullAdder_368_io_s; // @[wallace.scala 71:19]
  assign FullAdder_563_io_a = FullAdder_369_io_s; // @[wallace.scala 69:18]
  assign FullAdder_563_io_b = FullAdder_370_io_s; // @[wallace.scala 70:18]
  assign FullAdder_563_io_ci = FullAdder_371_io_s; // @[wallace.scala 71:19]
  assign FullAdder_564_io_a = FullAdder_372_io_co; // @[wallace.scala 69:18]
  assign FullAdder_564_io_b = FullAdder_373_io_co; // @[wallace.scala 70:18]
  assign FullAdder_564_io_ci = FullAdder_374_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_42_io_a = FullAdder_375_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_42_io_b = FullAdder_376_io_co; // @[wallace.scala 60:18]
  assign FullAdder_565_io_a = FullAdder_90_io_co; // @[wallace.scala 69:18]
  assign FullAdder_565_io_b = FullAdder_372_io_s; // @[wallace.scala 70:18]
  assign FullAdder_565_io_ci = FullAdder_373_io_s; // @[wallace.scala 71:19]
  assign FullAdder_566_io_a = FullAdder_374_io_s; // @[wallace.scala 69:18]
  assign FullAdder_566_io_b = FullAdder_375_io_s; // @[wallace.scala 70:18]
  assign FullAdder_566_io_ci = FullAdder_376_io_s; // @[wallace.scala 71:19]
  assign FullAdder_567_io_a = FullAdder_377_io_co; // @[wallace.scala 69:18]
  assign FullAdder_567_io_b = FullAdder_378_io_co; // @[wallace.scala 70:18]
  assign FullAdder_567_io_ci = FullAdder_379_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_43_io_a = FullAdder_380_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_43_io_b = FullAdder_381_io_co; // @[wallace.scala 60:18]
  assign FullAdder_568_io_a = FullAdder_98_io_co; // @[wallace.scala 69:18]
  assign FullAdder_568_io_b = FullAdder_377_io_s; // @[wallace.scala 70:18]
  assign FullAdder_568_io_ci = FullAdder_378_io_s; // @[wallace.scala 71:19]
  assign FullAdder_569_io_a = FullAdder_379_io_s; // @[wallace.scala 69:18]
  assign FullAdder_569_io_b = FullAdder_380_io_s; // @[wallace.scala 70:18]
  assign FullAdder_569_io_ci = FullAdder_381_io_s; // @[wallace.scala 71:19]
  assign FullAdder_570_io_a = FullAdder_382_io_co; // @[wallace.scala 69:18]
  assign FullAdder_570_io_b = FullAdder_383_io_co; // @[wallace.scala 70:18]
  assign FullAdder_570_io_ci = FullAdder_384_io_co; // @[wallace.scala 71:19]
  assign FullAdder_571_io_a = FullAdder_385_io_co; // @[wallace.scala 69:18]
  assign FullAdder_571_io_b = FullAdder_386_io_co; // @[wallace.scala 70:18]
  assign FullAdder_571_io_ci = HalfAdder_22_io_co; // @[wallace.scala 71:19]
  assign FullAdder_572_io_a = FullAdder_382_io_s; // @[wallace.scala 69:18]
  assign FullAdder_572_io_b = FullAdder_383_io_s; // @[wallace.scala 70:18]
  assign FullAdder_572_io_ci = FullAdder_384_io_s; // @[wallace.scala 71:19]
  assign FullAdder_573_io_a = FullAdder_385_io_s; // @[wallace.scala 69:18]
  assign FullAdder_573_io_b = FullAdder_386_io_s; // @[wallace.scala 70:18]
  assign FullAdder_573_io_ci = HalfAdder_22_io_s; // @[wallace.scala 71:19]
  assign FullAdder_574_io_a = FullAdder_387_io_co; // @[wallace.scala 69:18]
  assign FullAdder_574_io_b = FullAdder_388_io_co; // @[wallace.scala 70:18]
  assign FullAdder_574_io_ci = FullAdder_389_io_co; // @[wallace.scala 71:19]
  assign FullAdder_575_io_a = FullAdder_390_io_co; // @[wallace.scala 69:18]
  assign FullAdder_575_io_b = FullAdder_391_io_co; // @[wallace.scala 70:18]
  assign FullAdder_575_io_ci = FullAdder_392_io_co; // @[wallace.scala 71:19]
  assign FullAdder_576_io_a = FullAdder_115_io_co; // @[wallace.scala 69:18]
  assign FullAdder_576_io_b = FullAdder_387_io_s; // @[wallace.scala 70:18]
  assign FullAdder_576_io_ci = FullAdder_388_io_s; // @[wallace.scala 71:19]
  assign FullAdder_577_io_a = FullAdder_389_io_s; // @[wallace.scala 69:18]
  assign FullAdder_577_io_b = FullAdder_390_io_s; // @[wallace.scala 70:18]
  assign FullAdder_577_io_ci = FullAdder_391_io_s; // @[wallace.scala 71:19]
  assign FullAdder_578_io_a = FullAdder_392_io_s; // @[wallace.scala 69:18]
  assign FullAdder_578_io_b = FullAdder_393_io_co; // @[wallace.scala 70:18]
  assign FullAdder_578_io_ci = FullAdder_394_io_co; // @[wallace.scala 71:19]
  assign FullAdder_579_io_a = FullAdder_395_io_co; // @[wallace.scala 69:18]
  assign FullAdder_579_io_b = FullAdder_396_io_co; // @[wallace.scala 70:18]
  assign FullAdder_579_io_ci = FullAdder_397_io_co; // @[wallace.scala 71:19]
  assign FullAdder_580_io_a = FullAdder_393_io_s; // @[wallace.scala 69:18]
  assign FullAdder_580_io_b = FullAdder_394_io_s; // @[wallace.scala 70:18]
  assign FullAdder_580_io_ci = FullAdder_395_io_s; // @[wallace.scala 71:19]
  assign FullAdder_581_io_a = FullAdder_396_io_s; // @[wallace.scala 69:18]
  assign FullAdder_581_io_b = FullAdder_397_io_s; // @[wallace.scala 70:18]
  assign FullAdder_581_io_ci = FullAdder_398_io_s; // @[wallace.scala 71:19]
  assign FullAdder_582_io_a = FullAdder_399_io_co; // @[wallace.scala 69:18]
  assign FullAdder_582_io_b = FullAdder_400_io_co; // @[wallace.scala 70:18]
  assign FullAdder_582_io_ci = FullAdder_401_io_co; // @[wallace.scala 71:19]
  assign FullAdder_583_io_a = FullAdder_402_io_co; // @[wallace.scala 69:18]
  assign FullAdder_583_io_b = FullAdder_403_io_co; // @[wallace.scala 70:18]
  assign FullAdder_583_io_ci = FullAdder_404_io_co; // @[wallace.scala 71:19]
  assign FullAdder_584_io_a = FullAdder_399_io_s; // @[wallace.scala 69:18]
  assign FullAdder_584_io_b = FullAdder_400_io_s; // @[wallace.scala 70:18]
  assign FullAdder_584_io_ci = FullAdder_401_io_s; // @[wallace.scala 71:19]
  assign FullAdder_585_io_a = FullAdder_402_io_s; // @[wallace.scala 69:18]
  assign FullAdder_585_io_b = FullAdder_403_io_s; // @[wallace.scala 70:18]
  assign FullAdder_585_io_ci = FullAdder_404_io_s; // @[wallace.scala 71:19]
  assign FullAdder_586_io_a = HalfAdder_23_io_s; // @[wallace.scala 69:18]
  assign FullAdder_586_io_b = FullAdder_405_io_co; // @[wallace.scala 70:18]
  assign FullAdder_586_io_ci = FullAdder_406_io_co; // @[wallace.scala 71:19]
  assign FullAdder_587_io_a = FullAdder_407_io_co; // @[wallace.scala 69:18]
  assign FullAdder_587_io_b = FullAdder_408_io_co; // @[wallace.scala 70:18]
  assign FullAdder_587_io_ci = FullAdder_409_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_44_io_a = FullAdder_410_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_44_io_b = HalfAdder_24_io_co; // @[wallace.scala 60:18]
  assign FullAdder_588_io_a = FullAdder_405_io_s; // @[wallace.scala 69:18]
  assign FullAdder_588_io_b = FullAdder_406_io_s; // @[wallace.scala 70:18]
  assign FullAdder_588_io_ci = FullAdder_407_io_s; // @[wallace.scala 71:19]
  assign FullAdder_589_io_a = FullAdder_408_io_s; // @[wallace.scala 69:18]
  assign FullAdder_589_io_b = FullAdder_409_io_s; // @[wallace.scala 70:18]
  assign FullAdder_589_io_ci = FullAdder_410_io_s; // @[wallace.scala 71:19]
  assign FullAdder_590_io_a = HalfAdder_24_io_s; // @[wallace.scala 69:18]
  assign FullAdder_590_io_b = FullAdder_411_io_co; // @[wallace.scala 70:18]
  assign FullAdder_590_io_ci = FullAdder_412_io_co; // @[wallace.scala 71:19]
  assign FullAdder_591_io_a = FullAdder_413_io_co; // @[wallace.scala 69:18]
  assign FullAdder_591_io_b = FullAdder_414_io_co; // @[wallace.scala 70:18]
  assign FullAdder_591_io_ci = FullAdder_415_io_co; // @[wallace.scala 71:19]
  assign FullAdder_592_io_a = FullAdder_152_io_co; // @[wallace.scala 69:18]
  assign FullAdder_592_io_b = FullAdder_153_io_co; // @[wallace.scala 70:18]
  assign FullAdder_592_io_ci = FullAdder_411_io_s; // @[wallace.scala 71:19]
  assign FullAdder_593_io_a = FullAdder_412_io_s; // @[wallace.scala 69:18]
  assign FullAdder_593_io_b = FullAdder_413_io_s; // @[wallace.scala 70:18]
  assign FullAdder_593_io_ci = FullAdder_414_io_s; // @[wallace.scala 71:19]
  assign FullAdder_594_io_a = FullAdder_415_io_s; // @[wallace.scala 69:18]
  assign FullAdder_594_io_b = FullAdder_416_io_s; // @[wallace.scala 70:18]
  assign FullAdder_594_io_ci = FullAdder_417_io_co; // @[wallace.scala 71:19]
  assign FullAdder_595_io_a = FullAdder_418_io_co; // @[wallace.scala 69:18]
  assign FullAdder_595_io_b = FullAdder_419_io_co; // @[wallace.scala 70:18]
  assign FullAdder_595_io_ci = FullAdder_420_io_co; // @[wallace.scala 71:19]
  assign FullAdder_596_io_a = FullAdder_421_io_co; // @[wallace.scala 69:18]
  assign FullAdder_596_io_b = FullAdder_422_io_co; // @[wallace.scala 70:18]
  assign FullAdder_596_io_ci = FullAdder_423_io_co; // @[wallace.scala 71:19]
  assign FullAdder_597_io_a = FullAdder_417_io_s; // @[wallace.scala 69:18]
  assign FullAdder_597_io_b = FullAdder_418_io_s; // @[wallace.scala 70:18]
  assign FullAdder_597_io_ci = FullAdder_419_io_s; // @[wallace.scala 71:19]
  assign FullAdder_598_io_a = FullAdder_420_io_s; // @[wallace.scala 69:18]
  assign FullAdder_598_io_b = FullAdder_421_io_s; // @[wallace.scala 70:18]
  assign FullAdder_598_io_ci = FullAdder_422_io_s; // @[wallace.scala 71:19]
  assign FullAdder_599_io_a = FullAdder_423_io_s; // @[wallace.scala 69:18]
  assign FullAdder_599_io_b = FullAdder_424_io_co; // @[wallace.scala 70:18]
  assign FullAdder_599_io_ci = FullAdder_425_io_co; // @[wallace.scala 71:19]
  assign FullAdder_600_io_a = FullAdder_426_io_co; // @[wallace.scala 69:18]
  assign FullAdder_600_io_b = FullAdder_427_io_co; // @[wallace.scala 70:18]
  assign FullAdder_600_io_ci = FullAdder_428_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_45_io_a = FullAdder_429_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_45_io_b = FullAdder_430_io_co; // @[wallace.scala 60:18]
  assign FullAdder_601_io_a = FullAdder_173_io_co; // @[wallace.scala 69:18]
  assign FullAdder_601_io_b = FullAdder_424_io_s; // @[wallace.scala 70:18]
  assign FullAdder_601_io_ci = FullAdder_425_io_s; // @[wallace.scala 71:19]
  assign FullAdder_602_io_a = FullAdder_426_io_s; // @[wallace.scala 69:18]
  assign FullAdder_602_io_b = FullAdder_427_io_s; // @[wallace.scala 70:18]
  assign FullAdder_602_io_ci = FullAdder_428_io_s; // @[wallace.scala 71:19]
  assign FullAdder_603_io_a = FullAdder_429_io_s; // @[wallace.scala 69:18]
  assign FullAdder_603_io_b = FullAdder_430_io_s; // @[wallace.scala 70:18]
  assign FullAdder_603_io_ci = FullAdder_431_io_co; // @[wallace.scala 71:19]
  assign FullAdder_604_io_a = FullAdder_432_io_co; // @[wallace.scala 69:18]
  assign FullAdder_604_io_b = FullAdder_433_io_co; // @[wallace.scala 70:18]
  assign FullAdder_604_io_ci = FullAdder_434_io_co; // @[wallace.scala 71:19]
  assign FullAdder_605_io_a = FullAdder_435_io_co; // @[wallace.scala 69:18]
  assign FullAdder_605_io_b = FullAdder_436_io_co; // @[wallace.scala 70:18]
  assign FullAdder_605_io_ci = FullAdder_437_io_co; // @[wallace.scala 71:19]
  assign FullAdder_606_io_a = FullAdder_431_io_s; // @[wallace.scala 69:18]
  assign FullAdder_606_io_b = FullAdder_432_io_s; // @[wallace.scala 70:18]
  assign FullAdder_606_io_ci = FullAdder_433_io_s; // @[wallace.scala 71:19]
  assign FullAdder_607_io_a = FullAdder_434_io_s; // @[wallace.scala 69:18]
  assign FullAdder_607_io_b = FullAdder_435_io_s; // @[wallace.scala 70:18]
  assign FullAdder_607_io_ci = FullAdder_436_io_s; // @[wallace.scala 71:19]
  assign FullAdder_608_io_a = FullAdder_437_io_s; // @[wallace.scala 69:18]
  assign FullAdder_608_io_b = FullAdder_438_io_co; // @[wallace.scala 70:18]
  assign FullAdder_608_io_ci = FullAdder_439_io_co; // @[wallace.scala 71:19]
  assign FullAdder_609_io_a = FullAdder_440_io_co; // @[wallace.scala 69:18]
  assign FullAdder_609_io_b = FullAdder_441_io_co; // @[wallace.scala 70:18]
  assign FullAdder_609_io_ci = FullAdder_442_io_co; // @[wallace.scala 71:19]
  assign FullAdder_610_io_a = FullAdder_192_io_co; // @[wallace.scala 69:18]
  assign FullAdder_610_io_b = HalfAdder_8_io_co; // @[wallace.scala 70:18]
  assign FullAdder_610_io_ci = FullAdder_438_io_s; // @[wallace.scala 71:19]
  assign FullAdder_611_io_a = FullAdder_439_io_s; // @[wallace.scala 69:18]
  assign FullAdder_611_io_b = FullAdder_440_io_s; // @[wallace.scala 70:18]
  assign FullAdder_611_io_ci = FullAdder_441_io_s; // @[wallace.scala 71:19]
  assign FullAdder_612_io_a = FullAdder_442_io_s; // @[wallace.scala 69:18]
  assign FullAdder_612_io_b = FullAdder_443_io_s; // @[wallace.scala 70:18]
  assign FullAdder_612_io_ci = FullAdder_444_io_co; // @[wallace.scala 71:19]
  assign FullAdder_613_io_a = FullAdder_445_io_co; // @[wallace.scala 69:18]
  assign FullAdder_613_io_b = FullAdder_446_io_co; // @[wallace.scala 70:18]
  assign FullAdder_613_io_ci = FullAdder_447_io_co; // @[wallace.scala 71:19]
  assign FullAdder_614_io_a = FullAdder_201_io_co; // @[wallace.scala 69:18]
  assign FullAdder_614_io_b = FullAdder_444_io_s; // @[wallace.scala 70:18]
  assign FullAdder_614_io_ci = FullAdder_445_io_s; // @[wallace.scala 71:19]
  assign FullAdder_615_io_a = FullAdder_446_io_s; // @[wallace.scala 69:18]
  assign FullAdder_615_io_b = FullAdder_447_io_s; // @[wallace.scala 70:18]
  assign FullAdder_615_io_ci = FullAdder_448_io_s; // @[wallace.scala 71:19]
  assign FullAdder_616_io_a = FullAdder_449_io_s; // @[wallace.scala 69:18]
  assign FullAdder_616_io_b = FullAdder_450_io_co; // @[wallace.scala 70:18]
  assign FullAdder_616_io_ci = FullAdder_451_io_co; // @[wallace.scala 71:19]
  assign FullAdder_617_io_a = FullAdder_452_io_co; // @[wallace.scala 69:18]
  assign FullAdder_617_io_b = FullAdder_453_io_co; // @[wallace.scala 70:18]
  assign FullAdder_617_io_ci = FullAdder_454_io_co; // @[wallace.scala 71:19]
  assign FullAdder_618_io_a = FullAdder_210_io_co; // @[wallace.scala 69:18]
  assign FullAdder_618_io_b = FullAdder_450_io_s; // @[wallace.scala 70:18]
  assign FullAdder_618_io_ci = FullAdder_451_io_s; // @[wallace.scala 71:19]
  assign FullAdder_619_io_a = FullAdder_452_io_s; // @[wallace.scala 69:18]
  assign FullAdder_619_io_b = FullAdder_453_io_s; // @[wallace.scala 70:18]
  assign FullAdder_619_io_ci = FullAdder_454_io_s; // @[wallace.scala 71:19]
  assign FullAdder_620_io_a = FullAdder_455_io_s; // @[wallace.scala 69:18]
  assign FullAdder_620_io_b = FullAdder_456_io_co; // @[wallace.scala 70:18]
  assign FullAdder_620_io_ci = FullAdder_457_io_co; // @[wallace.scala 71:19]
  assign FullAdder_621_io_a = FullAdder_458_io_co; // @[wallace.scala 69:18]
  assign FullAdder_621_io_b = FullAdder_459_io_co; // @[wallace.scala 70:18]
  assign FullAdder_621_io_ci = FullAdder_460_io_co; // @[wallace.scala 71:19]
  assign FullAdder_622_io_a = FullAdder_456_io_s; // @[wallace.scala 69:18]
  assign FullAdder_622_io_b = FullAdder_457_io_s; // @[wallace.scala 70:18]
  assign FullAdder_622_io_ci = FullAdder_458_io_s; // @[wallace.scala 71:19]
  assign FullAdder_623_io_a = FullAdder_459_io_s; // @[wallace.scala 69:18]
  assign FullAdder_623_io_b = FullAdder_460_io_s; // @[wallace.scala 70:18]
  assign FullAdder_623_io_ci = FullAdder_461_io_s; // @[wallace.scala 71:19]
  assign FullAdder_624_io_a = FullAdder_462_io_co; // @[wallace.scala 69:18]
  assign FullAdder_624_io_b = FullAdder_463_io_co; // @[wallace.scala 70:18]
  assign FullAdder_624_io_ci = FullAdder_464_io_co; // @[wallace.scala 71:19]
  assign FullAdder_625_io_a = FullAdder_465_io_co; // @[wallace.scala 69:18]
  assign FullAdder_625_io_b = FullAdder_466_io_co; // @[wallace.scala 70:18]
  assign FullAdder_625_io_ci = HalfAdder_25_io_co; // @[wallace.scala 71:19]
  assign FullAdder_626_io_a = FullAdder_462_io_s; // @[wallace.scala 69:18]
  assign FullAdder_626_io_b = FullAdder_463_io_s; // @[wallace.scala 70:18]
  assign FullAdder_626_io_ci = FullAdder_464_io_s; // @[wallace.scala 71:19]
  assign FullAdder_627_io_a = FullAdder_465_io_s; // @[wallace.scala 69:18]
  assign FullAdder_627_io_b = FullAdder_466_io_s; // @[wallace.scala 70:18]
  assign FullAdder_627_io_ci = HalfAdder_25_io_s; // @[wallace.scala 71:19]
  assign FullAdder_628_io_a = FullAdder_467_io_co; // @[wallace.scala 69:18]
  assign FullAdder_628_io_b = FullAdder_468_io_co; // @[wallace.scala 70:18]
  assign FullAdder_628_io_ci = FullAdder_469_io_co; // @[wallace.scala 71:19]
  assign FullAdder_629_io_a = FullAdder_470_io_co; // @[wallace.scala 69:18]
  assign FullAdder_629_io_b = FullAdder_471_io_co; // @[wallace.scala 70:18]
  assign FullAdder_629_io_ci = HalfAdder_26_io_co; // @[wallace.scala 71:19]
  assign FullAdder_630_io_a = FullAdder_467_io_s; // @[wallace.scala 69:18]
  assign FullAdder_630_io_b = FullAdder_468_io_s; // @[wallace.scala 70:18]
  assign FullAdder_630_io_ci = FullAdder_469_io_s; // @[wallace.scala 71:19]
  assign FullAdder_631_io_a = FullAdder_470_io_s; // @[wallace.scala 69:18]
  assign FullAdder_631_io_b = FullAdder_471_io_s; // @[wallace.scala 70:18]
  assign FullAdder_631_io_ci = HalfAdder_26_io_s; // @[wallace.scala 71:19]
  assign FullAdder_632_io_a = FullAdder_472_io_co; // @[wallace.scala 69:18]
  assign FullAdder_632_io_b = FullAdder_473_io_co; // @[wallace.scala 70:18]
  assign FullAdder_632_io_ci = FullAdder_474_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_46_io_a = FullAdder_475_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_46_io_b = FullAdder_476_io_co; // @[wallace.scala 60:18]
  assign FullAdder_633_io_a = FullAdder_472_io_s; // @[wallace.scala 69:18]
  assign FullAdder_633_io_b = FullAdder_473_io_s; // @[wallace.scala 70:18]
  assign FullAdder_633_io_ci = FullAdder_474_io_s; // @[wallace.scala 71:19]
  assign FullAdder_634_io_a = FullAdder_475_io_s; // @[wallace.scala 69:18]
  assign FullAdder_634_io_b = FullAdder_476_io_s; // @[wallace.scala 70:18]
  assign FullAdder_634_io_ci = FullAdder_477_io_co; // @[wallace.scala 71:19]
  assign FullAdder_635_io_a = FullAdder_478_io_co; // @[wallace.scala 69:18]
  assign FullAdder_635_io_b = FullAdder_479_io_co; // @[wallace.scala 70:18]
  assign FullAdder_635_io_ci = FullAdder_480_io_co; // @[wallace.scala 71:19]
  assign FullAdder_636_io_a = FullAdder_248_io_co; // @[wallace.scala 69:18]
  assign FullAdder_636_io_b = FullAdder_477_io_s; // @[wallace.scala 70:18]
  assign FullAdder_636_io_ci = FullAdder_478_io_s; // @[wallace.scala 71:19]
  assign FullAdder_637_io_a = FullAdder_479_io_s; // @[wallace.scala 69:18]
  assign FullAdder_637_io_b = FullAdder_480_io_s; // @[wallace.scala 70:18]
  assign FullAdder_637_io_ci = FullAdder_481_io_s; // @[wallace.scala 71:19]
  assign FullAdder_638_io_a = FullAdder_482_io_co; // @[wallace.scala 69:18]
  assign FullAdder_638_io_b = FullAdder_483_io_co; // @[wallace.scala 70:18]
  assign FullAdder_638_io_ci = FullAdder_484_io_co; // @[wallace.scala 71:19]
  assign FullAdder_639_io_a = FullAdder_482_io_s; // @[wallace.scala 69:18]
  assign FullAdder_639_io_b = FullAdder_483_io_s; // @[wallace.scala 70:18]
  assign FullAdder_639_io_ci = FullAdder_484_io_s; // @[wallace.scala 71:19]
  assign FullAdder_640_io_a = FullAdder_485_io_s; // @[wallace.scala 69:18]
  assign FullAdder_640_io_b = FullAdder_486_io_s; // @[wallace.scala 70:18]
  assign FullAdder_640_io_ci = FullAdder_487_io_co; // @[wallace.scala 71:19]
  assign FullAdder_641_io_a = FullAdder_488_io_co; // @[wallace.scala 69:18]
  assign FullAdder_641_io_b = FullAdder_489_io_co; // @[wallace.scala 70:18]
  assign FullAdder_641_io_ci = FullAdder_490_io_co; // @[wallace.scala 71:19]
  assign FullAdder_642_io_a = FullAdder_261_io_co; // @[wallace.scala 69:18]
  assign FullAdder_642_io_b = FullAdder_487_io_s; // @[wallace.scala 70:18]
  assign FullAdder_642_io_ci = FullAdder_488_io_s; // @[wallace.scala 71:19]
  assign FullAdder_643_io_a = FullAdder_489_io_s; // @[wallace.scala 69:18]
  assign FullAdder_643_io_b = FullAdder_490_io_s; // @[wallace.scala 70:18]
  assign FullAdder_643_io_ci = FullAdder_491_io_co; // @[wallace.scala 71:19]
  assign FullAdder_644_io_a = FullAdder_492_io_co; // @[wallace.scala 69:18]
  assign FullAdder_644_io_b = FullAdder_493_io_co; // @[wallace.scala 70:18]
  assign FullAdder_644_io_ci = FullAdder_494_io_co; // @[wallace.scala 71:19]
  assign FullAdder_645_io_a = FullAdder_266_io_co; // @[wallace.scala 69:18]
  assign FullAdder_645_io_b = FullAdder_267_io_co; // @[wallace.scala 70:18]
  assign FullAdder_645_io_ci = FullAdder_491_io_s; // @[wallace.scala 71:19]
  assign FullAdder_646_io_a = FullAdder_492_io_s; // @[wallace.scala 69:18]
  assign FullAdder_646_io_b = FullAdder_493_io_s; // @[wallace.scala 70:18]
  assign FullAdder_646_io_ci = FullAdder_494_io_s; // @[wallace.scala 71:19]
  assign FullAdder_647_io_a = FullAdder_495_io_co; // @[wallace.scala 69:18]
  assign FullAdder_647_io_b = FullAdder_496_io_co; // @[wallace.scala 70:18]
  assign FullAdder_647_io_ci = FullAdder_497_io_co; // @[wallace.scala 71:19]
  assign FullAdder_648_io_a = FullAdder_273_io_co; // @[wallace.scala 69:18]
  assign FullAdder_648_io_b = FullAdder_495_io_s; // @[wallace.scala 70:18]
  assign FullAdder_648_io_ci = FullAdder_496_io_s; // @[wallace.scala 71:19]
  assign FullAdder_649_io_a = FullAdder_497_io_s; // @[wallace.scala 69:18]
  assign FullAdder_649_io_b = FullAdder_498_io_s; // @[wallace.scala 70:18]
  assign FullAdder_649_io_ci = FullAdder_499_io_co; // @[wallace.scala 71:19]
  assign FullAdder_650_io_a = FullAdder_500_io_co; // @[wallace.scala 69:18]
  assign FullAdder_650_io_b = FullAdder_501_io_co; // @[wallace.scala 70:18]
  assign FullAdder_650_io_ci = FullAdder_502_io_co; // @[wallace.scala 71:19]
  assign FullAdder_651_io_a = FullAdder_499_io_s; // @[wallace.scala 69:18]
  assign FullAdder_651_io_b = FullAdder_500_io_s; // @[wallace.scala 70:18]
  assign FullAdder_651_io_ci = FullAdder_501_io_s; // @[wallace.scala 71:19]
  assign FullAdder_652_io_a = FullAdder_502_io_s; // @[wallace.scala 69:18]
  assign FullAdder_652_io_b = FullAdder_503_io_co; // @[wallace.scala 70:18]
  assign FullAdder_652_io_ci = FullAdder_504_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_47_io_a = FullAdder_505_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_47_io_b = HalfAdder_27_io_co; // @[wallace.scala 60:18]
  assign FullAdder_653_io_a = FullAdder_503_io_s; // @[wallace.scala 69:18]
  assign FullAdder_653_io_b = FullAdder_504_io_s; // @[wallace.scala 70:18]
  assign FullAdder_653_io_ci = FullAdder_505_io_s; // @[wallace.scala 71:19]
  assign FullAdder_654_io_a = HalfAdder_27_io_s; // @[wallace.scala 69:18]
  assign FullAdder_654_io_b = FullAdder_506_io_co; // @[wallace.scala 70:18]
  assign FullAdder_654_io_ci = FullAdder_507_io_co; // @[wallace.scala 71:19]
  assign FullAdder_655_io_a = FullAdder_287_io_co; // @[wallace.scala 69:18]
  assign FullAdder_655_io_b = FullAdder_288_io_co; // @[wallace.scala 70:18]
  assign FullAdder_655_io_ci = FullAdder_506_io_s; // @[wallace.scala 71:19]
  assign FullAdder_656_io_a = FullAdder_507_io_s; // @[wallace.scala 69:18]
  assign FullAdder_656_io_b = FullAdder_508_io_s; // @[wallace.scala 70:18]
  assign FullAdder_656_io_ci = FullAdder_509_io_co; // @[wallace.scala 71:19]
  assign FullAdder_657_io_a = FullAdder_509_io_s; // @[wallace.scala 69:18]
  assign FullAdder_657_io_b = FullAdder_510_io_s; // @[wallace.scala 70:18]
  assign FullAdder_657_io_ci = FullAdder_511_io_s; // @[wallace.scala 71:19]
  assign FullAdder_658_io_a = FullAdder_512_io_co; // @[wallace.scala 69:18]
  assign FullAdder_658_io_b = FullAdder_513_io_co; // @[wallace.scala 70:18]
  assign FullAdder_658_io_ci = FullAdder_514_io_co; // @[wallace.scala 71:19]
  assign FullAdder_659_io_a = FullAdder_296_io_co; // @[wallace.scala 69:18]
  assign FullAdder_659_io_b = FullAdder_512_io_s; // @[wallace.scala 70:18]
  assign FullAdder_659_io_ci = FullAdder_513_io_s; // @[wallace.scala 71:19]
  assign FullAdder_660_io_a = FullAdder_514_io_s; // @[wallace.scala 69:18]
  assign FullAdder_660_io_b = FullAdder_515_io_co; // @[wallace.scala 70:18]
  assign FullAdder_660_io_ci = FullAdder_516_io_co; // @[wallace.scala 71:19]
  assign FullAdder_661_io_a = FullAdder_515_io_s; // @[wallace.scala 69:18]
  assign FullAdder_661_io_b = FullAdder_516_io_s; // @[wallace.scala 70:18]
  assign FullAdder_661_io_ci = FullAdder_517_io_s; // @[wallace.scala 71:19]
  assign FullAdder_662_io_a = FullAdder_518_io_co; // @[wallace.scala 69:18]
  assign FullAdder_662_io_b = FullAdder_519_io_co; // @[wallace.scala 70:18]
  assign FullAdder_662_io_ci = HalfAdder_28_io_co; // @[wallace.scala 71:19]
  assign FullAdder_663_io_a = FullAdder_518_io_s; // @[wallace.scala 69:18]
  assign FullAdder_663_io_b = FullAdder_519_io_s; // @[wallace.scala 70:18]
  assign FullAdder_663_io_ci = HalfAdder_28_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_48_io_a = FullAdder_520_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_48_io_b = FullAdder_521_io_co; // @[wallace.scala 60:18]
  assign FullAdder_664_io_a = FullAdder_306_io_co; // @[wallace.scala 69:18]
  assign FullAdder_664_io_b = FullAdder_520_io_s; // @[wallace.scala 70:18]
  assign FullAdder_664_io_ci = FullAdder_521_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_49_io_a = FullAdder_522_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_49_io_b = FullAdder_523_io_co; // @[wallace.scala 60:18]
  assign FullAdder_665_io_a = FullAdder_309_io_co; // @[wallace.scala 69:18]
  assign FullAdder_665_io_b = FullAdder_522_io_s; // @[wallace.scala 70:18]
  assign FullAdder_665_io_ci = FullAdder_523_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_50_io_a = FullAdder_524_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_50_io_b = FullAdder_525_io_co; // @[wallace.scala 60:18]
  assign FullAdder_666_io_a = FullAdder_524_io_s; // @[wallace.scala 69:18]
  assign FullAdder_666_io_b = FullAdder_525_io_s; // @[wallace.scala 70:18]
  assign FullAdder_666_io_ci = FullAdder_526_io_co; // @[wallace.scala 71:19]
  assign FullAdder_667_io_a = FullAdder_526_io_s; // @[wallace.scala 69:18]
  assign FullAdder_667_io_b = HalfAdder_29_io_s; // @[wallace.scala 70:18]
  assign FullAdder_667_io_ci = FullAdder_527_io_co; // @[wallace.scala 71:19]
  assign FullAdder_668_io_a = FullAdder_527_io_s; // @[wallace.scala 69:18]
  assign FullAdder_668_io_b = HalfAdder_30_io_s; // @[wallace.scala 70:18]
  assign FullAdder_668_io_ci = HalfAdder_31_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_51_io_a = HalfAdder_31_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_51_io_b = HalfAdder_32_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_52_io_a = FullAdder_317_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_52_io_b = HalfAdder_33_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_53_io_a = HalfAdder_34_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_53_io_b = HalfAdder_35_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_54_io_a = HalfAdder_35_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_54_io_b = HalfAdder_36_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_55_io_a = FullAdder_319_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_55_io_b = HalfAdder_36_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_56_io_a = FullAdder_529_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_56_io_b = FullAdder_530_io_co; // @[wallace.scala 60:18]
  assign FullAdder_669_io_a = HalfAdder_17_io_co; // @[wallace.scala 69:18]
  assign FullAdder_669_io_b = FullAdder_531_io_s; // @[wallace.scala 70:18]
  assign FullAdder_669_io_ci = FullAdder_532_io_co; // @[wallace.scala 71:19]
  assign FullAdder_670_io_a = FullAdder_324_io_co; // @[wallace.scala 69:18]
  assign FullAdder_670_io_b = FullAdder_532_io_s; // @[wallace.scala 70:18]
  assign FullAdder_670_io_ci = FullAdder_533_io_co; // @[wallace.scala 71:19]
  assign FullAdder_671_io_a = FullAdder_325_io_co; // @[wallace.scala 69:18]
  assign FullAdder_671_io_b = FullAdder_326_io_co; // @[wallace.scala 70:18]
  assign FullAdder_671_io_ci = FullAdder_533_io_s; // @[wallace.scala 71:19]
  assign FullAdder_672_io_a = FullAdder_534_io_s; // @[wallace.scala 69:18]
  assign FullAdder_672_io_b = HalfAdder_37_io_s; // @[wallace.scala 70:18]
  assign FullAdder_672_io_ci = FullAdder_535_io_co; // @[wallace.scala 71:19]
  assign FullAdder_673_io_a = FullAdder_535_io_s; // @[wallace.scala 69:18]
  assign FullAdder_673_io_b = FullAdder_536_io_s; // @[wallace.scala 70:18]
  assign FullAdder_673_io_ci = FullAdder_537_io_co; // @[wallace.scala 71:19]
  assign FullAdder_674_io_a = FullAdder_537_io_s; // @[wallace.scala 69:18]
  assign FullAdder_674_io_b = FullAdder_538_io_s; // @[wallace.scala 70:18]
  assign FullAdder_674_io_ci = FullAdder_539_io_co; // @[wallace.scala 71:19]
  assign FullAdder_675_io_a = FullAdder_539_io_s; // @[wallace.scala 69:18]
  assign FullAdder_675_io_b = FullAdder_540_io_s; // @[wallace.scala 70:18]
  assign FullAdder_675_io_ci = FullAdder_541_io_co; // @[wallace.scala 71:19]
  assign FullAdder_676_io_a = FullAdder_338_io_co; // @[wallace.scala 69:18]
  assign FullAdder_676_io_b = FullAdder_541_io_s; // @[wallace.scala 70:18]
  assign FullAdder_676_io_ci = FullAdder_542_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_57_io_a = FullAdder_543_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_57_io_b = FullAdder_544_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_58_io_a = FullAdder_341_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_58_io_b = FullAdder_543_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_59_io_a = FullAdder_544_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_59_io_b = FullAdder_545_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_60_io_a = FullAdder_546_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_60_io_b = HalfAdder_38_io_co; // @[wallace.scala 60:18]
  assign FullAdder_677_io_a = FullAdder_545_io_s; // @[wallace.scala 69:18]
  assign FullAdder_677_io_b = FullAdder_546_io_s; // @[wallace.scala 70:18]
  assign FullAdder_677_io_ci = HalfAdder_38_io_s; // @[wallace.scala 71:19]
  assign FullAdder_678_io_a = FullAdder_547_io_co; // @[wallace.scala 69:18]
  assign FullAdder_678_io_b = FullAdder_548_io_co; // @[wallace.scala 70:18]
  assign FullAdder_678_io_ci = HalfAdder_39_io_co; // @[wallace.scala 71:19]
  assign FullAdder_679_io_a = FullAdder_547_io_s; // @[wallace.scala 69:18]
  assign FullAdder_679_io_b = FullAdder_548_io_s; // @[wallace.scala 70:18]
  assign FullAdder_679_io_ci = HalfAdder_39_io_s; // @[wallace.scala 71:19]
  assign FullAdder_680_io_a = FullAdder_549_io_co; // @[wallace.scala 69:18]
  assign FullAdder_680_io_b = FullAdder_550_io_co; // @[wallace.scala 70:18]
  assign FullAdder_680_io_ci = HalfAdder_40_io_co; // @[wallace.scala 71:19]
  assign FullAdder_681_io_a = FullAdder_549_io_s; // @[wallace.scala 69:18]
  assign FullAdder_681_io_b = FullAdder_550_io_s; // @[wallace.scala 70:18]
  assign FullAdder_681_io_ci = HalfAdder_40_io_s; // @[wallace.scala 71:19]
  assign FullAdder_682_io_a = FullAdder_551_io_co; // @[wallace.scala 69:18]
  assign FullAdder_682_io_b = FullAdder_552_io_co; // @[wallace.scala 70:18]
  assign FullAdder_682_io_ci = HalfAdder_41_io_co; // @[wallace.scala 71:19]
  assign FullAdder_683_io_a = FullAdder_551_io_s; // @[wallace.scala 69:18]
  assign FullAdder_683_io_b = FullAdder_552_io_s; // @[wallace.scala 70:18]
  assign FullAdder_683_io_ci = HalfAdder_41_io_s; // @[wallace.scala 71:19]
  assign FullAdder_684_io_a = FullAdder_553_io_co; // @[wallace.scala 69:18]
  assign FullAdder_684_io_b = FullAdder_554_io_co; // @[wallace.scala 70:18]
  assign FullAdder_684_io_ci = FullAdder_555_io_co; // @[wallace.scala 71:19]
  assign FullAdder_685_io_a = FullAdder_362_io_co; // @[wallace.scala 69:18]
  assign FullAdder_685_io_b = FullAdder_553_io_s; // @[wallace.scala 70:18]
  assign FullAdder_685_io_ci = FullAdder_554_io_s; // @[wallace.scala 71:19]
  assign FullAdder_686_io_a = FullAdder_555_io_s; // @[wallace.scala 69:18]
  assign FullAdder_686_io_b = FullAdder_556_io_co; // @[wallace.scala 70:18]
  assign FullAdder_686_io_ci = FullAdder_557_io_co; // @[wallace.scala 71:19]
  assign FullAdder_687_io_a = HalfAdder_21_io_co; // @[wallace.scala 69:18]
  assign FullAdder_687_io_b = FullAdder_556_io_s; // @[wallace.scala 70:18]
  assign FullAdder_687_io_ci = FullAdder_557_io_s; // @[wallace.scala 71:19]
  assign FullAdder_688_io_a = FullAdder_558_io_s; // @[wallace.scala 69:18]
  assign FullAdder_688_io_b = FullAdder_559_io_co; // @[wallace.scala 70:18]
  assign FullAdder_688_io_ci = FullAdder_560_io_co; // @[wallace.scala 71:19]
  assign FullAdder_689_io_a = FullAdder_371_io_co; // @[wallace.scala 69:18]
  assign FullAdder_689_io_b = FullAdder_559_io_s; // @[wallace.scala 70:18]
  assign FullAdder_689_io_ci = FullAdder_560_io_s; // @[wallace.scala 71:19]
  assign FullAdder_690_io_a = FullAdder_561_io_s; // @[wallace.scala 69:18]
  assign FullAdder_690_io_b = FullAdder_562_io_co; // @[wallace.scala 70:18]
  assign FullAdder_690_io_ci = FullAdder_563_io_co; // @[wallace.scala 71:19]
  assign FullAdder_691_io_a = FullAdder_562_io_s; // @[wallace.scala 69:18]
  assign FullAdder_691_io_b = FullAdder_563_io_s; // @[wallace.scala 70:18]
  assign FullAdder_691_io_ci = FullAdder_564_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_61_io_a = HalfAdder_42_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_61_io_b = FullAdder_565_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_62_io_a = FullAdder_566_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_62_io_b = FullAdder_567_io_co; // @[wallace.scala 60:18]
  assign FullAdder_692_io_a = FullAdder_565_io_s; // @[wallace.scala 69:18]
  assign FullAdder_692_io_b = FullAdder_566_io_s; // @[wallace.scala 70:18]
  assign FullAdder_692_io_ci = FullAdder_567_io_s; // @[wallace.scala 71:19]
  assign FullAdder_693_io_a = HalfAdder_43_io_s; // @[wallace.scala 69:18]
  assign FullAdder_693_io_b = FullAdder_568_io_co; // @[wallace.scala 70:18]
  assign FullAdder_693_io_ci = FullAdder_569_io_co; // @[wallace.scala 71:19]
  assign FullAdder_694_io_a = FullAdder_568_io_s; // @[wallace.scala 69:18]
  assign FullAdder_694_io_b = FullAdder_569_io_s; // @[wallace.scala 70:18]
  assign FullAdder_694_io_ci = FullAdder_570_io_s; // @[wallace.scala 71:19]
  assign FullAdder_695_io_a = FullAdder_571_io_s; // @[wallace.scala 69:18]
  assign FullAdder_695_io_b = FullAdder_572_io_co; // @[wallace.scala 70:18]
  assign FullAdder_695_io_ci = FullAdder_573_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_63_io_a = FullAdder_574_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_63_io_b = FullAdder_575_io_co; // @[wallace.scala 60:18]
  assign FullAdder_696_io_a = FullAdder_572_io_s; // @[wallace.scala 69:18]
  assign FullAdder_696_io_b = FullAdder_573_io_s; // @[wallace.scala 70:18]
  assign FullAdder_696_io_ci = FullAdder_574_io_s; // @[wallace.scala 71:19]
  assign FullAdder_697_io_a = FullAdder_575_io_s; // @[wallace.scala 69:18]
  assign FullAdder_697_io_b = FullAdder_576_io_co; // @[wallace.scala 70:18]
  assign FullAdder_697_io_ci = FullAdder_577_io_co; // @[wallace.scala 71:19]
  assign FullAdder_698_io_a = FullAdder_398_io_co; // @[wallace.scala 69:18]
  assign FullAdder_698_io_b = FullAdder_576_io_s; // @[wallace.scala 70:18]
  assign FullAdder_698_io_ci = FullAdder_577_io_s; // @[wallace.scala 71:19]
  assign FullAdder_699_io_a = FullAdder_578_io_s; // @[wallace.scala 69:18]
  assign FullAdder_699_io_b = FullAdder_579_io_s; // @[wallace.scala 70:18]
  assign FullAdder_699_io_ci = FullAdder_580_io_co; // @[wallace.scala 71:19]
  assign FullAdder_700_io_a = FullAdder_581_io_co; // @[wallace.scala 69:18]
  assign FullAdder_700_io_b = FullAdder_582_io_co; // @[wallace.scala 70:18]
  assign FullAdder_700_io_ci = FullAdder_583_io_co; // @[wallace.scala 71:19]
  assign FullAdder_701_io_a = HalfAdder_23_io_co; // @[wallace.scala 69:18]
  assign FullAdder_701_io_b = FullAdder_580_io_s; // @[wallace.scala 70:18]
  assign FullAdder_701_io_ci = FullAdder_581_io_s; // @[wallace.scala 71:19]
  assign FullAdder_702_io_a = FullAdder_582_io_s; // @[wallace.scala 69:18]
  assign FullAdder_702_io_b = FullAdder_583_io_s; // @[wallace.scala 70:18]
  assign FullAdder_702_io_ci = FullAdder_584_io_co; // @[wallace.scala 71:19]
  assign FullAdder_703_io_a = FullAdder_585_io_co; // @[wallace.scala 69:18]
  assign FullAdder_703_io_b = FullAdder_586_io_co; // @[wallace.scala 70:18]
  assign FullAdder_703_io_ci = FullAdder_587_io_co; // @[wallace.scala 71:19]
  assign FullAdder_704_io_a = FullAdder_584_io_s; // @[wallace.scala 69:18]
  assign FullAdder_704_io_b = FullAdder_585_io_s; // @[wallace.scala 70:18]
  assign FullAdder_704_io_ci = FullAdder_586_io_s; // @[wallace.scala 71:19]
  assign FullAdder_705_io_a = FullAdder_587_io_s; // @[wallace.scala 69:18]
  assign FullAdder_705_io_b = HalfAdder_44_io_s; // @[wallace.scala 70:18]
  assign FullAdder_705_io_ci = FullAdder_588_io_co; // @[wallace.scala 71:19]
  assign FullAdder_706_io_a = FullAdder_589_io_co; // @[wallace.scala 69:18]
  assign FullAdder_706_io_b = FullAdder_590_io_co; // @[wallace.scala 70:18]
  assign FullAdder_706_io_ci = FullAdder_591_io_co; // @[wallace.scala 71:19]
  assign FullAdder_707_io_a = FullAdder_416_io_co; // @[wallace.scala 69:18]
  assign FullAdder_707_io_b = FullAdder_588_io_s; // @[wallace.scala 70:18]
  assign FullAdder_707_io_ci = FullAdder_589_io_s; // @[wallace.scala 71:19]
  assign FullAdder_708_io_a = FullAdder_590_io_s; // @[wallace.scala 69:18]
  assign FullAdder_708_io_b = FullAdder_591_io_s; // @[wallace.scala 70:18]
  assign FullAdder_708_io_ci = FullAdder_592_io_co; // @[wallace.scala 71:19]
  assign FullAdder_709_io_a = FullAdder_593_io_co; // @[wallace.scala 69:18]
  assign FullAdder_709_io_b = FullAdder_594_io_co; // @[wallace.scala 70:18]
  assign FullAdder_709_io_ci = FullAdder_595_io_co; // @[wallace.scala 71:19]
  assign FullAdder_710_io_a = FullAdder_592_io_s; // @[wallace.scala 69:18]
  assign FullAdder_710_io_b = FullAdder_593_io_s; // @[wallace.scala 70:18]
  assign FullAdder_710_io_ci = FullAdder_594_io_s; // @[wallace.scala 71:19]
  assign FullAdder_711_io_a = FullAdder_595_io_s; // @[wallace.scala 69:18]
  assign FullAdder_711_io_b = FullAdder_596_io_s; // @[wallace.scala 70:18]
  assign FullAdder_711_io_ci = FullAdder_597_io_co; // @[wallace.scala 71:19]
  assign FullAdder_712_io_a = FullAdder_598_io_co; // @[wallace.scala 69:18]
  assign FullAdder_712_io_b = FullAdder_599_io_co; // @[wallace.scala 70:18]
  assign FullAdder_712_io_ci = FullAdder_600_io_co; // @[wallace.scala 71:19]
  assign FullAdder_713_io_a = FullAdder_597_io_s; // @[wallace.scala 69:18]
  assign FullAdder_713_io_b = FullAdder_598_io_s; // @[wallace.scala 70:18]
  assign FullAdder_713_io_ci = FullAdder_599_io_s; // @[wallace.scala 71:19]
  assign FullAdder_714_io_a = FullAdder_600_io_s; // @[wallace.scala 69:18]
  assign FullAdder_714_io_b = HalfAdder_45_io_s; // @[wallace.scala 70:18]
  assign FullAdder_714_io_ci = FullAdder_601_io_co; // @[wallace.scala 71:19]
  assign FullAdder_715_io_a = FullAdder_602_io_co; // @[wallace.scala 69:18]
  assign FullAdder_715_io_b = FullAdder_603_io_co; // @[wallace.scala 70:18]
  assign FullAdder_715_io_ci = FullAdder_604_io_co; // @[wallace.scala 71:19]
  assign FullAdder_716_io_a = FullAdder_601_io_s; // @[wallace.scala 69:18]
  assign FullAdder_716_io_b = FullAdder_602_io_s; // @[wallace.scala 70:18]
  assign FullAdder_716_io_ci = FullAdder_603_io_s; // @[wallace.scala 71:19]
  assign FullAdder_717_io_a = FullAdder_604_io_s; // @[wallace.scala 69:18]
  assign FullAdder_717_io_b = FullAdder_605_io_s; // @[wallace.scala 70:18]
  assign FullAdder_717_io_ci = FullAdder_606_io_co; // @[wallace.scala 71:19]
  assign FullAdder_718_io_a = FullAdder_607_io_co; // @[wallace.scala 69:18]
  assign FullAdder_718_io_b = FullAdder_608_io_co; // @[wallace.scala 70:18]
  assign FullAdder_718_io_ci = FullAdder_609_io_co; // @[wallace.scala 71:19]
  assign FullAdder_719_io_a = FullAdder_443_io_co; // @[wallace.scala 69:18]
  assign FullAdder_719_io_b = FullAdder_606_io_s; // @[wallace.scala 70:18]
  assign FullAdder_719_io_ci = FullAdder_607_io_s; // @[wallace.scala 71:19]
  assign FullAdder_720_io_a = FullAdder_608_io_s; // @[wallace.scala 69:18]
  assign FullAdder_720_io_b = FullAdder_609_io_s; // @[wallace.scala 70:18]
  assign FullAdder_720_io_ci = FullAdder_610_io_co; // @[wallace.scala 71:19]
  assign FullAdder_721_io_a = FullAdder_611_io_co; // @[wallace.scala 69:18]
  assign FullAdder_721_io_b = FullAdder_612_io_co; // @[wallace.scala 70:18]
  assign FullAdder_721_io_ci = FullAdder_613_io_co; // @[wallace.scala 71:19]
  assign FullAdder_722_io_a = FullAdder_448_io_co; // @[wallace.scala 69:18]
  assign FullAdder_722_io_b = FullAdder_449_io_co; // @[wallace.scala 70:18]
  assign FullAdder_722_io_ci = FullAdder_610_io_s; // @[wallace.scala 71:19]
  assign FullAdder_723_io_a = FullAdder_611_io_s; // @[wallace.scala 69:18]
  assign FullAdder_723_io_b = FullAdder_612_io_s; // @[wallace.scala 70:18]
  assign FullAdder_723_io_ci = FullAdder_613_io_s; // @[wallace.scala 71:19]
  assign FullAdder_724_io_a = FullAdder_614_io_co; // @[wallace.scala 69:18]
  assign FullAdder_724_io_b = FullAdder_615_io_co; // @[wallace.scala 70:18]
  assign FullAdder_724_io_ci = FullAdder_616_io_co; // @[wallace.scala 71:19]
  assign FullAdder_725_io_a = FullAdder_455_io_co; // @[wallace.scala 69:18]
  assign FullAdder_725_io_b = FullAdder_614_io_s; // @[wallace.scala 70:18]
  assign FullAdder_725_io_ci = FullAdder_615_io_s; // @[wallace.scala 71:19]
  assign FullAdder_726_io_a = FullAdder_616_io_s; // @[wallace.scala 69:18]
  assign FullAdder_726_io_b = FullAdder_617_io_s; // @[wallace.scala 70:18]
  assign FullAdder_726_io_ci = FullAdder_618_io_co; // @[wallace.scala 71:19]
  assign FullAdder_727_io_a = FullAdder_619_io_co; // @[wallace.scala 69:18]
  assign FullAdder_727_io_b = FullAdder_620_io_co; // @[wallace.scala 70:18]
  assign FullAdder_727_io_ci = FullAdder_621_io_co; // @[wallace.scala 71:19]
  assign FullAdder_728_io_a = FullAdder_461_io_co; // @[wallace.scala 69:18]
  assign FullAdder_728_io_b = FullAdder_618_io_s; // @[wallace.scala 70:18]
  assign FullAdder_728_io_ci = FullAdder_619_io_s; // @[wallace.scala 71:19]
  assign FullAdder_729_io_a = FullAdder_620_io_s; // @[wallace.scala 69:18]
  assign FullAdder_729_io_b = FullAdder_621_io_s; // @[wallace.scala 70:18]
  assign FullAdder_729_io_ci = FullAdder_622_io_co; // @[wallace.scala 71:19]
  assign FullAdder_730_io_a = FullAdder_623_io_co; // @[wallace.scala 69:18]
  assign FullAdder_730_io_b = FullAdder_624_io_co; // @[wallace.scala 70:18]
  assign FullAdder_730_io_ci = FullAdder_625_io_co; // @[wallace.scala 71:19]
  assign FullAdder_731_io_a = FullAdder_622_io_s; // @[wallace.scala 69:18]
  assign FullAdder_731_io_b = FullAdder_623_io_s; // @[wallace.scala 70:18]
  assign FullAdder_731_io_ci = FullAdder_624_io_s; // @[wallace.scala 71:19]
  assign FullAdder_732_io_a = FullAdder_625_io_s; // @[wallace.scala 69:18]
  assign FullAdder_732_io_b = FullAdder_626_io_co; // @[wallace.scala 70:18]
  assign FullAdder_732_io_ci = FullAdder_627_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_64_io_a = FullAdder_628_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_64_io_b = FullAdder_629_io_co; // @[wallace.scala 60:18]
  assign FullAdder_733_io_a = FullAdder_626_io_s; // @[wallace.scala 69:18]
  assign FullAdder_733_io_b = FullAdder_627_io_s; // @[wallace.scala 70:18]
  assign FullAdder_733_io_ci = FullAdder_628_io_s; // @[wallace.scala 71:19]
  assign FullAdder_734_io_a = FullAdder_629_io_s; // @[wallace.scala 69:18]
  assign FullAdder_734_io_b = FullAdder_630_io_co; // @[wallace.scala 70:18]
  assign FullAdder_734_io_ci = FullAdder_631_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_65_io_a = FullAdder_632_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_65_io_b = HalfAdder_46_io_co; // @[wallace.scala 60:18]
  assign FullAdder_735_io_a = FullAdder_630_io_s; // @[wallace.scala 69:18]
  assign FullAdder_735_io_b = FullAdder_631_io_s; // @[wallace.scala 70:18]
  assign FullAdder_735_io_ci = FullAdder_632_io_s; // @[wallace.scala 71:19]
  assign FullAdder_736_io_a = HalfAdder_46_io_s; // @[wallace.scala 69:18]
  assign FullAdder_736_io_b = FullAdder_633_io_co; // @[wallace.scala 70:18]
  assign FullAdder_736_io_ci = FullAdder_634_io_co; // @[wallace.scala 71:19]
  assign FullAdder_737_io_a = FullAdder_481_io_co; // @[wallace.scala 69:18]
  assign FullAdder_737_io_b = FullAdder_633_io_s; // @[wallace.scala 70:18]
  assign FullAdder_737_io_ci = FullAdder_634_io_s; // @[wallace.scala 71:19]
  assign FullAdder_738_io_a = FullAdder_635_io_s; // @[wallace.scala 69:18]
  assign FullAdder_738_io_b = FullAdder_636_io_co; // @[wallace.scala 70:18]
  assign FullAdder_738_io_ci = FullAdder_637_io_co; // @[wallace.scala 71:19]
  assign FullAdder_739_io_a = FullAdder_485_io_co; // @[wallace.scala 69:18]
  assign FullAdder_739_io_b = FullAdder_486_io_co; // @[wallace.scala 70:18]
  assign FullAdder_739_io_ci = FullAdder_636_io_s; // @[wallace.scala 71:19]
  assign FullAdder_740_io_a = FullAdder_637_io_s; // @[wallace.scala 69:18]
  assign FullAdder_740_io_b = FullAdder_638_io_s; // @[wallace.scala 70:18]
  assign FullAdder_740_io_ci = FullAdder_639_io_co; // @[wallace.scala 71:19]
  assign FullAdder_741_io_a = FullAdder_639_io_s; // @[wallace.scala 69:18]
  assign FullAdder_741_io_b = FullAdder_640_io_s; // @[wallace.scala 70:18]
  assign FullAdder_741_io_ci = FullAdder_641_io_s; // @[wallace.scala 71:19]
  assign FullAdder_742_io_a = FullAdder_642_io_co; // @[wallace.scala 69:18]
  assign FullAdder_742_io_b = FullAdder_643_io_co; // @[wallace.scala 70:18]
  assign FullAdder_742_io_ci = FullAdder_644_io_co; // @[wallace.scala 71:19]
  assign FullAdder_743_io_a = FullAdder_642_io_s; // @[wallace.scala 69:18]
  assign FullAdder_743_io_b = FullAdder_643_io_s; // @[wallace.scala 70:18]
  assign FullAdder_743_io_ci = FullAdder_644_io_s; // @[wallace.scala 71:19]
  assign FullAdder_744_io_a = FullAdder_645_io_co; // @[wallace.scala 69:18]
  assign FullAdder_744_io_b = FullAdder_646_io_co; // @[wallace.scala 70:18]
  assign FullAdder_744_io_ci = FullAdder_647_io_co; // @[wallace.scala 71:19]
  assign FullAdder_745_io_a = FullAdder_498_io_co; // @[wallace.scala 69:18]
  assign FullAdder_745_io_b = FullAdder_645_io_s; // @[wallace.scala 70:18]
  assign FullAdder_745_io_ci = FullAdder_646_io_s; // @[wallace.scala 71:19]
  assign FullAdder_746_io_a = FullAdder_647_io_s; // @[wallace.scala 69:18]
  assign FullAdder_746_io_b = FullAdder_648_io_co; // @[wallace.scala 70:18]
  assign FullAdder_746_io_ci = FullAdder_649_io_co; // @[wallace.scala 71:19]
  assign FullAdder_747_io_a = FullAdder_648_io_s; // @[wallace.scala 69:18]
  assign FullAdder_747_io_b = FullAdder_649_io_s; // @[wallace.scala 70:18]
  assign FullAdder_747_io_ci = FullAdder_650_io_s; // @[wallace.scala 71:19]
  assign FullAdder_748_io_a = FullAdder_651_io_co; // @[wallace.scala 69:18]
  assign FullAdder_748_io_b = FullAdder_652_io_co; // @[wallace.scala 70:18]
  assign FullAdder_748_io_ci = HalfAdder_47_io_co; // @[wallace.scala 71:19]
  assign FullAdder_749_io_a = FullAdder_651_io_s; // @[wallace.scala 69:18]
  assign FullAdder_749_io_b = FullAdder_652_io_s; // @[wallace.scala 70:18]
  assign FullAdder_749_io_ci = HalfAdder_47_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_66_io_a = FullAdder_653_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_66_io_b = FullAdder_654_io_co; // @[wallace.scala 60:18]
  assign FullAdder_750_io_a = FullAdder_508_io_co; // @[wallace.scala 69:18]
  assign FullAdder_750_io_b = FullAdder_653_io_s; // @[wallace.scala 70:18]
  assign FullAdder_750_io_ci = FullAdder_654_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_67_io_a = FullAdder_655_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_67_io_b = FullAdder_656_io_co; // @[wallace.scala 60:18]
  assign FullAdder_751_io_a = FullAdder_510_io_co; // @[wallace.scala 69:18]
  assign FullAdder_751_io_b = FullAdder_511_io_co; // @[wallace.scala 70:18]
  assign FullAdder_751_io_ci = FullAdder_655_io_s; // @[wallace.scala 71:19]
  assign FullAdder_752_io_a = FullAdder_656_io_s; // @[wallace.scala 69:18]
  assign FullAdder_752_io_b = FullAdder_657_io_co; // @[wallace.scala 70:18]
  assign FullAdder_752_io_ci = FullAdder_658_io_co; // @[wallace.scala 71:19]
  assign FullAdder_753_io_a = FullAdder_657_io_s; // @[wallace.scala 69:18]
  assign FullAdder_753_io_b = FullAdder_658_io_s; // @[wallace.scala 70:18]
  assign FullAdder_753_io_ci = FullAdder_659_io_co; // @[wallace.scala 71:19]
  assign FullAdder_754_io_a = FullAdder_517_io_co; // @[wallace.scala 69:18]
  assign FullAdder_754_io_b = FullAdder_659_io_s; // @[wallace.scala 70:18]
  assign FullAdder_754_io_ci = FullAdder_660_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_68_io_a = FullAdder_661_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_68_io_b = FullAdder_662_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_69_io_a = FullAdder_663_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_69_io_b = HalfAdder_48_io_co; // @[wallace.scala 60:18]
  assign FullAdder_755_io_a = FullAdder_663_io_s; // @[wallace.scala 69:18]
  assign FullAdder_755_io_b = HalfAdder_48_io_s; // @[wallace.scala 70:18]
  assign FullAdder_755_io_ci = FullAdder_664_io_co; // @[wallace.scala 71:19]
  assign FullAdder_756_io_a = FullAdder_664_io_s; // @[wallace.scala 69:18]
  assign FullAdder_756_io_b = HalfAdder_49_io_s; // @[wallace.scala 70:18]
  assign FullAdder_756_io_ci = FullAdder_665_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_70_io_a = FullAdder_665_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_70_io_b = HalfAdder_50_io_s; // @[wallace.scala 60:18]
  assign FullAdder_757_io_a = HalfAdder_29_io_co; // @[wallace.scala 69:18]
  assign FullAdder_757_io_b = FullAdder_666_io_s; // @[wallace.scala 70:18]
  assign FullAdder_757_io_ci = FullAdder_667_io_co; // @[wallace.scala 71:19]
  assign FullAdder_758_io_a = HalfAdder_30_io_co; // @[wallace.scala 69:18]
  assign FullAdder_758_io_b = FullAdder_667_io_s; // @[wallace.scala 70:18]
  assign FullAdder_758_io_ci = FullAdder_668_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_71_io_a = HalfAdder_32_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_71_io_b = FullAdder_668_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_72_io_a = HalfAdder_33_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_72_io_b = HalfAdder_51_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_73_io_a = HalfAdder_53_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_73_io_b = HalfAdder_54_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_74_io_a = HalfAdder_54_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_74_io_b = HalfAdder_55_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_75_io_a = FullAdder_529_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_75_io_b = HalfAdder_55_io_s; // @[wallace.scala 60:18]
  assign FullAdder_759_io_a = FullAdder_530_io_s; // @[wallace.scala 69:18]
  assign FullAdder_759_io_b = FullAdder_531_io_co; // @[wallace.scala 70:18]
  assign FullAdder_759_io_ci = FullAdder_669_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_76_io_a = FullAdder_669_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_76_io_b = FullAdder_670_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_77_io_a = FullAdder_670_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_77_io_b = FullAdder_671_io_co; // @[wallace.scala 60:18]
  assign FullAdder_760_io_a = FullAdder_534_io_co; // @[wallace.scala 69:18]
  assign FullAdder_760_io_b = HalfAdder_37_io_co; // @[wallace.scala 70:18]
  assign FullAdder_760_io_ci = FullAdder_671_io_s; // @[wallace.scala 71:19]
  assign FullAdder_761_io_a = FullAdder_536_io_co; // @[wallace.scala 69:18]
  assign FullAdder_761_io_b = FullAdder_672_io_s; // @[wallace.scala 70:18]
  assign FullAdder_761_io_ci = FullAdder_673_io_co; // @[wallace.scala 71:19]
  assign FullAdder_762_io_a = FullAdder_538_io_co; // @[wallace.scala 69:18]
  assign FullAdder_762_io_b = FullAdder_673_io_s; // @[wallace.scala 70:18]
  assign FullAdder_762_io_ci = FullAdder_674_io_co; // @[wallace.scala 71:19]
  assign FullAdder_763_io_a = FullAdder_540_io_co; // @[wallace.scala 69:18]
  assign FullAdder_763_io_b = FullAdder_674_io_s; // @[wallace.scala 70:18]
  assign FullAdder_763_io_ci = FullAdder_675_io_co; // @[wallace.scala 71:19]
  assign FullAdder_764_io_a = FullAdder_542_io_co; // @[wallace.scala 69:18]
  assign FullAdder_764_io_b = FullAdder_675_io_s; // @[wallace.scala 70:18]
  assign FullAdder_764_io_ci = FullAdder_676_io_co; // @[wallace.scala 71:19]
  assign FullAdder_765_io_a = FullAdder_676_io_s; // @[wallace.scala 69:18]
  assign FullAdder_765_io_b = HalfAdder_57_io_s; // @[wallace.scala 70:18]
  assign FullAdder_765_io_ci = HalfAdder_58_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_78_io_a = HalfAdder_59_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_78_io_b = HalfAdder_60_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_79_io_a = HalfAdder_58_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_79_io_b = HalfAdder_59_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_80_io_a = HalfAdder_60_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_80_io_b = FullAdder_677_io_co; // @[wallace.scala 60:18]
  assign FullAdder_766_io_a = FullAdder_677_io_s; // @[wallace.scala 69:18]
  assign FullAdder_766_io_b = FullAdder_678_io_s; // @[wallace.scala 70:18]
  assign FullAdder_766_io_ci = FullAdder_679_io_co; // @[wallace.scala 71:19]
  assign FullAdder_767_io_a = FullAdder_679_io_s; // @[wallace.scala 69:18]
  assign FullAdder_767_io_b = FullAdder_680_io_s; // @[wallace.scala 70:18]
  assign FullAdder_767_io_ci = FullAdder_681_io_co; // @[wallace.scala 71:19]
  assign FullAdder_768_io_a = FullAdder_681_io_s; // @[wallace.scala 69:18]
  assign FullAdder_768_io_b = FullAdder_682_io_s; // @[wallace.scala 70:18]
  assign FullAdder_768_io_ci = FullAdder_683_io_co; // @[wallace.scala 71:19]
  assign FullAdder_769_io_a = FullAdder_683_io_s; // @[wallace.scala 69:18]
  assign FullAdder_769_io_b = FullAdder_684_io_s; // @[wallace.scala 70:18]
  assign FullAdder_769_io_ci = FullAdder_685_io_co; // @[wallace.scala 71:19]
  assign FullAdder_770_io_a = FullAdder_558_io_co; // @[wallace.scala 69:18]
  assign FullAdder_770_io_b = FullAdder_685_io_s; // @[wallace.scala 70:18]
  assign FullAdder_770_io_ci = FullAdder_686_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_81_io_a = FullAdder_687_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_81_io_b = FullAdder_688_io_co; // @[wallace.scala 60:18]
  assign FullAdder_771_io_a = FullAdder_561_io_co; // @[wallace.scala 69:18]
  assign FullAdder_771_io_b = FullAdder_687_io_s; // @[wallace.scala 70:18]
  assign FullAdder_771_io_ci = FullAdder_688_io_s; // @[wallace.scala 71:19]
  assign FullAdder_772_io_a = FullAdder_564_io_co; // @[wallace.scala 69:18]
  assign FullAdder_772_io_b = HalfAdder_42_io_co; // @[wallace.scala 70:18]
  assign FullAdder_772_io_ci = FullAdder_689_io_s; // @[wallace.scala 71:19]
  assign FullAdder_773_io_a = FullAdder_690_io_s; // @[wallace.scala 69:18]
  assign FullAdder_773_io_b = FullAdder_691_io_co; // @[wallace.scala 70:18]
  assign FullAdder_773_io_ci = HalfAdder_61_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_82_io_a = HalfAdder_43_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_82_io_b = FullAdder_691_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_83_io_a = HalfAdder_61_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_83_io_b = HalfAdder_62_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_84_io_a = FullAdder_692_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_84_io_b = FullAdder_693_io_co; // @[wallace.scala 60:18]
  assign FullAdder_774_io_a = FullAdder_570_io_co; // @[wallace.scala 69:18]
  assign FullAdder_774_io_b = FullAdder_571_io_co; // @[wallace.scala 70:18]
  assign FullAdder_774_io_ci = FullAdder_692_io_s; // @[wallace.scala 71:19]
  assign FullAdder_775_io_a = FullAdder_693_io_s; // @[wallace.scala 69:18]
  assign FullAdder_775_io_b = FullAdder_694_io_co; // @[wallace.scala 70:18]
  assign FullAdder_775_io_ci = FullAdder_695_io_co; // @[wallace.scala 71:19]
  assign FullAdder_776_io_a = FullAdder_694_io_s; // @[wallace.scala 69:18]
  assign FullAdder_776_io_b = FullAdder_695_io_s; // @[wallace.scala 70:18]
  assign FullAdder_776_io_ci = HalfAdder_63_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_85_io_a = FullAdder_696_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_85_io_b = FullAdder_697_io_co; // @[wallace.scala 60:18]
  assign FullAdder_777_io_a = FullAdder_578_io_co; // @[wallace.scala 69:18]
  assign FullAdder_777_io_b = FullAdder_579_io_co; // @[wallace.scala 70:18]
  assign FullAdder_777_io_ci = FullAdder_696_io_s; // @[wallace.scala 71:19]
  assign FullAdder_778_io_a = FullAdder_697_io_s; // @[wallace.scala 69:18]
  assign FullAdder_778_io_b = FullAdder_698_io_co; // @[wallace.scala 70:18]
  assign FullAdder_778_io_ci = FullAdder_699_io_co; // @[wallace.scala 71:19]
  assign FullAdder_779_io_a = FullAdder_698_io_s; // @[wallace.scala 69:18]
  assign FullAdder_779_io_b = FullAdder_699_io_s; // @[wallace.scala 70:18]
  assign FullAdder_779_io_ci = FullAdder_700_io_s; // @[wallace.scala 71:19]
  assign FullAdder_780_io_a = FullAdder_701_io_co; // @[wallace.scala 69:18]
  assign FullAdder_780_io_b = FullAdder_702_io_co; // @[wallace.scala 70:18]
  assign FullAdder_780_io_ci = FullAdder_703_io_co; // @[wallace.scala 71:19]
  assign FullAdder_781_io_a = HalfAdder_44_io_co; // @[wallace.scala 69:18]
  assign FullAdder_781_io_b = FullAdder_701_io_s; // @[wallace.scala 70:18]
  assign FullAdder_781_io_ci = FullAdder_702_io_s; // @[wallace.scala 71:19]
  assign FullAdder_782_io_a = FullAdder_703_io_s; // @[wallace.scala 69:18]
  assign FullAdder_782_io_b = FullAdder_704_io_co; // @[wallace.scala 70:18]
  assign FullAdder_782_io_ci = FullAdder_705_io_co; // @[wallace.scala 71:19]
  assign FullAdder_783_io_a = FullAdder_704_io_s; // @[wallace.scala 69:18]
  assign FullAdder_783_io_b = FullAdder_705_io_s; // @[wallace.scala 70:18]
  assign FullAdder_783_io_ci = FullAdder_706_io_s; // @[wallace.scala 71:19]
  assign FullAdder_784_io_a = FullAdder_707_io_co; // @[wallace.scala 69:18]
  assign FullAdder_784_io_b = FullAdder_708_io_co; // @[wallace.scala 70:18]
  assign FullAdder_784_io_ci = FullAdder_709_io_co; // @[wallace.scala 71:19]
  assign FullAdder_785_io_a = FullAdder_596_io_co; // @[wallace.scala 69:18]
  assign FullAdder_785_io_b = FullAdder_707_io_s; // @[wallace.scala 70:18]
  assign FullAdder_785_io_ci = FullAdder_708_io_s; // @[wallace.scala 71:19]
  assign FullAdder_786_io_a = FullAdder_709_io_s; // @[wallace.scala 69:18]
  assign FullAdder_786_io_b = FullAdder_710_io_co; // @[wallace.scala 70:18]
  assign FullAdder_786_io_ci = FullAdder_711_io_co; // @[wallace.scala 71:19]
  assign FullAdder_787_io_a = HalfAdder_45_io_co; // @[wallace.scala 69:18]
  assign FullAdder_787_io_b = FullAdder_710_io_s; // @[wallace.scala 70:18]
  assign FullAdder_787_io_ci = FullAdder_711_io_s; // @[wallace.scala 71:19]
  assign FullAdder_788_io_a = FullAdder_712_io_s; // @[wallace.scala 69:18]
  assign FullAdder_788_io_b = FullAdder_713_io_co; // @[wallace.scala 70:18]
  assign FullAdder_788_io_ci = FullAdder_714_io_co; // @[wallace.scala 71:19]
  assign FullAdder_789_io_a = FullAdder_605_io_co; // @[wallace.scala 69:18]
  assign FullAdder_789_io_b = FullAdder_713_io_s; // @[wallace.scala 70:18]
  assign FullAdder_789_io_ci = FullAdder_714_io_s; // @[wallace.scala 71:19]
  assign FullAdder_790_io_a = FullAdder_715_io_s; // @[wallace.scala 69:18]
  assign FullAdder_790_io_b = FullAdder_716_io_co; // @[wallace.scala 70:18]
  assign FullAdder_790_io_ci = FullAdder_717_io_co; // @[wallace.scala 71:19]
  assign FullAdder_791_io_a = FullAdder_716_io_s; // @[wallace.scala 69:18]
  assign FullAdder_791_io_b = FullAdder_717_io_s; // @[wallace.scala 70:18]
  assign FullAdder_791_io_ci = FullAdder_718_io_s; // @[wallace.scala 71:19]
  assign FullAdder_792_io_a = FullAdder_719_io_co; // @[wallace.scala 69:18]
  assign FullAdder_792_io_b = FullAdder_720_io_co; // @[wallace.scala 70:18]
  assign FullAdder_792_io_ci = FullAdder_721_io_co; // @[wallace.scala 71:19]
  assign FullAdder_793_io_a = FullAdder_719_io_s; // @[wallace.scala 69:18]
  assign FullAdder_793_io_b = FullAdder_720_io_s; // @[wallace.scala 70:18]
  assign FullAdder_793_io_ci = FullAdder_721_io_s; // @[wallace.scala 71:19]
  assign FullAdder_794_io_a = FullAdder_722_io_co; // @[wallace.scala 69:18]
  assign FullAdder_794_io_b = FullAdder_723_io_co; // @[wallace.scala 70:18]
  assign FullAdder_794_io_ci = FullAdder_724_io_co; // @[wallace.scala 71:19]
  assign FullAdder_795_io_a = FullAdder_617_io_co; // @[wallace.scala 69:18]
  assign FullAdder_795_io_b = FullAdder_722_io_s; // @[wallace.scala 70:18]
  assign FullAdder_795_io_ci = FullAdder_723_io_s; // @[wallace.scala 71:19]
  assign FullAdder_796_io_a = FullAdder_724_io_s; // @[wallace.scala 69:18]
  assign FullAdder_796_io_b = FullAdder_725_io_co; // @[wallace.scala 70:18]
  assign FullAdder_796_io_ci = FullAdder_726_io_co; // @[wallace.scala 71:19]
  assign FullAdder_797_io_a = FullAdder_725_io_s; // @[wallace.scala 69:18]
  assign FullAdder_797_io_b = FullAdder_726_io_s; // @[wallace.scala 70:18]
  assign FullAdder_797_io_ci = FullAdder_727_io_s; // @[wallace.scala 71:19]
  assign FullAdder_798_io_a = FullAdder_728_io_co; // @[wallace.scala 69:18]
  assign FullAdder_798_io_b = FullAdder_729_io_co; // @[wallace.scala 70:18]
  assign FullAdder_798_io_ci = FullAdder_730_io_co; // @[wallace.scala 71:19]
  assign FullAdder_799_io_a = FullAdder_728_io_s; // @[wallace.scala 69:18]
  assign FullAdder_799_io_b = FullAdder_729_io_s; // @[wallace.scala 70:18]
  assign FullAdder_799_io_ci = FullAdder_730_io_s; // @[wallace.scala 71:19]
  assign FullAdder_800_io_a = FullAdder_731_io_co; // @[wallace.scala 69:18]
  assign FullAdder_800_io_b = FullAdder_732_io_co; // @[wallace.scala 70:18]
  assign FullAdder_800_io_ci = HalfAdder_64_io_co; // @[wallace.scala 71:19]
  assign FullAdder_801_io_a = FullAdder_731_io_s; // @[wallace.scala 69:18]
  assign FullAdder_801_io_b = FullAdder_732_io_s; // @[wallace.scala 70:18]
  assign FullAdder_801_io_ci = HalfAdder_64_io_s; // @[wallace.scala 71:19]
  assign FullAdder_802_io_a = FullAdder_733_io_co; // @[wallace.scala 69:18]
  assign FullAdder_802_io_b = FullAdder_734_io_co; // @[wallace.scala 70:18]
  assign FullAdder_802_io_ci = HalfAdder_65_io_co; // @[wallace.scala 71:19]
  assign FullAdder_803_io_a = FullAdder_733_io_s; // @[wallace.scala 69:18]
  assign FullAdder_803_io_b = FullAdder_734_io_s; // @[wallace.scala 70:18]
  assign FullAdder_803_io_ci = HalfAdder_65_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_86_io_a = FullAdder_735_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_86_io_b = FullAdder_736_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_87_io_a = FullAdder_635_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_87_io_b = FullAdder_735_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_88_io_a = FullAdder_736_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_88_io_b = FullAdder_737_io_co; // @[wallace.scala 60:18]
  assign FullAdder_804_io_a = FullAdder_638_io_co; // @[wallace.scala 69:18]
  assign FullAdder_804_io_b = FullAdder_737_io_s; // @[wallace.scala 70:18]
  assign FullAdder_804_io_ci = FullAdder_738_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_89_io_a = FullAdder_739_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_89_io_b = FullAdder_740_io_co; // @[wallace.scala 60:18]
  assign FullAdder_805_io_a = FullAdder_640_io_co; // @[wallace.scala 69:18]
  assign FullAdder_805_io_b = FullAdder_641_io_co; // @[wallace.scala 70:18]
  assign FullAdder_805_io_ci = FullAdder_739_io_s; // @[wallace.scala 71:19]
  assign FullAdder_806_io_a = FullAdder_740_io_s; // @[wallace.scala 69:18]
  assign FullAdder_806_io_b = FullAdder_741_io_co; // @[wallace.scala 70:18]
  assign FullAdder_806_io_ci = FullAdder_742_io_co; // @[wallace.scala 71:19]
  assign FullAdder_807_io_a = FullAdder_741_io_s; // @[wallace.scala 69:18]
  assign FullAdder_807_io_b = FullAdder_742_io_s; // @[wallace.scala 70:18]
  assign FullAdder_807_io_ci = FullAdder_743_io_co; // @[wallace.scala 71:19]
  assign FullAdder_808_io_a = FullAdder_743_io_s; // @[wallace.scala 69:18]
  assign FullAdder_808_io_b = FullAdder_744_io_s; // @[wallace.scala 70:18]
  assign FullAdder_808_io_ci = FullAdder_745_io_co; // @[wallace.scala 71:19]
  assign FullAdder_809_io_a = FullAdder_650_io_co; // @[wallace.scala 69:18]
  assign FullAdder_809_io_b = FullAdder_745_io_s; // @[wallace.scala 70:18]
  assign FullAdder_809_io_ci = FullAdder_746_io_s; // @[wallace.scala 71:19]
  assign FullAdder_810_io_a = FullAdder_747_io_s; // @[wallace.scala 69:18]
  assign FullAdder_810_io_b = FullAdder_748_io_s; // @[wallace.scala 70:18]
  assign FullAdder_810_io_ci = FullAdder_749_io_co; // @[wallace.scala 71:19]
  assign FullAdder_811_io_a = FullAdder_749_io_s; // @[wallace.scala 69:18]
  assign FullAdder_811_io_b = HalfAdder_66_io_s; // @[wallace.scala 70:18]
  assign FullAdder_811_io_ci = FullAdder_750_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_90_io_a = FullAdder_750_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_90_io_b = HalfAdder_67_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_91_io_a = FullAdder_751_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_91_io_b = FullAdder_752_io_co; // @[wallace.scala 60:18]
  assign FullAdder_812_io_a = FullAdder_751_io_s; // @[wallace.scala 69:18]
  assign FullAdder_812_io_b = FullAdder_752_io_s; // @[wallace.scala 70:18]
  assign FullAdder_812_io_ci = FullAdder_753_io_co; // @[wallace.scala 71:19]
  assign FullAdder_813_io_a = FullAdder_660_io_co; // @[wallace.scala 69:18]
  assign FullAdder_813_io_b = FullAdder_753_io_s; // @[wallace.scala 70:18]
  assign FullAdder_813_io_ci = FullAdder_754_io_co; // @[wallace.scala 71:19]
  assign FullAdder_814_io_a = FullAdder_661_io_co; // @[wallace.scala 69:18]
  assign FullAdder_814_io_b = FullAdder_662_io_co; // @[wallace.scala 70:18]
  assign FullAdder_814_io_ci = FullAdder_754_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_92_io_a = HalfAdder_68_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_92_io_b = HalfAdder_69_io_s; // @[wallace.scala 60:18]
  assign FullAdder_815_io_a = HalfAdder_49_io_co; // @[wallace.scala 69:18]
  assign FullAdder_815_io_b = FullAdder_755_io_s; // @[wallace.scala 70:18]
  assign FullAdder_815_io_ci = FullAdder_756_io_co; // @[wallace.scala 71:19]
  assign FullAdder_816_io_a = HalfAdder_50_io_co; // @[wallace.scala 69:18]
  assign FullAdder_816_io_b = FullAdder_756_io_s; // @[wallace.scala 70:18]
  assign FullAdder_816_io_ci = HalfAdder_70_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_93_io_a = FullAdder_666_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_93_io_b = HalfAdder_70_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_94_io_a = FullAdder_757_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_94_io_b = FullAdder_758_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_95_io_a = HalfAdder_51_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_95_io_b = HalfAdder_71_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_96_io_a = HalfAdder_52_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_96_io_b = HalfAdder_72_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_97_io_a = HalfAdder_73_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_97_io_b = HalfAdder_74_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_98_io_a = HalfAdder_56_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_98_io_b = HalfAdder_75_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_99_io_a = HalfAdder_56_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_99_io_b = FullAdder_759_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_100_io_a = HalfAdder_76_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_100_io_b = HalfAdder_77_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_101_io_a = HalfAdder_77_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_101_io_b = FullAdder_760_io_co; // @[wallace.scala 60:18]
  assign FullAdder_817_io_a = FullAdder_672_io_co; // @[wallace.scala 69:18]
  assign FullAdder_817_io_b = FullAdder_760_io_s; // @[wallace.scala 70:18]
  assign FullAdder_817_io_ci = FullAdder_761_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_102_io_a = FullAdder_761_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_102_io_b = FullAdder_762_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_103_io_a = FullAdder_762_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_103_io_b = FullAdder_763_io_co; // @[wallace.scala 60:18]
  assign FullAdder_818_io_a = HalfAdder_57_io_co; // @[wallace.scala 69:18]
  assign FullAdder_818_io_b = FullAdder_764_io_s; // @[wallace.scala 70:18]
  assign FullAdder_818_io_ci = FullAdder_765_io_co; // @[wallace.scala 71:19]
  assign FullAdder_819_io_a = FullAdder_765_io_s; // @[wallace.scala 69:18]
  assign FullAdder_819_io_b = HalfAdder_78_io_s; // @[wallace.scala 70:18]
  assign FullAdder_819_io_ci = HalfAdder_79_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_104_io_a = FullAdder_678_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_104_io_b = HalfAdder_79_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_105_io_a = HalfAdder_80_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_105_io_b = FullAdder_766_io_co; // @[wallace.scala 60:18]
  assign FullAdder_820_io_a = FullAdder_680_io_co; // @[wallace.scala 69:18]
  assign FullAdder_820_io_b = FullAdder_766_io_s; // @[wallace.scala 70:18]
  assign FullAdder_820_io_ci = FullAdder_767_io_co; // @[wallace.scala 71:19]
  assign FullAdder_821_io_a = FullAdder_682_io_co; // @[wallace.scala 69:18]
  assign FullAdder_821_io_b = FullAdder_767_io_s; // @[wallace.scala 70:18]
  assign FullAdder_821_io_ci = FullAdder_768_io_co; // @[wallace.scala 71:19]
  assign FullAdder_822_io_a = FullAdder_684_io_co; // @[wallace.scala 69:18]
  assign FullAdder_822_io_b = FullAdder_768_io_s; // @[wallace.scala 70:18]
  assign FullAdder_822_io_ci = FullAdder_769_io_co; // @[wallace.scala 71:19]
  assign FullAdder_823_io_a = FullAdder_686_io_co; // @[wallace.scala 69:18]
  assign FullAdder_823_io_b = FullAdder_769_io_s; // @[wallace.scala 70:18]
  assign FullAdder_823_io_ci = FullAdder_770_io_co; // @[wallace.scala 71:19]
  assign FullAdder_824_io_a = FullAdder_770_io_s; // @[wallace.scala 69:18]
  assign FullAdder_824_io_b = HalfAdder_81_io_s; // @[wallace.scala 70:18]
  assign FullAdder_824_io_ci = FullAdder_771_io_co; // @[wallace.scala 71:19]
  assign FullAdder_825_io_a = FullAdder_689_io_co; // @[wallace.scala 69:18]
  assign FullAdder_825_io_b = FullAdder_690_io_co; // @[wallace.scala 70:18]
  assign FullAdder_825_io_ci = FullAdder_771_io_s; // @[wallace.scala 71:19]
  assign FullAdder_826_io_a = HalfAdder_62_io_co; // @[wallace.scala 69:18]
  assign FullAdder_826_io_b = FullAdder_772_io_s; // @[wallace.scala 70:18]
  assign FullAdder_826_io_ci = FullAdder_773_io_s; // @[wallace.scala 71:19]
  assign FullAdder_827_io_a = HalfAdder_82_io_co; // @[wallace.scala 69:18]
  assign FullAdder_827_io_b = HalfAdder_83_io_co; // @[wallace.scala 70:18]
  assign FullAdder_827_io_ci = HalfAdder_84_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_106_io_a = HalfAdder_82_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_106_io_b = HalfAdder_83_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_107_io_a = HalfAdder_84_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_107_io_b = FullAdder_774_io_co; // @[wallace.scala 60:18]
  assign FullAdder_828_io_a = HalfAdder_63_io_co; // @[wallace.scala 69:18]
  assign FullAdder_828_io_b = FullAdder_774_io_s; // @[wallace.scala 70:18]
  assign FullAdder_828_io_ci = FullAdder_775_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_108_io_a = FullAdder_776_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_108_io_b = HalfAdder_85_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_109_io_a = FullAdder_777_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_109_io_b = FullAdder_778_io_co; // @[wallace.scala 60:18]
  assign FullAdder_829_io_a = FullAdder_700_io_co; // @[wallace.scala 69:18]
  assign FullAdder_829_io_b = FullAdder_777_io_s; // @[wallace.scala 70:18]
  assign FullAdder_829_io_ci = FullAdder_778_io_s; // @[wallace.scala 71:19]
  assign FullAdder_830_io_a = FullAdder_779_io_s; // @[wallace.scala 69:18]
  assign FullAdder_830_io_b = FullAdder_780_io_s; // @[wallace.scala 70:18]
  assign FullAdder_830_io_ci = FullAdder_781_io_co; // @[wallace.scala 71:19]
  assign FullAdder_831_io_a = FullAdder_706_io_co; // @[wallace.scala 69:18]
  assign FullAdder_831_io_b = FullAdder_781_io_s; // @[wallace.scala 70:18]
  assign FullAdder_831_io_ci = FullAdder_782_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_110_io_a = FullAdder_783_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_110_io_b = FullAdder_784_io_co; // @[wallace.scala 60:18]
  assign FullAdder_832_io_a = FullAdder_783_io_s; // @[wallace.scala 69:18]
  assign FullAdder_832_io_b = FullAdder_784_io_s; // @[wallace.scala 70:18]
  assign FullAdder_832_io_ci = FullAdder_785_io_co; // @[wallace.scala 71:19]
  assign FullAdder_833_io_a = FullAdder_712_io_co; // @[wallace.scala 69:18]
  assign FullAdder_833_io_b = FullAdder_785_io_s; // @[wallace.scala 70:18]
  assign FullAdder_833_io_ci = FullAdder_786_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_111_io_a = FullAdder_787_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_111_io_b = FullAdder_788_io_co; // @[wallace.scala 60:18]
  assign FullAdder_834_io_a = FullAdder_715_io_co; // @[wallace.scala 69:18]
  assign FullAdder_834_io_b = FullAdder_787_io_s; // @[wallace.scala 70:18]
  assign FullAdder_834_io_ci = FullAdder_788_io_s; // @[wallace.scala 71:19]
  assign FullAdder_835_io_a = FullAdder_718_io_co; // @[wallace.scala 69:18]
  assign FullAdder_835_io_b = FullAdder_789_io_s; // @[wallace.scala 70:18]
  assign FullAdder_835_io_ci = FullAdder_790_io_s; // @[wallace.scala 71:19]
  assign FullAdder_836_io_a = FullAdder_791_io_s; // @[wallace.scala 69:18]
  assign FullAdder_836_io_b = FullAdder_792_io_s; // @[wallace.scala 70:18]
  assign FullAdder_836_io_ci = FullAdder_793_io_co; // @[wallace.scala 71:19]
  assign FullAdder_837_io_a = FullAdder_793_io_s; // @[wallace.scala 69:18]
  assign FullAdder_837_io_b = FullAdder_794_io_s; // @[wallace.scala 70:18]
  assign FullAdder_837_io_ci = FullAdder_795_io_co; // @[wallace.scala 71:19]
  assign FullAdder_838_io_a = FullAdder_727_io_co; // @[wallace.scala 69:18]
  assign FullAdder_838_io_b = FullAdder_795_io_s; // @[wallace.scala 70:18]
  assign FullAdder_838_io_ci = FullAdder_796_io_s; // @[wallace.scala 71:19]
  assign FullAdder_839_io_a = FullAdder_797_io_s; // @[wallace.scala 69:18]
  assign FullAdder_839_io_b = FullAdder_798_io_s; // @[wallace.scala 70:18]
  assign FullAdder_839_io_ci = FullAdder_799_io_co; // @[wallace.scala 71:19]
  assign FullAdder_840_io_a = FullAdder_799_io_s; // @[wallace.scala 69:18]
  assign FullAdder_840_io_b = FullAdder_800_io_s; // @[wallace.scala 70:18]
  assign FullAdder_840_io_ci = FullAdder_801_io_co; // @[wallace.scala 71:19]
  assign FullAdder_841_io_a = FullAdder_801_io_s; // @[wallace.scala 69:18]
  assign FullAdder_841_io_b = FullAdder_802_io_s; // @[wallace.scala 70:18]
  assign FullAdder_841_io_ci = FullAdder_803_io_co; // @[wallace.scala 71:19]
  assign FullAdder_842_io_a = FullAdder_803_io_s; // @[wallace.scala 69:18]
  assign FullAdder_842_io_b = HalfAdder_86_io_s; // @[wallace.scala 70:18]
  assign FullAdder_842_io_ci = HalfAdder_87_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_112_io_a = FullAdder_738_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_112_io_b = HalfAdder_87_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_113_io_a = HalfAdder_88_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_113_io_b = FullAdder_804_io_co; // @[wallace.scala 60:18]
  assign FullAdder_843_io_a = FullAdder_804_io_s; // @[wallace.scala 69:18]
  assign FullAdder_843_io_b = HalfAdder_89_io_s; // @[wallace.scala 70:18]
  assign FullAdder_843_io_ci = FullAdder_805_io_co; // @[wallace.scala 71:19]
  assign FullAdder_844_io_a = FullAdder_805_io_s; // @[wallace.scala 69:18]
  assign FullAdder_844_io_b = FullAdder_806_io_s; // @[wallace.scala 70:18]
  assign FullAdder_844_io_ci = FullAdder_807_io_co; // @[wallace.scala 71:19]
  assign FullAdder_845_io_a = FullAdder_744_io_co; // @[wallace.scala 69:18]
  assign FullAdder_845_io_b = FullAdder_807_io_s; // @[wallace.scala 70:18]
  assign FullAdder_845_io_ci = FullAdder_808_io_co; // @[wallace.scala 71:19]
  assign FullAdder_846_io_a = FullAdder_746_io_co; // @[wallace.scala 69:18]
  assign FullAdder_846_io_b = FullAdder_808_io_s; // @[wallace.scala 70:18]
  assign FullAdder_846_io_ci = FullAdder_809_io_co; // @[wallace.scala 71:19]
  assign FullAdder_847_io_a = FullAdder_747_io_co; // @[wallace.scala 69:18]
  assign FullAdder_847_io_b = FullAdder_748_io_co; // @[wallace.scala 70:18]
  assign FullAdder_847_io_ci = FullAdder_809_io_s; // @[wallace.scala 71:19]
  assign FullAdder_848_io_a = HalfAdder_66_io_co; // @[wallace.scala 69:18]
  assign FullAdder_848_io_b = FullAdder_810_io_s; // @[wallace.scala 70:18]
  assign FullAdder_848_io_ci = FullAdder_811_io_co; // @[wallace.scala 71:19]
  assign FullAdder_849_io_a = HalfAdder_67_io_co; // @[wallace.scala 69:18]
  assign FullAdder_849_io_b = FullAdder_811_io_s; // @[wallace.scala 70:18]
  assign FullAdder_849_io_ci = HalfAdder_90_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_114_io_a = HalfAdder_90_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_114_io_b = HalfAdder_91_io_s; // @[wallace.scala 60:18]
  assign FullAdder_850_io_a = HalfAdder_68_io_co; // @[wallace.scala 69:18]
  assign FullAdder_850_io_b = HalfAdder_69_io_co; // @[wallace.scala 70:18]
  assign FullAdder_850_io_ci = FullAdder_814_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_115_io_a = FullAdder_755_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_115_io_b = HalfAdder_92_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_116_io_a = FullAdder_816_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_116_io_b = HalfAdder_93_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_117_io_a = FullAdder_757_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_117_io_b = HalfAdder_93_io_s; // @[wallace.scala 60:18]
  assign FullAdder_851_io_a = FullAdder_758_io_s; // @[wallace.scala 69:18]
  assign FullAdder_851_io_b = HalfAdder_71_io_co; // @[wallace.scala 70:18]
  assign FullAdder_851_io_ci = HalfAdder_95_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_118_io_a = HalfAdder_72_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_118_io_b = HalfAdder_95_io_s; // @[wallace.scala 60:18]
  assign FullAdder_852_io_a = HalfAdder_74_io_s; // @[wallace.scala 69:18]
  assign FullAdder_852_io_b = HalfAdder_75_io_co; // @[wallace.scala 70:18]
  assign FullAdder_852_io_ci = HalfAdder_98_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_119_io_a = HalfAdder_98_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_119_io_b = HalfAdder_99_io_co; // @[wallace.scala 60:18]
  assign FullAdder_853_io_a = FullAdder_759_io_s; // @[wallace.scala 69:18]
  assign FullAdder_853_io_b = HalfAdder_76_io_co; // @[wallace.scala 70:18]
  assign FullAdder_853_io_ci = HalfAdder_100_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_120_io_a = HalfAdder_100_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_120_io_b = HalfAdder_101_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_121_io_a = HalfAdder_101_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_121_io_b = FullAdder_817_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_122_io_a = HalfAdder_102_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_122_io_b = HalfAdder_103_io_co; // @[wallace.scala 60:18]
  assign FullAdder_854_io_a = FullAdder_763_io_s; // @[wallace.scala 69:18]
  assign FullAdder_854_io_b = FullAdder_764_io_co; // @[wallace.scala 70:18]
  assign FullAdder_854_io_ci = FullAdder_818_io_co; // @[wallace.scala 71:19]
  assign FullAdder_855_io_a = HalfAdder_78_io_co; // @[wallace.scala 69:18]
  assign FullAdder_855_io_b = FullAdder_818_io_s; // @[wallace.scala 70:18]
  assign FullAdder_855_io_ci = FullAdder_819_io_co; // @[wallace.scala 71:19]
  assign FullAdder_856_io_a = HalfAdder_80_io_co; // @[wallace.scala 69:18]
  assign FullAdder_856_io_b = FullAdder_819_io_s; // @[wallace.scala 70:18]
  assign FullAdder_856_io_ci = HalfAdder_104_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_123_io_a = HalfAdder_104_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_123_io_b = HalfAdder_105_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_124_io_a = FullAdder_820_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_124_io_b = FullAdder_821_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_125_io_a = HalfAdder_81_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_125_io_b = FullAdder_823_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_126_io_a = FullAdder_824_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_126_io_b = FullAdder_825_io_co; // @[wallace.scala 60:18]
  assign FullAdder_857_io_a = FullAdder_772_io_co; // @[wallace.scala 69:18]
  assign FullAdder_857_io_b = FullAdder_773_io_co; // @[wallace.scala 70:18]
  assign FullAdder_857_io_ci = FullAdder_825_io_s; // @[wallace.scala 71:19]
  assign FullAdder_858_io_a = FullAdder_826_io_s; // @[wallace.scala 69:18]
  assign FullAdder_858_io_b = FullAdder_827_io_s; // @[wallace.scala 70:18]
  assign FullAdder_858_io_ci = HalfAdder_106_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_127_io_a = FullAdder_775_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_127_io_b = HalfAdder_106_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_128_io_a = HalfAdder_107_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_128_io_b = FullAdder_828_io_co; // @[wallace.scala 60:18]
  assign FullAdder_859_io_a = FullAdder_776_io_co; // @[wallace.scala 69:18]
  assign FullAdder_859_io_b = HalfAdder_85_io_co; // @[wallace.scala 70:18]
  assign FullAdder_859_io_ci = FullAdder_828_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_129_io_a = HalfAdder_108_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_129_io_b = HalfAdder_109_io_s; // @[wallace.scala 60:18]
  assign FullAdder_860_io_a = FullAdder_779_io_co; // @[wallace.scala 69:18]
  assign FullAdder_860_io_b = FullAdder_780_io_co; // @[wallace.scala 70:18]
  assign FullAdder_860_io_ci = FullAdder_829_io_s; // @[wallace.scala 71:19]
  assign FullAdder_861_io_a = FullAdder_782_io_co; // @[wallace.scala 69:18]
  assign FullAdder_861_io_b = FullAdder_830_io_s; // @[wallace.scala 70:18]
  assign FullAdder_861_io_ci = FullAdder_831_io_co; // @[wallace.scala 71:19]
  assign FullAdder_862_io_a = FullAdder_831_io_s; // @[wallace.scala 69:18]
  assign FullAdder_862_io_b = HalfAdder_110_io_s; // @[wallace.scala 70:18]
  assign FullAdder_862_io_ci = FullAdder_832_io_co; // @[wallace.scala 71:19]
  assign FullAdder_863_io_a = FullAdder_786_io_co; // @[wallace.scala 69:18]
  assign FullAdder_863_io_b = FullAdder_832_io_s; // @[wallace.scala 70:18]
  assign FullAdder_863_io_ci = FullAdder_833_io_co; // @[wallace.scala 71:19]
  assign FullAdder_864_io_a = FullAdder_833_io_s; // @[wallace.scala 69:18]
  assign FullAdder_864_io_b = HalfAdder_111_io_s; // @[wallace.scala 70:18]
  assign FullAdder_864_io_ci = FullAdder_834_io_co; // @[wallace.scala 71:19]
  assign FullAdder_865_io_a = FullAdder_789_io_co; // @[wallace.scala 69:18]
  assign FullAdder_865_io_b = FullAdder_790_io_co; // @[wallace.scala 70:18]
  assign FullAdder_865_io_ci = FullAdder_834_io_s; // @[wallace.scala 71:19]
  assign FullAdder_866_io_a = FullAdder_791_io_co; // @[wallace.scala 69:18]
  assign FullAdder_866_io_b = FullAdder_792_io_co; // @[wallace.scala 70:18]
  assign FullAdder_866_io_ci = FullAdder_835_io_s; // @[wallace.scala 71:19]
  assign FullAdder_867_io_a = FullAdder_794_io_co; // @[wallace.scala 69:18]
  assign FullAdder_867_io_b = FullAdder_836_io_s; // @[wallace.scala 70:18]
  assign FullAdder_867_io_ci = FullAdder_837_io_co; // @[wallace.scala 71:19]
  assign FullAdder_868_io_a = FullAdder_796_io_co; // @[wallace.scala 69:18]
  assign FullAdder_868_io_b = FullAdder_837_io_s; // @[wallace.scala 70:18]
  assign FullAdder_868_io_ci = FullAdder_838_io_co; // @[wallace.scala 71:19]
  assign FullAdder_869_io_a = FullAdder_797_io_co; // @[wallace.scala 69:18]
  assign FullAdder_869_io_b = FullAdder_798_io_co; // @[wallace.scala 70:18]
  assign FullAdder_869_io_ci = FullAdder_838_io_s; // @[wallace.scala 71:19]
  assign FullAdder_870_io_a = FullAdder_800_io_co; // @[wallace.scala 69:18]
  assign FullAdder_870_io_b = FullAdder_839_io_s; // @[wallace.scala 70:18]
  assign FullAdder_870_io_ci = FullAdder_840_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_130_io_a = FullAdder_802_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_130_io_b = FullAdder_840_io_s; // @[wallace.scala 60:18]
  assign FullAdder_871_io_a = HalfAdder_86_io_co; // @[wallace.scala 69:18]
  assign FullAdder_871_io_b = FullAdder_841_io_s; // @[wallace.scala 70:18]
  assign FullAdder_871_io_ci = FullAdder_842_io_co; // @[wallace.scala 71:19]
  assign FullAdder_872_io_a = HalfAdder_88_io_co; // @[wallace.scala 69:18]
  assign FullAdder_872_io_b = FullAdder_842_io_s; // @[wallace.scala 70:18]
  assign FullAdder_872_io_ci = HalfAdder_112_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_131_io_a = HalfAdder_89_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_131_io_b = HalfAdder_112_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_132_io_a = HalfAdder_113_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_132_io_b = FullAdder_843_io_co; // @[wallace.scala 60:18]
  assign FullAdder_873_io_a = FullAdder_806_io_co; // @[wallace.scala 69:18]
  assign FullAdder_873_io_b = FullAdder_843_io_s; // @[wallace.scala 70:18]
  assign FullAdder_873_io_ci = FullAdder_844_io_co; // @[wallace.scala 71:19]
  assign FullAdder_874_io_a = FullAdder_810_io_co; // @[wallace.scala 69:18]
  assign FullAdder_874_io_b = FullAdder_847_io_s; // @[wallace.scala 70:18]
  assign FullAdder_874_io_ci = FullAdder_848_io_co; // @[wallace.scala 71:19]
  assign FullAdder_875_io_a = HalfAdder_91_io_co; // @[wallace.scala 69:18]
  assign FullAdder_875_io_b = FullAdder_849_io_s; // @[wallace.scala 70:18]
  assign FullAdder_875_io_ci = HalfAdder_114_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_133_io_a = FullAdder_812_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_133_io_b = HalfAdder_114_io_s; // @[wallace.scala 60:18]
  assign FullAdder_876_io_a = FullAdder_813_io_s; // @[wallace.scala 69:18]
  assign FullAdder_876_io_b = FullAdder_814_io_co; // @[wallace.scala 70:18]
  assign FullAdder_876_io_ci = FullAdder_850_io_co; // @[wallace.scala 71:19]
  assign FullAdder_877_io_a = HalfAdder_92_io_co; // @[wallace.scala 69:18]
  assign FullAdder_877_io_b = FullAdder_850_io_s; // @[wallace.scala 70:18]
  assign FullAdder_877_io_ci = HalfAdder_115_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_134_io_a = FullAdder_815_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_134_io_b = HalfAdder_115_io_s; // @[wallace.scala 60:18]
  assign FullAdder_878_io_a = FullAdder_815_io_s; // @[wallace.scala 69:18]
  assign FullAdder_878_io_b = FullAdder_816_io_co; // @[wallace.scala 70:18]
  assign FullAdder_878_io_ci = HalfAdder_116_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_135_io_a = HalfAdder_116_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_135_io_b = HalfAdder_117_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_136_io_a = HalfAdder_94_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_136_io_b = HalfAdder_117_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_137_io_a = HalfAdder_94_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_137_io_b = FullAdder_851_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_138_io_a = HalfAdder_96_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_138_io_b = HalfAdder_118_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_139_io_a = HalfAdder_97_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_139_io_b = FullAdder_852_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_140_io_a = HalfAdder_99_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_140_io_b = FullAdder_853_io_co; // @[wallace.scala 60:18]
  assign FullAdder_879_io_a = FullAdder_817_io_s; // @[wallace.scala 69:18]
  assign FullAdder_879_io_b = HalfAdder_102_io_co; // @[wallace.scala 70:18]
  assign FullAdder_879_io_ci = HalfAdder_122_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_141_io_a = HalfAdder_103_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_141_io_b = FullAdder_854_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_142_io_a = FullAdder_855_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_142_io_b = FullAdder_856_io_co; // @[wallace.scala 60:18]
  assign FullAdder_880_io_a = HalfAdder_105_io_co; // @[wallace.scala 69:18]
  assign FullAdder_880_io_b = FullAdder_856_io_s; // @[wallace.scala 70:18]
  assign FullAdder_880_io_ci = HalfAdder_123_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_143_io_a = FullAdder_820_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_143_io_b = HalfAdder_123_io_s; // @[wallace.scala 60:18]
  assign FullAdder_881_io_a = FullAdder_822_io_s; // @[wallace.scala 69:18]
  assign FullAdder_881_io_b = FullAdder_823_io_co; // @[wallace.scala 70:18]
  assign FullAdder_881_io_ci = HalfAdder_125_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_144_io_a = FullAdder_824_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_144_io_b = HalfAdder_125_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_145_io_a = HalfAdder_126_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_145_io_b = FullAdder_857_io_co; // @[wallace.scala 60:18]
  assign FullAdder_882_io_a = FullAdder_826_io_co; // @[wallace.scala 69:18]
  assign FullAdder_882_io_b = FullAdder_827_io_co; // @[wallace.scala 70:18]
  assign FullAdder_882_io_ci = FullAdder_857_io_s; // @[wallace.scala 71:19]
  assign FullAdder_883_io_a = HalfAdder_107_io_co; // @[wallace.scala 69:18]
  assign FullAdder_883_io_b = FullAdder_858_io_s; // @[wallace.scala 70:18]
  assign FullAdder_883_io_ci = HalfAdder_127_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_146_io_a = HalfAdder_127_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_146_io_b = HalfAdder_128_io_s; // @[wallace.scala 60:18]
  assign FullAdder_884_io_a = HalfAdder_108_io_co; // @[wallace.scala 69:18]
  assign FullAdder_884_io_b = HalfAdder_109_io_co; // @[wallace.scala 70:18]
  assign FullAdder_884_io_ci = FullAdder_859_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_147_io_a = FullAdder_829_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_147_io_b = HalfAdder_129_io_s; // @[wallace.scala 60:18]
  assign FullAdder_885_io_a = FullAdder_830_io_co; // @[wallace.scala 69:18]
  assign FullAdder_885_io_b = FullAdder_860_io_s; // @[wallace.scala 70:18]
  assign FullAdder_885_io_ci = FullAdder_861_io_co; // @[wallace.scala 71:19]
  assign FullAdder_886_io_a = HalfAdder_110_io_co; // @[wallace.scala 69:18]
  assign FullAdder_886_io_b = FullAdder_861_io_s; // @[wallace.scala 70:18]
  assign FullAdder_886_io_ci = FullAdder_862_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_148_io_a = FullAdder_862_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_148_io_b = FullAdder_863_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_149_io_a = HalfAdder_111_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_149_io_b = FullAdder_863_io_s; // @[wallace.scala 60:18]
  assign FullAdder_887_io_a = FullAdder_835_io_co; // @[wallace.scala 69:18]
  assign FullAdder_887_io_b = FullAdder_865_io_s; // @[wallace.scala 70:18]
  assign FullAdder_887_io_ci = FullAdder_866_io_co; // @[wallace.scala 71:19]
  assign FullAdder_888_io_a = FullAdder_836_io_co; // @[wallace.scala 69:18]
  assign FullAdder_888_io_b = FullAdder_866_io_s; // @[wallace.scala 70:18]
  assign FullAdder_888_io_ci = FullAdder_867_io_co; // @[wallace.scala 71:19]
  assign FullAdder_889_io_a = FullAdder_839_io_co; // @[wallace.scala 69:18]
  assign FullAdder_889_io_b = FullAdder_869_io_s; // @[wallace.scala 70:18]
  assign FullAdder_889_io_ci = FullAdder_870_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_150_io_a = FullAdder_870_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_150_io_b = HalfAdder_130_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_151_io_a = FullAdder_841_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_151_io_b = HalfAdder_130_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_152_io_a = FullAdder_871_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_152_io_b = FullAdder_872_io_co; // @[wallace.scala 60:18]
  assign FullAdder_890_io_a = HalfAdder_113_io_co; // @[wallace.scala 69:18]
  assign FullAdder_890_io_b = FullAdder_872_io_s; // @[wallace.scala 70:18]
  assign FullAdder_890_io_ci = HalfAdder_131_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_153_io_a = HalfAdder_131_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_153_io_b = HalfAdder_132_io_s; // @[wallace.scala 60:18]
  assign FullAdder_891_io_a = FullAdder_846_io_s; // @[wallace.scala 69:18]
  assign FullAdder_891_io_b = FullAdder_847_io_co; // @[wallace.scala 70:18]
  assign FullAdder_891_io_ci = FullAdder_874_io_co; // @[wallace.scala 71:19]
  assign FullAdder_892_io_a = FullAdder_848_io_s; // @[wallace.scala 69:18]
  assign FullAdder_892_io_b = FullAdder_849_io_co; // @[wallace.scala 70:18]
  assign FullAdder_892_io_ci = FullAdder_875_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_154_io_a = FullAdder_875_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_154_io_b = HalfAdder_133_io_co; // @[wallace.scala 60:18]
  assign FullAdder_893_io_a = FullAdder_812_io_s; // @[wallace.scala 69:18]
  assign FullAdder_893_io_b = FullAdder_813_io_co; // @[wallace.scala 70:18]
  assign FullAdder_893_io_ci = FullAdder_876_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_155_io_a = HalfAdder_134_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_155_io_b = FullAdder_878_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_156_io_a = HalfAdder_135_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_156_io_b = HalfAdder_136_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_157_io_a = HalfAdder_136_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_157_io_b = HalfAdder_137_io_co; // @[wallace.scala 60:18]
  assign FullAdder_894_io_a = FullAdder_851_io_s; // @[wallace.scala 69:18]
  assign FullAdder_894_io_b = HalfAdder_118_io_co; // @[wallace.scala 70:18]
  assign FullAdder_894_io_ci = HalfAdder_138_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_158_io_a = HalfAdder_119_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_158_io_b = HalfAdder_140_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_159_io_a = HalfAdder_121_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_159_io_b = FullAdder_879_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_160_io_a = HalfAdder_122_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_160_io_b = HalfAdder_141_io_co; // @[wallace.scala 60:18]
  assign FullAdder_895_io_a = FullAdder_854_io_s; // @[wallace.scala 69:18]
  assign FullAdder_895_io_b = FullAdder_855_io_co; // @[wallace.scala 70:18]
  assign FullAdder_895_io_ci = HalfAdder_142_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_161_io_a = FullAdder_880_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_161_io_b = HalfAdder_143_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_162_io_a = HalfAdder_124_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_162_io_b = HalfAdder_143_io_s; // @[wallace.scala 60:18]
  assign FullAdder_896_io_a = FullAdder_821_io_s; // @[wallace.scala 69:18]
  assign FullAdder_896_io_b = FullAdder_822_io_co; // @[wallace.scala 70:18]
  assign FullAdder_896_io_ci = FullAdder_881_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_163_io_a = HalfAdder_126_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_163_io_b = HalfAdder_144_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_164_io_a = HalfAdder_145_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_164_io_b = FullAdder_882_io_co; // @[wallace.scala 60:18]
  assign FullAdder_897_io_a = FullAdder_858_io_co; // @[wallace.scala 69:18]
  assign FullAdder_897_io_b = FullAdder_882_io_s; // @[wallace.scala 70:18]
  assign FullAdder_897_io_ci = FullAdder_883_io_co; // @[wallace.scala 71:19]
  assign FullAdder_898_io_a = HalfAdder_128_io_co; // @[wallace.scala 69:18]
  assign FullAdder_898_io_b = FullAdder_883_io_s; // @[wallace.scala 70:18]
  assign FullAdder_898_io_ci = HalfAdder_146_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_165_io_a = FullAdder_859_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_165_io_b = HalfAdder_146_io_s; // @[wallace.scala 60:18]
  assign FullAdder_899_io_a = HalfAdder_129_io_co; // @[wallace.scala 69:18]
  assign FullAdder_899_io_b = FullAdder_884_io_s; // @[wallace.scala 70:18]
  assign FullAdder_899_io_ci = HalfAdder_147_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_166_io_a = FullAdder_860_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_166_io_b = HalfAdder_147_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_167_io_a = FullAdder_864_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_167_io_b = HalfAdder_149_io_s; // @[wallace.scala 60:18]
  assign FullAdder_900_io_a = FullAdder_864_io_s; // @[wallace.scala 69:18]
  assign FullAdder_900_io_b = FullAdder_865_io_co; // @[wallace.scala 70:18]
  assign FullAdder_900_io_ci = FullAdder_887_io_co; // @[wallace.scala 71:19]
  assign FullAdder_901_io_a = FullAdder_868_io_s; // @[wallace.scala 69:18]
  assign FullAdder_901_io_b = FullAdder_869_io_co; // @[wallace.scala 70:18]
  assign FullAdder_901_io_ci = FullAdder_889_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_168_io_a = FullAdder_871_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_168_io_b = HalfAdder_151_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_169_io_a = HalfAdder_152_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_169_io_b = FullAdder_890_io_co; // @[wallace.scala 60:18]
  assign FullAdder_902_io_a = HalfAdder_132_io_co; // @[wallace.scala 69:18]
  assign FullAdder_902_io_b = FullAdder_890_io_s; // @[wallace.scala 70:18]
  assign FullAdder_902_io_ci = HalfAdder_153_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_170_io_a = FullAdder_873_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_170_io_b = HalfAdder_153_io_s; // @[wallace.scala 60:18]
  assign FullAdder_903_io_a = FullAdder_845_io_s; // @[wallace.scala 69:18]
  assign FullAdder_903_io_b = FullAdder_846_io_co; // @[wallace.scala 70:18]
  assign FullAdder_903_io_ci = FullAdder_891_io_co; // @[wallace.scala 71:19]
  assign FullAdder_904_io_a = FullAdder_877_io_s; // @[wallace.scala 69:18]
  assign FullAdder_904_io_b = HalfAdder_134_io_co; // @[wallace.scala 70:18]
  assign FullAdder_904_io_ci = HalfAdder_155_io_co; // @[wallace.scala 71:19]
  assign FullAdder_905_io_a = FullAdder_878_io_s; // @[wallace.scala 69:18]
  assign FullAdder_905_io_b = HalfAdder_135_io_co; // @[wallace.scala 70:18]
  assign FullAdder_905_io_ci = HalfAdder_156_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_171_io_a = HalfAdder_137_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_171_io_b = FullAdder_894_io_co; // @[wallace.scala 60:18]
  assign FullAdder_906_io_a = FullAdder_852_io_s; // @[wallace.scala 69:18]
  assign FullAdder_906_io_b = HalfAdder_119_io_co; // @[wallace.scala 70:18]
  assign FullAdder_906_io_ci = HalfAdder_158_io_co; // @[wallace.scala 71:19]
  assign FullAdder_907_io_a = HalfAdder_120_io_s; // @[wallace.scala 69:18]
  assign FullAdder_907_io_b = HalfAdder_121_io_co; // @[wallace.scala 70:18]
  assign FullAdder_907_io_ci = HalfAdder_159_io_co; // @[wallace.scala 71:19]
  assign FullAdder_908_io_a = HalfAdder_142_io_s; // @[wallace.scala 69:18]
  assign FullAdder_908_io_b = FullAdder_880_io_co; // @[wallace.scala 70:18]
  assign FullAdder_908_io_ci = HalfAdder_161_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_172_io_a = HalfAdder_161_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_172_io_b = HalfAdder_162_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_173_io_a = HalfAdder_124_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_173_io_b = FullAdder_896_io_co; // @[wallace.scala 60:18]
  assign FullAdder_909_io_a = FullAdder_881_io_s; // @[wallace.scala 69:18]
  assign FullAdder_909_io_b = HalfAdder_144_io_co; // @[wallace.scala 70:18]
  assign FullAdder_909_io_ci = HalfAdder_163_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_174_io_a = HalfAdder_145_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_174_io_b = HalfAdder_163_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_175_io_a = FullAdder_884_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_175_io_b = HalfAdder_165_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_176_io_a = FullAdder_885_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_176_io_b = HalfAdder_166_io_s; // @[wallace.scala 60:18]
  assign FullAdder_910_io_a = HalfAdder_148_io_s; // @[wallace.scala 69:18]
  assign FullAdder_910_io_b = HalfAdder_149_io_co; // @[wallace.scala 70:18]
  assign FullAdder_910_io_ci = HalfAdder_167_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_177_io_a = HalfAdder_167_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_177_io_b = FullAdder_900_io_co; // @[wallace.scala 60:18]
  assign FullAdder_911_io_a = FullAdder_867_io_s; // @[wallace.scala 69:18]
  assign FullAdder_911_io_b = FullAdder_868_io_co; // @[wallace.scala 70:18]
  assign FullAdder_911_io_ci = FullAdder_901_io_co; // @[wallace.scala 71:19]
  assign FullAdder_912_io_a = HalfAdder_150_io_s; // @[wallace.scala 69:18]
  assign FullAdder_912_io_b = HalfAdder_151_io_co; // @[wallace.scala 70:18]
  assign FullAdder_912_io_ci = HalfAdder_168_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_178_io_a = HalfAdder_152_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_178_io_b = HalfAdder_168_io_s; // @[wallace.scala 60:18]
  assign FullAdder_913_io_a = FullAdder_844_io_s; // @[wallace.scala 69:18]
  assign FullAdder_913_io_b = FullAdder_845_io_co; // @[wallace.scala 70:18]
  assign FullAdder_913_io_ci = FullAdder_903_io_co; // @[wallace.scala 71:19]
  assign FullAdder_914_io_a = FullAdder_876_io_s; // @[wallace.scala 69:18]
  assign FullAdder_914_io_b = FullAdder_877_io_co; // @[wallace.scala 70:18]
  assign FullAdder_914_io_ci = FullAdder_904_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_179_io_a = HalfAdder_155_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_179_io_b = FullAdder_905_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_180_io_a = HalfAdder_157_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_180_io_b = HalfAdder_171_io_co; // @[wallace.scala 60:18]
  assign FullAdder_915_io_a = FullAdder_853_io_s; // @[wallace.scala 69:18]
  assign FullAdder_915_io_b = HalfAdder_120_io_co; // @[wallace.scala 70:18]
  assign FullAdder_915_io_ci = FullAdder_907_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_181_io_a = HalfAdder_162_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_181_io_b = HalfAdder_173_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_182_io_a = HalfAdder_164_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_182_io_b = HalfAdder_174_io_s; // @[wallace.scala 60:18]
  assign FullAdder_916_io_a = FullAdder_898_io_s; // @[wallace.scala 69:18]
  assign FullAdder_916_io_b = HalfAdder_165_io_co; // @[wallace.scala 70:18]
  assign FullAdder_916_io_ci = HalfAdder_175_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_183_io_a = FullAdder_899_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_183_io_b = HalfAdder_175_io_s; // @[wallace.scala 60:18]
  assign FullAdder_917_io_a = FullAdder_899_io_s; // @[wallace.scala 69:18]
  assign FullAdder_917_io_b = HalfAdder_166_io_co; // @[wallace.scala 70:18]
  assign FullAdder_917_io_ci = HalfAdder_176_io_co; // @[wallace.scala 71:19]
  assign FullAdder_918_io_a = FullAdder_886_io_s; // @[wallace.scala 69:18]
  assign FullAdder_918_io_b = HalfAdder_148_io_co; // @[wallace.scala 70:18]
  assign FullAdder_918_io_ci = FullAdder_910_io_co; // @[wallace.scala 71:19]
  assign FullAdder_919_io_a = FullAdder_889_io_s; // @[wallace.scala 69:18]
  assign FullAdder_919_io_b = HalfAdder_150_io_co; // @[wallace.scala 70:18]
  assign FullAdder_919_io_ci = FullAdder_912_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_184_io_a = HalfAdder_169_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_184_io_b = HalfAdder_178_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_185_io_a = FullAdder_873_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_185_io_b = FullAdder_913_io_co; // @[wallace.scala 60:18]
  assign FullAdder_920_io_a = HalfAdder_156_io_s; // @[wallace.scala 69:18]
  assign FullAdder_920_io_b = HalfAdder_157_io_co; // @[wallace.scala 70:18]
  assign FullAdder_920_io_ci = HalfAdder_180_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_186_io_a = HalfAdder_172_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_186_io_b = HalfAdder_181_io_co; // @[wallace.scala 60:18]
  assign FullAdder_921_io_a = FullAdder_909_io_s; // @[wallace.scala 69:18]
  assign FullAdder_921_io_b = HalfAdder_174_io_co; // @[wallace.scala 70:18]
  assign FullAdder_921_io_ci = HalfAdder_182_io_co; // @[wallace.scala 71:19]
  assign FullAdder_922_io_a = FullAdder_897_io_s; // @[wallace.scala 69:18]
  assign FullAdder_922_io_b = FullAdder_898_io_co; // @[wallace.scala 70:18]
  assign FullAdder_922_io_ci = FullAdder_916_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_187_io_a = HalfAdder_183_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_187_io_b = FullAdder_917_io_co; // @[wallace.scala 60:18]
  assign FullAdder_923_io_a = FullAdder_885_io_s; // @[wallace.scala 69:18]
  assign FullAdder_923_io_b = FullAdder_886_io_co; // @[wallace.scala 70:18]
  assign FullAdder_923_io_ci = FullAdder_918_io_co; // @[wallace.scala 71:19]
  assign FullAdder_924_io_a = FullAdder_912_io_s; // @[wallace.scala 69:18]
  assign FullAdder_924_io_b = HalfAdder_178_io_co; // @[wallace.scala 70:18]
  assign FullAdder_924_io_ci = HalfAdder_184_io_co; // @[wallace.scala 71:19]
  assign FullAdder_925_io_a = FullAdder_908_io_s; // @[wallace.scala 69:18]
  assign FullAdder_925_io_b = HalfAdder_172_io_co; // @[wallace.scala 70:18]
  assign FullAdder_925_io_ci = HalfAdder_186_io_co; // @[wallace.scala 71:19]
  assign FullAdder_926_io_a = FullAdder_896_io_s; // @[wallace.scala 69:18]
  assign FullAdder_926_io_b = FullAdder_909_io_co; // @[wallace.scala 70:18]
  assign FullAdder_926_io_ci = FullAdder_921_io_co; // @[wallace.scala 71:19]
  assign FullAdder_927_io_a = HalfAdder_164_io_s; // @[wallace.scala 69:18]
  assign FullAdder_927_io_b = FullAdder_897_io_co; // @[wallace.scala 70:18]
  assign FullAdder_927_io_ci = FullAdder_922_io_co; // @[wallace.scala 71:19]
  assign FullAdder_928_io_a = FullAdder_916_io_s; // @[wallace.scala 69:18]
  assign FullAdder_928_io_b = HalfAdder_183_io_co; // @[wallace.scala 70:18]
  assign FullAdder_928_io_ci = HalfAdder_187_io_co; // @[wallace.scala 71:19]
  assign FullAdder_929_io_a = FullAdder_895_io_s; // @[wallace.scala 69:18]
  assign FullAdder_929_io_b = FullAdder_908_io_co; // @[wallace.scala 70:18]
  assign FullAdder_929_io_ci = FullAdder_925_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_188_io_a = HalfAdder_173_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_188_io_b = FullAdder_926_io_co; // @[wallace.scala 60:18]
  assign FullAdder_930_io_a = HalfAdder_141_io_s; // @[wallace.scala 69:18]
  assign FullAdder_930_io_b = FullAdder_895_io_co; // @[wallace.scala 70:18]
  assign FullAdder_930_io_ci = FullAdder_929_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_189_io_a = HalfAdder_181_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_189_io_b = HalfAdder_188_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_190_io_a = HalfAdder_186_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_190_io_b = HalfAdder_189_io_co; // @[wallace.scala 60:18]
endmodule
module MUL(
  input  [31:0] io_multiplicand,
  input  [31:0] io_multiplier,
  output [62:0] io_outs
);
  wire [31:0] pp_io_multiplicand; // @[mul.scala 26:18]
  wire [31:0] pp_io_multiplier; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_0; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_1; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_2; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_3; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_4; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_5; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_6; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_7; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_8; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_9; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_10; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_11; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_12; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_13; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_14; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_15; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_16; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_17; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_18; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_19; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_20; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_21; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_22; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_23; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_24; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_25; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_26; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_27; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_28; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_29; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_30; // @[mul.scala 26:18]
  wire [31:0] pp_io_outs_31; // @[mul.scala 26:18]
  wire [31:0] wt_io_pp_0; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_1; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_2; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_3; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_4; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_5; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_6; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_7; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_8; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_9; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_10; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_11; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_12; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_13; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_14; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_15; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_16; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_17; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_18; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_19; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_20; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_21; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_22; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_23; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_24; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_25; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_26; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_27; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_28; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_29; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_30; // @[mul.scala 30:18]
  wire [31:0] wt_io_pp_31; // @[mul.scala 30:18]
  wire [63:0] wt_io_augend; // @[mul.scala 30:18]
  wire [63:0] wt_io_addend; // @[mul.scala 30:18]
  wire [63:0] _T_1 = wt_io_augend + wt_io_addend; // @[mul.scala 37:27]
  PartialProd pp ( // @[mul.scala 26:18]
    .io_multiplicand(pp_io_multiplicand),
    .io_multiplier(pp_io_multiplier),
    .io_outs_0(pp_io_outs_0),
    .io_outs_1(pp_io_outs_1),
    .io_outs_2(pp_io_outs_2),
    .io_outs_3(pp_io_outs_3),
    .io_outs_4(pp_io_outs_4),
    .io_outs_5(pp_io_outs_5),
    .io_outs_6(pp_io_outs_6),
    .io_outs_7(pp_io_outs_7),
    .io_outs_8(pp_io_outs_8),
    .io_outs_9(pp_io_outs_9),
    .io_outs_10(pp_io_outs_10),
    .io_outs_11(pp_io_outs_11),
    .io_outs_12(pp_io_outs_12),
    .io_outs_13(pp_io_outs_13),
    .io_outs_14(pp_io_outs_14),
    .io_outs_15(pp_io_outs_15),
    .io_outs_16(pp_io_outs_16),
    .io_outs_17(pp_io_outs_17),
    .io_outs_18(pp_io_outs_18),
    .io_outs_19(pp_io_outs_19),
    .io_outs_20(pp_io_outs_20),
    .io_outs_21(pp_io_outs_21),
    .io_outs_22(pp_io_outs_22),
    .io_outs_23(pp_io_outs_23),
    .io_outs_24(pp_io_outs_24),
    .io_outs_25(pp_io_outs_25),
    .io_outs_26(pp_io_outs_26),
    .io_outs_27(pp_io_outs_27),
    .io_outs_28(pp_io_outs_28),
    .io_outs_29(pp_io_outs_29),
    .io_outs_30(pp_io_outs_30),
    .io_outs_31(pp_io_outs_31)
  );
  Wallace wt ( // @[mul.scala 30:18]
    .io_pp_0(wt_io_pp_0),
    .io_pp_1(wt_io_pp_1),
    .io_pp_2(wt_io_pp_2),
    .io_pp_3(wt_io_pp_3),
    .io_pp_4(wt_io_pp_4),
    .io_pp_5(wt_io_pp_5),
    .io_pp_6(wt_io_pp_6),
    .io_pp_7(wt_io_pp_7),
    .io_pp_8(wt_io_pp_8),
    .io_pp_9(wt_io_pp_9),
    .io_pp_10(wt_io_pp_10),
    .io_pp_11(wt_io_pp_11),
    .io_pp_12(wt_io_pp_12),
    .io_pp_13(wt_io_pp_13),
    .io_pp_14(wt_io_pp_14),
    .io_pp_15(wt_io_pp_15),
    .io_pp_16(wt_io_pp_16),
    .io_pp_17(wt_io_pp_17),
    .io_pp_18(wt_io_pp_18),
    .io_pp_19(wt_io_pp_19),
    .io_pp_20(wt_io_pp_20),
    .io_pp_21(wt_io_pp_21),
    .io_pp_22(wt_io_pp_22),
    .io_pp_23(wt_io_pp_23),
    .io_pp_24(wt_io_pp_24),
    .io_pp_25(wt_io_pp_25),
    .io_pp_26(wt_io_pp_26),
    .io_pp_27(wt_io_pp_27),
    .io_pp_28(wt_io_pp_28),
    .io_pp_29(wt_io_pp_29),
    .io_pp_30(wt_io_pp_30),
    .io_pp_31(wt_io_pp_31),
    .io_augend(wt_io_augend),
    .io_addend(wt_io_addend)
  );
  assign io_outs = _T_1[62:0]; // @[mul.scala 37:11]
  assign pp_io_multiplicand = io_multiplicand; // @[mul.scala 27:22]
  assign pp_io_multiplier = io_multiplier; // @[mul.scala 28:20]
  assign wt_io_pp_0 = pp_io_outs_0; // @[mul.scala 31:12]
  assign wt_io_pp_1 = pp_io_outs_1; // @[mul.scala 31:12]
  assign wt_io_pp_2 = pp_io_outs_2; // @[mul.scala 31:12]
  assign wt_io_pp_3 = pp_io_outs_3; // @[mul.scala 31:12]
  assign wt_io_pp_4 = pp_io_outs_4; // @[mul.scala 31:12]
  assign wt_io_pp_5 = pp_io_outs_5; // @[mul.scala 31:12]
  assign wt_io_pp_6 = pp_io_outs_6; // @[mul.scala 31:12]
  assign wt_io_pp_7 = pp_io_outs_7; // @[mul.scala 31:12]
  assign wt_io_pp_8 = pp_io_outs_8; // @[mul.scala 31:12]
  assign wt_io_pp_9 = pp_io_outs_9; // @[mul.scala 31:12]
  assign wt_io_pp_10 = pp_io_outs_10; // @[mul.scala 31:12]
  assign wt_io_pp_11 = pp_io_outs_11; // @[mul.scala 31:12]
  assign wt_io_pp_12 = pp_io_outs_12; // @[mul.scala 31:12]
  assign wt_io_pp_13 = pp_io_outs_13; // @[mul.scala 31:12]
  assign wt_io_pp_14 = pp_io_outs_14; // @[mul.scala 31:12]
  assign wt_io_pp_15 = pp_io_outs_15; // @[mul.scala 31:12]
  assign wt_io_pp_16 = pp_io_outs_16; // @[mul.scala 31:12]
  assign wt_io_pp_17 = pp_io_outs_17; // @[mul.scala 31:12]
  assign wt_io_pp_18 = pp_io_outs_18; // @[mul.scala 31:12]
  assign wt_io_pp_19 = pp_io_outs_19; // @[mul.scala 31:12]
  assign wt_io_pp_20 = pp_io_outs_20; // @[mul.scala 31:12]
  assign wt_io_pp_21 = pp_io_outs_21; // @[mul.scala 31:12]
  assign wt_io_pp_22 = pp_io_outs_22; // @[mul.scala 31:12]
  assign wt_io_pp_23 = pp_io_outs_23; // @[mul.scala 31:12]
  assign wt_io_pp_24 = pp_io_outs_24; // @[mul.scala 31:12]
  assign wt_io_pp_25 = pp_io_outs_25; // @[mul.scala 31:12]
  assign wt_io_pp_26 = pp_io_outs_26; // @[mul.scala 31:12]
  assign wt_io_pp_27 = pp_io_outs_27; // @[mul.scala 31:12]
  assign wt_io_pp_28 = pp_io_outs_28; // @[mul.scala 31:12]
  assign wt_io_pp_29 = pp_io_outs_29; // @[mul.scala 31:12]
  assign wt_io_pp_30 = pp_io_outs_30; // @[mul.scala 31:12]
  assign wt_io_pp_31 = pp_io_outs_31; // @[mul.scala 31:12]
endmodule
