module ks64 (in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, in100, in101, in102, in103, in104, in105, in106, in107, in108, in109, in110, in111, in112, in113, in114, in115, in116, in117, in118, in119, in120, in121, in122, in123, in124, in125, in126, in127, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, out30, out31, out32, out33, out34, out35, out36, out37, out38, out39, out40, out41, out42, out43, out44, out45, out46, out47, out48, out49, out50, out51, out52, out53, out54, out55, out56, out57, out58, out59, out60, out61, out62, out63, out64, );
input in0;
input in1;
input in2;
input in3;
input in4;
input in5;
input in6;
input in7;
input in8;
input in9;
input in10;
input in11;
input in12;
input in13;
input in14;
input in15;
input in16;
input in17;
input in18;
input in19;
input in20;
input in21;
input in22;
input in23;
input in24;
input in25;
input in26;
input in27;
input in28;
input in29;
input in30;
input in31;
input in32;
input in33;
input in34;
input in35;
input in36;
input in37;
input in38;
input in39;
input in40;
input in41;
input in42;
input in43;
input in44;
input in45;
input in46;
input in47;
input in48;
input in49;
input in50;
input in51;
input in52;
input in53;
input in54;
input in55;
input in56;
input in57;
input in58;
input in59;
input in60;
input in61;
input in62;
input in63;
input in64;
input in65;
input in66;
input in67;
input in68;
input in69;
input in70;
input in71;
input in72;
input in73;
input in74;
input in75;
input in76;
input in77;
input in78;
input in79;
input in80;
input in81;
input in82;
input in83;
input in84;
input in85;
input in86;
input in87;
input in88;
input in89;
input in90;
input in91;
input in92;
input in93;
input in94;
input in95;
input in96;
input in97;
input in98;
input in99;
input in100;
input in101;
input in102;
input in103;
input in104;
input in105;
input in106;
input in107;
input in108;
input in109;
input in110;
input in111;
input in112;
input in113;
input in114;
input in115;
input in116;
input in117;
input in118;
input in119;
input in120;
input in121;
input in122;
input in123;
input in124;
input in125;
input in126;
input in127;
output out0;
output out1;
output out2;
output out3;
output out4;
output out5;
output out6;
output out7;
output out8;
output out9;
output out10;
output out11;
output out12;
output out13;
output out14;
output out15;
output out16;
output out17;
output out18;
output out19;
output out20;
output out21;
output out22;
output out23;
output out24;
output out25;
output out26;
output out27;
output out28;
output out29;
output out30;
output out31;
output out32;
output out33;
output out34;
output out35;
output out36;
output out37;
output out38;
output out39;
output out40;
output out41;
output out42;
output out43;
output out44;
output out45;
output out46;
output out47;
output out48;
output out49;
output out50;
output out51;
output out52;
output out53;
output out54;
output out55;
output out56;
output out57;
output out58;
output out59;
output out60;
output out61;
output out62;
output out63;
output out64;
wire var0;
wire var1;
wire var2;
wire var3;
wire var4;
wire var5;
wire var6;
wire var7;
wire var8;
wire var9;
wire var10;
wire var11;
wire var12;
wire var13;
wire var14;
wire var15;
wire var16;
wire var17;
wire var18;
wire var19;
wire var20;
wire var21;
wire var22;
wire var23;
wire var24;
wire var25;
wire var26;
wire var27;
wire var28;
wire var29;
wire var30;
wire var31;
wire var32;
wire var33;
wire var34;
wire var35;
wire var36;
wire var37;
wire var38;
wire var39;
wire var40;
wire var41;
wire var42;
wire var43;
wire var44;
wire var45;
wire var46;
wire var47;
wire var48;
wire var49;
wire var50;
wire var51;
wire var52;
wire var53;
wire var54;
wire var55;
wire var56;
wire var57;
wire var58;
wire var59;
wire var60;
wire var61;
wire var62;
wire var63;
wire var64;
wire var65;
wire var66;
wire var67;
wire var68;
wire var69;
wire var70;
wire var71;
wire var72;
wire var73;
wire var74;
wire var75;
wire var76;
wire var77;
wire var78;
wire var79;
wire var80;
wire var81;
wire var82;
wire var83;
wire var84;
wire var85;
wire var86;
wire var87;
wire var88;
wire var89;
wire var90;
wire var91;
wire var92;
wire var93;
wire var94;
wire var95;
wire var96;
wire var97;
wire var98;
wire var99;
wire var100;
wire var101;
wire var102;
wire var103;
wire var104;
wire var105;
wire var106;
wire var107;
wire var108;
wire var109;
wire var110;
wire var111;
wire var112;
wire var113;
wire var114;
wire var115;
wire var116;
wire var117;
wire var118;
wire var119;
wire var120;
wire var121;
wire var122;
wire var123;
wire var124;
wire var125;
wire var126;
wire var127;
wire var128;
wire var129;
wire var130;
wire var131;
wire var132;
wire var133;
wire var134;
wire var135;
wire var136;
wire var137;
wire var138;
wire var139;
wire var140;
wire var141;
wire var142;
wire var143;
wire var144;
wire var145;
wire var146;
wire var147;
wire var148;
wire var149;
wire var150;
wire var151;
wire var152;
wire var153;
wire var154;
wire var155;
wire var156;
wire var157;
wire var158;
wire var159;
wire var160;
wire var161;
wire var162;
wire var163;
wire var164;
wire var165;
wire var166;
wire var167;
wire var168;
wire var169;
wire var170;
wire var171;
wire var172;
wire var173;
wire var174;
wire var175;
wire var176;
wire var177;
wire var178;
wire var179;
wire var180;
wire var181;
wire var182;
wire var183;
wire var184;
wire var185;
wire var186;
wire var187;
wire var188;
wire var189;
wire var190;
wire var191;
wire var192;
wire var193;
wire var194;
wire var195;
wire var196;
wire var197;
wire var198;
wire var199;
wire var200;
wire var201;
wire var202;
wire var203;
wire var204;
wire var205;
wire var206;
wire var207;
wire var208;
wire var209;
wire var210;
wire var211;
wire var212;
wire var213;
wire var214;
wire var215;
wire var216;
wire var217;
wire var218;
wire var219;
wire var220;
wire var221;
wire var222;
wire var223;
wire var224;
wire var225;
wire var226;
wire var227;
wire var228;
wire var229;
wire var230;
wire var231;
wire var232;
wire var233;
wire var234;
wire var235;
wire var236;
wire var237;
wire var238;
wire var239;
wire var240;
wire var241;
wire var242;
wire var243;
wire var244;
wire var245;
wire var246;
wire var247;
wire var248;
wire var249;
wire var250;
wire var251;
wire var252;
wire var253;
wire var254;
wire var255;
wire var256;
wire var257;
wire var258;
wire var259;
wire var260;
wire var261;
wire var262;
wire var263;
wire var264;
wire var265;
wire var266;
wire var267;
wire var268;
wire var269;
wire var270;
wire var271;
wire var272;
wire var273;
wire var274;
wire var275;
wire var276;
wire var277;
wire var278;
wire var279;
wire var280;
wire var281;
wire var282;
wire var283;
wire var284;
wire var285;
wire var286;
wire var287;
wire var288;
wire var289;
wire var290;
wire var291;
wire var292;
wire var293;
wire var294;
wire var295;
wire var296;
wire var297;
wire var298;
wire var299;
wire var300;
wire var301;
wire var302;
wire var303;
wire var304;
wire var305;
wire var306;
wire var307;
wire var308;
wire var309;
wire var310;
wire var311;
wire var312;
wire var313;
wire var314;
wire var315;
wire var316;
wire var317;
wire var318;
wire var319;
wire var320;
wire var321;
wire var322;
wire var323;
wire var324;
wire var325;
wire var326;
wire var327;
wire var328;
wire var329;
wire var330;
wire var331;
wire var332;
wire var333;
wire var334;
wire var335;
wire var336;
wire var337;
wire var338;
wire var339;
wire var340;
wire var341;
wire var342;
wire var343;
wire var344;
wire var345;
wire var346;
wire var347;
wire var348;
wire var349;
wire var350;
wire var351;
wire var352;
wire var353;
wire var354;
wire var355;
wire var356;
wire var357;
wire var358;
wire var359;
wire var360;
wire var361;
wire var362;
wire var363;
wire var364;
wire var365;
wire var366;
wire var367;
wire var368;
wire var369;
wire var370;
wire var371;
wire var372;
wire var373;
wire var374;
wire var375;
wire var376;
wire var377;
wire var378;
wire var379;
wire var380;
wire var381;
wire var382;
wire var383;
wire var384;
wire var385;
wire var386;
wire var387;
wire var388;
wire var389;
wire var390;
wire var391;
wire var392;
wire var393;
wire var394;
wire var395;
wire var396;
wire var397;
wire var398;
wire var399;
wire var400;
wire var401;
wire var402;
wire var403;
wire var404;
wire var405;
wire var406;
wire var407;
wire var408;
wire var409;
wire var410;
wire var411;
wire var412;
wire var413;
wire var414;
wire var415;
wire var416;
wire var417;
wire var418;
wire var419;
wire var420;
wire var421;
wire var422;
wire var423;
wire var424;
wire var425;
wire var426;
wire var427;
wire var428;
wire var429;
wire var430;
wire var431;
wire var432;
wire var433;
wire var434;
wire var435;
wire var436;
wire var437;
wire var438;
wire var439;
wire var440;
wire var441;
wire var442;
wire var443;
wire var444;
wire var445;
wire var446;
wire var447;
wire var448;
wire var449;
wire var450;
wire var451;
wire var452;
wire var453;
wire var454;
wire var455;
wire var456;
wire var457;
wire var458;
wire var459;
wire var460;
wire var461;
wire var462;
wire var463;
wire var464;
wire var465;
wire var466;
wire var467;
wire var468;
wire var469;
wire var470;
wire var471;
wire var472;
wire var473;
wire var474;
wire var475;
wire var476;
wire var477;
wire var478;
wire var479;
wire var480;
wire var481;
wire var482;
wire var483;
wire var484;
wire var485;
wire var486;
wire var487;
wire var488;
wire var489;
wire var490;
wire var491;
wire var492;
wire var493;
wire var494;
wire var495;
wire var496;
wire var497;
wire var498;
wire var499;
wire var500;
wire var501;
wire var502;
wire var503;
wire var504;
wire var505;
wire var506;
wire var507;
wire var508;
wire var509;
wire var510;
wire var511;
wire var512;
wire var513;
wire var514;
wire var515;
wire var516;
wire var517;
wire var518;
wire var519;
wire var520;
wire var521;
wire var522;
wire var523;
wire var524;
wire var525;
wire var526;
wire var527;
wire var528;
wire var529;
wire var530;
wire var531;
wire var532;
wire var533;
wire var534;
wire var535;
wire var536;
wire var537;
wire var538;
wire var539;
wire var540;
wire var541;
wire var542;
wire var543;
wire var544;
wire var545;
wire var546;
wire var547;
wire var548;
wire var549;
wire var550;
wire var551;
wire var552;
wire var553;
wire var554;
wire var555;
wire var556;
wire var557;
wire var558;
wire var559;
wire var560;
wire var561;
wire var562;
wire var563;
wire var564;
wire var565;
wire var566;
wire var567;
wire var568;
wire var569;
wire var570;
wire var571;
wire var572;
wire var573;
wire var574;
wire var575;
wire var576;
wire var577;
wire var578;
wire var579;
wire var580;
wire var581;
wire var582;
wire var583;
wire var584;
wire var585;
wire var586;
wire var587;
wire var588;
wire var589;
wire var590;
wire var591;
wire var592;
wire var593;
wire var594;
wire var595;
wire var596;
wire var597;
wire var598;
wire var599;
wire var600;
wire var601;
wire var602;
wire var603;
wire var604;
wire var605;
wire var606;
wire var607;
wire var608;
wire var609;
wire var610;
wire var611;
wire var612;
wire var613;
wire var614;
wire var615;
wire var616;
wire var617;
wire var618;
wire var619;
wire var620;
wire var621;
wire var622;
wire var623;
wire var624;
wire var625;
wire var626;
wire var627;
wire var628;
wire var629;
wire var630;
wire var631;
wire var632;
wire var633;
wire var634;
wire var635;
wire var636;
wire var637;
wire var638;
wire var639;
wire var640;
wire var641;
wire var642;
wire var643;
wire var644;
wire var645;
wire var646;
wire var647;
wire var648;
wire var649;
wire var650;
wire var651;
wire var652;
wire var653;
wire var654;
wire var655;
wire var656;
wire var657;
wire var658;
wire var659;
wire var660;
wire var661;
wire var662;
wire var663;
wire var664;
wire var665;
wire var666;
wire var667;
wire var668;
wire var669;
wire var670;
wire var671;
wire var672;
wire var673;
wire var674;
wire var675;
wire var676;
wire var677;
wire var678;
wire var679;
wire var680;
wire var681;
wire var682;
wire var683;
wire var684;
wire var685;
wire var686;
wire var687;
wire var688;
wire var689;
wire var690;
wire var691;
wire var692;
wire var693;
wire var694;
wire var695;
wire var696;
wire var697;
wire var698;
wire var699;
wire var700;
wire var701;
wire var702;
wire var703;
wire var704;
wire var705;
wire var706;
wire var707;
wire var708;
wire var709;
wire var710;
wire var711;
wire var712;
wire var713;
wire var714;
wire var715;
wire var716;
wire var717;
wire var718;
wire var719;
wire var720;
wire var721;
wire var722;
wire var723;
wire var724;
wire var725;
wire var726;
wire var727;
wire var728;
wire var729;
wire var730;
wire var731;
wire var732;
wire var733;
wire var734;
wire var735;
wire var736;
wire var737;
wire var738;
wire var739;
wire var740;
wire var741;
wire var742;
wire var743;
wire var744;
wire var745;
wire var746;
wire var747;
wire var748;
wire var749;
wire var750;
wire var751;
wire var752;
wire var753;
wire var754;
wire var755;
wire var756;
wire var757;
wire var758;
wire var759;
wire var760;
wire var761;
wire var762;
wire var763;
wire var764;
wire var765;
wire var766;
wire var767;
wire var768;
wire var769;
wire var770;
wire var771;
wire var772;
wire var773;
wire var774;
wire var775;
wire var776;
wire var777;
wire var778;
wire var779;
wire var780;
wire var781;
wire var782;
wire var783;
wire var784;
wire var785;
wire var786;
wire var787;
wire var788;
wire var789;
wire var790;
wire var791;
wire var792;
wire var793;
wire var794;
wire var795;
wire var796;
wire var797;
wire var798;
wire var799;
wire var800;
wire var801;
wire var802;
wire var803;
wire var804;
wire var805;
wire var806;
wire var807;
wire var808;
wire var809;
wire var810;
wire var811;
wire var812;
wire var813;
wire var814;
wire var815;
wire var816;
wire var817;
wire var818;
wire var819;
wire var820;
wire var821;
wire var822;
wire var823;
wire var824;
wire var825;
wire var826;
wire var827;
wire var828;
wire var829;
wire var830;
wire var831;
wire var832;
wire var833;
wire var834;
wire var835;
wire var836;
wire var837;
wire var838;
wire var839;
wire var840;
wire var841;
wire var842;
wire var843;
wire var844;
wire var845;
wire var846;
wire var847;
wire var848;
wire var849;
wire var850;
wire var851;
wire var852;
wire var853;
wire var854;
wire var855;
wire var856;
wire var857;
wire var858;
wire var859;
wire var860;
wire var861;
wire var862;
wire var863;
wire var864;
wire var865;
wire var866;
wire var867;
wire var868;
wire var869;
wire var870;
wire var871;
wire var872;
wire var873;
wire var874;
wire var875;
wire var876;
wire var877;
wire var878;
wire var879;
wire var880;
wire var881;
wire var882;
wire var883;
wire var884;
wire var885;
wire var886;
wire var887;
wire var888;
wire var889;
wire var890;
wire var891;
wire var892;
wire var893;
wire var894;
wire var895;
wire var896;
wire var897;
wire var898;
wire var899;
wire var900;
wire var901;
wire var902;
wire var903;
wire var904;
wire var905;
wire var906;
wire var907;
wire var908;
wire var909;
wire var910;
wire var911;
wire var912;
wire var913;
wire var914;
wire var915;
wire var916;
wire var917;
wire var918;
wire var919;
wire var920;
wire var921;
wire var922;
wire var923;
wire var924;
wire var925;
wire var926;
wire var927;
wire var928;
wire var929;
wire var930;
wire var931;
wire var932;
wire var933;
wire var934;
wire var935;
wire var936;
wire var937;
wire var938;
wire var939;
wire var940;
wire var941;
wire var942;
wire var943;
wire var944;
wire var945;
wire var946;
wire var947;
wire var948;
wire var949;
wire var950;
wire var951;
wire var952;
wire var953;
wire var954;
wire var955;
wire var956;
wire var957;
wire var958;
wire var959;
wire var960;
wire var961;
wire var962;
wire var963;
wire var964;
wire var965;
wire var966;
wire var967;
wire var968;
wire var969;
wire var970;
wire var971;
wire var972;
wire var973;
wire var974;
wire var975;
wire var976;
wire var977;
wire var978;
wire var979;
wire var980;
wire var981;
wire var982;
wire var983;
wire var984;
wire var985;
wire var986;
wire var987;
wire var988;
wire var989;
wire var990;
wire var991;
wire var992;
wire var993;
wire var994;
wire var995;
wire var996;
wire var997;
wire var998;
wire var999;
wire var1000;
wire var1001;
wire var1002;
wire var1003;
wire var1004;
wire var1005;
wire var1006;
wire var1007;
wire var1008;
wire var1009;
wire var1010;
wire var1011;
wire var1012;
wire var1013;
wire var1014;
wire var1015;
wire var1016;
wire var1017;
wire var1018;
wire var1019;
wire var1020;
wire var1021;
wire var1022;
wire var1023;
wire var1024;
wire var1025;
wire var1026;
wire var1027;
wire var1028;
wire var1029;
wire var1030;
wire var1031;
wire var1032;
wire var1033;
wire var1034;
wire var1035;
wire var1036;
wire var1037;
wire var1038;
wire var1039;
wire var1040;
wire var1041;
wire var1042;
wire var1043;
wire var1044;
wire var1045;
wire var1046;
wire var1047;
wire var1048;
wire var1049;
wire var1050;
wire var1051;
wire var1052;
wire var1053;
wire var1054;
wire var1055;
wire var1056;
wire var1057;
wire var1058;
wire var1059;
wire var1060;
wire var1061;
wire var1062;
wire var1063;
wire var1064;
wire var1065;
wire var1066;
wire var1067;
wire var1068;
wire var1069;
wire var1070;
wire var1071;
wire var1072;
wire var1073;
wire var1074;
wire var1075;
wire var1076;
wire var1077;
wire var1078;
wire var1079;
wire var1080;
wire var1081;
wire var1082;
wire var1083;
wire var1084;
wire var1085;
wire var1086;
wire var1087;
wire var1088;
wire var1089;
wire var1090;
assign var0 = in127 & in63;
assign var1 = in126 & in62;
assign var2 = in125 & in61;
assign var3 = in124 & in60;
assign var4 = in123 & in59;
assign var5 = in122 & in58;
assign var6 = in121 & in57;
assign var7 = in120 & in56;
assign var8 = in119 & in55;
assign var9 = in118 & in54;
assign var10 = in117 & in53;
assign var11 = in116 & in52;
assign var12 = in115 & in51;
assign var13 = in114 & in50;
assign var14 = in113 & in49;
assign var15 = in112 & in48;
assign var16 = in111 & in47;
assign var17 = in110 & in46;
assign var18 = in109 & in45;
assign var19 = in108 & in44;
assign var20 = in107 & in43;
assign var21 = in106 & in42;
assign var22 = in105 & in41;
assign var23 = in104 & in40;
assign var24 = in103 & in39;
assign var25 = in102 & in38;
assign var26 = in101 & in37;
assign var27 = in100 & in36;
assign var28 = in99 & in35;
assign var29 = in98 & in34;
assign var30 = in97 & in33;
assign var31 = in96 & in32;
assign var32 = in95 & in31;
assign var33 = in94 & in30;
assign var34 = in93 & in29;
assign var35 = in92 & in28;
assign var36 = in91 & in27;
assign var37 = in90 & in26;
assign var38 = in89 & in25;
assign var39 = in88 & in24;
assign var40 = in87 & in23;
assign var41 = in86 & in22;
assign var42 = in85 & in21;
assign var43 = in84 & in20;
assign var44 = in83 & in19;
assign var45 = in82 & in18;
assign var46 = in81 & in17;
assign var47 = in80 & in16;
assign var48 = in79 & in15;
assign var49 = in78 & in14;
assign var50 = in77 & in13;
assign var51 = in76 & in12;
assign var52 = in75 & in11;
assign var53 = in74 & in10;
assign var54 = in73 & in9;
assign var55 = in72 & in8;
assign var56 = in71 & in7;
assign var57 = in70 & in6;
assign var58 = in69 & in5;
assign var59 = in68 & in4;
assign var60 = in67 & in3;
assign var61 = in66 & in2;
assign var62 = in65 & in1;
assign var63 = in64 & in0;
assign var64 = in127 ^ in63;
assign var65 = in126 ^ in62;
assign var66 = in125 ^ in61;
assign var67 = in124 ^ in60;
assign var68 = in123 ^ in59;
assign var69 = in122 ^ in58;
assign var70 = in121 ^ in57;
assign var71 = in120 ^ in56;
assign var72 = in119 ^ in55;
assign var73 = in118 ^ in54;
assign var74 = in117 ^ in53;
assign var75 = in116 ^ in52;
assign var76 = in115 ^ in51;
assign var77 = in114 ^ in50;
assign var78 = in113 ^ in49;
assign var79 = in112 ^ in48;
assign var80 = in111 ^ in47;
assign var81 = in110 ^ in46;
assign var82 = in109 ^ in45;
assign var83 = in108 ^ in44;
assign var84 = in107 ^ in43;
assign var85 = in106 ^ in42;
assign var86 = in105 ^ in41;
assign var87 = in104 ^ in40;
assign var88 = in103 ^ in39;
assign var89 = in102 ^ in38;
assign var90 = in101 ^ in37;
assign var91 = in100 ^ in36;
assign var92 = in99 ^ in35;
assign var93 = in98 ^ in34;
assign var94 = in97 ^ in33;
assign var95 = in96 ^ in32;
assign var96 = in95 ^ in31;
assign var97 = in94 ^ in30;
assign var98 = in93 ^ in29;
assign var99 = in92 ^ in28;
assign var100 = in91 ^ in27;
assign var101 = in90 ^ in26;
assign var102 = in89 ^ in25;
assign var103 = in88 ^ in24;
assign var104 = in87 ^ in23;
assign var105 = in86 ^ in22;
assign var106 = in85 ^ in21;
assign var107 = in84 ^ in20;
assign var108 = in83 ^ in19;
assign var109 = in82 ^ in18;
assign var110 = in81 ^ in17;
assign var111 = in80 ^ in16;
assign var112 = in79 ^ in15;
assign var113 = in78 ^ in14;
assign var114 = in77 ^ in13;
assign var115 = in76 ^ in12;
assign var116 = in75 ^ in11;
assign var117 = in74 ^ in10;
assign var118 = in73 ^ in9;
assign var119 = in72 ^ in8;
assign var120 = in71 ^ in7;
assign var121 = in70 ^ in6;
assign var122 = in69 ^ in5;
assign var123 = in68 ^ in4;
assign var124 = in67 ^ in3;
assign var125 = in66 ^ in2;
assign var126 = in65 ^ in1;
assign var127 = in64 ^ in0;
assign var128 = var127 & var62;
assign var129 = var63 | var128;
assign var130 = var127 & var126;
assign var131 = var126 & var61;
assign var132 = var62 | var131;
assign var133 = var126 & var125;
assign var134 = var125 & var60;
assign var135 = var61 | var134;
assign var136 = var125 & var124;
assign var137 = var124 & var59;
assign var138 = var60 | var137;
assign var139 = var124 & var123;
assign var140 = var123 & var58;
assign var141 = var59 | var140;
assign var142 = var123 & var122;
assign var143 = var122 & var57;
assign var144 = var58 | var143;
assign var145 = var122 & var121;
assign var146 = var121 & var56;
assign var147 = var57 | var146;
assign var148 = var121 & var120;
assign var149 = var120 & var55;
assign var150 = var56 | var149;
assign var151 = var120 & var119;
assign var152 = var119 & var54;
assign var153 = var55 | var152;
assign var154 = var119 & var118;
assign var155 = var118 & var53;
assign var156 = var54 | var155;
assign var157 = var118 & var117;
assign var158 = var117 & var52;
assign var159 = var53 | var158;
assign var160 = var117 & var116;
assign var161 = var116 & var51;
assign var162 = var52 | var161;
assign var163 = var116 & var115;
assign var164 = var115 & var50;
assign var165 = var51 | var164;
assign var166 = var115 & var114;
assign var167 = var114 & var49;
assign var168 = var50 | var167;
assign var169 = var114 & var113;
assign var170 = var113 & var48;
assign var171 = var49 | var170;
assign var172 = var113 & var112;
assign var173 = var112 & var47;
assign var174 = var48 | var173;
assign var175 = var112 & var111;
assign var176 = var111 & var46;
assign var177 = var47 | var176;
assign var178 = var111 & var110;
assign var179 = var110 & var45;
assign var180 = var46 | var179;
assign var181 = var110 & var109;
assign var182 = var109 & var44;
assign var183 = var45 | var182;
assign var184 = var109 & var108;
assign var185 = var108 & var43;
assign var186 = var44 | var185;
assign var187 = var108 & var107;
assign var188 = var107 & var42;
assign var189 = var43 | var188;
assign var190 = var107 & var106;
assign var191 = var106 & var41;
assign var192 = var42 | var191;
assign var193 = var106 & var105;
assign var194 = var105 & var40;
assign var195 = var41 | var194;
assign var196 = var105 & var104;
assign var197 = var104 & var39;
assign var198 = var40 | var197;
assign var199 = var104 & var103;
assign var200 = var103 & var38;
assign var201 = var39 | var200;
assign var202 = var103 & var102;
assign var203 = var102 & var37;
assign var204 = var38 | var203;
assign var205 = var102 & var101;
assign var206 = var101 & var36;
assign var207 = var37 | var206;
assign var208 = var101 & var100;
assign var209 = var100 & var35;
assign var210 = var36 | var209;
assign var211 = var100 & var99;
assign var212 = var99 & var34;
assign var213 = var35 | var212;
assign var214 = var99 & var98;
assign var215 = var98 & var33;
assign var216 = var34 | var215;
assign var217 = var98 & var97;
assign var218 = var97 & var32;
assign var219 = var33 | var218;
assign var220 = var97 & var96;
assign var221 = var96 & var31;
assign var222 = var32 | var221;
assign var223 = var96 & var95;
assign var224 = var95 & var30;
assign var225 = var31 | var224;
assign var226 = var95 & var94;
assign var227 = var94 & var29;
assign var228 = var30 | var227;
assign var229 = var94 & var93;
assign var230 = var93 & var28;
assign var231 = var29 | var230;
assign var232 = var93 & var92;
assign var233 = var92 & var27;
assign var234 = var28 | var233;
assign var235 = var92 & var91;
assign var236 = var91 & var26;
assign var237 = var27 | var236;
assign var238 = var91 & var90;
assign var239 = var90 & var25;
assign var240 = var26 | var239;
assign var241 = var90 & var89;
assign var242 = var89 & var24;
assign var243 = var25 | var242;
assign var244 = var89 & var88;
assign var245 = var88 & var23;
assign var246 = var24 | var245;
assign var247 = var88 & var87;
assign var248 = var87 & var22;
assign var249 = var23 | var248;
assign var250 = var87 & var86;
assign var251 = var86 & var21;
assign var252 = var22 | var251;
assign var253 = var86 & var85;
assign var254 = var85 & var20;
assign var255 = var21 | var254;
assign var256 = var85 & var84;
assign var257 = var84 & var19;
assign var258 = var20 | var257;
assign var259 = var84 & var83;
assign var260 = var83 & var18;
assign var261 = var19 | var260;
assign var262 = var83 & var82;
assign var263 = var82 & var17;
assign var264 = var18 | var263;
assign var265 = var82 & var81;
assign var266 = var81 & var16;
assign var267 = var17 | var266;
assign var268 = var81 & var80;
assign var269 = var80 & var15;
assign var270 = var16 | var269;
assign var271 = var80 & var79;
assign var272 = var79 & var14;
assign var273 = var15 | var272;
assign var274 = var79 & var78;
assign var275 = var78 & var13;
assign var276 = var14 | var275;
assign var277 = var78 & var77;
assign var278 = var77 & var12;
assign var279 = var13 | var278;
assign var280 = var77 & var76;
assign var281 = var76 & var11;
assign var282 = var12 | var281;
assign var283 = var76 & var75;
assign var284 = var75 & var10;
assign var285 = var11 | var284;
assign var286 = var75 & var74;
assign var287 = var74 & var9;
assign var288 = var10 | var287;
assign var289 = var74 & var73;
assign var290 = var73 & var8;
assign var291 = var9 | var290;
assign var292 = var73 & var72;
assign var293 = var72 & var7;
assign var294 = var8 | var293;
assign var295 = var72 & var71;
assign var296 = var71 & var6;
assign var297 = var7 | var296;
assign var298 = var71 & var70;
assign var299 = var70 & var5;
assign var300 = var6 | var299;
assign var301 = var70 & var69;
assign var302 = var69 & var4;
assign var303 = var5 | var302;
assign var304 = var69 & var68;
assign var305 = var68 & var3;
assign var306 = var4 | var305;
assign var307 = var68 & var67;
assign var308 = var67 & var2;
assign var309 = var3 | var308;
assign var310 = var67 & var66;
assign var311 = var66 & var1;
assign var312 = var2 | var311;
assign var313 = var66 & var65;
assign var314 = var65 & var0;
assign var315 = var1 | var314;
assign var316 = var130 & var135;
assign var317 = var129 | var316;
assign var318 = var130 & var136;
assign var319 = var133 & var138;
assign var320 = var132 | var319;
assign var321 = var133 & var139;
assign var322 = var136 & var141;
assign var323 = var135 | var322;
assign var324 = var136 & var142;
assign var325 = var139 & var144;
assign var326 = var138 | var325;
assign var327 = var139 & var145;
assign var328 = var142 & var147;
assign var329 = var141 | var328;
assign var330 = var142 & var148;
assign var331 = var145 & var150;
assign var332 = var144 | var331;
assign var333 = var145 & var151;
assign var334 = var148 & var153;
assign var335 = var147 | var334;
assign var336 = var148 & var154;
assign var337 = var151 & var156;
assign var338 = var150 | var337;
assign var339 = var151 & var157;
assign var340 = var154 & var159;
assign var341 = var153 | var340;
assign var342 = var154 & var160;
assign var343 = var157 & var162;
assign var344 = var156 | var343;
assign var345 = var157 & var163;
assign var346 = var160 & var165;
assign var347 = var159 | var346;
assign var348 = var160 & var166;
assign var349 = var163 & var168;
assign var350 = var162 | var349;
assign var351 = var163 & var169;
assign var352 = var166 & var171;
assign var353 = var165 | var352;
assign var354 = var166 & var172;
assign var355 = var169 & var174;
assign var356 = var168 | var355;
assign var357 = var169 & var175;
assign var358 = var172 & var177;
assign var359 = var171 | var358;
assign var360 = var172 & var178;
assign var361 = var175 & var180;
assign var362 = var174 | var361;
assign var363 = var175 & var181;
assign var364 = var178 & var183;
assign var365 = var177 | var364;
assign var366 = var178 & var184;
assign var367 = var181 & var186;
assign var368 = var180 | var367;
assign var369 = var181 & var187;
assign var370 = var184 & var189;
assign var371 = var183 | var370;
assign var372 = var184 & var190;
assign var373 = var187 & var192;
assign var374 = var186 | var373;
assign var375 = var187 & var193;
assign var376 = var190 & var195;
assign var377 = var189 | var376;
assign var378 = var190 & var196;
assign var379 = var193 & var198;
assign var380 = var192 | var379;
assign var381 = var193 & var199;
assign var382 = var196 & var201;
assign var383 = var195 | var382;
assign var384 = var196 & var202;
assign var385 = var199 & var204;
assign var386 = var198 | var385;
assign var387 = var199 & var205;
assign var388 = var202 & var207;
assign var389 = var201 | var388;
assign var390 = var202 & var208;
assign var391 = var205 & var210;
assign var392 = var204 | var391;
assign var393 = var205 & var211;
assign var394 = var208 & var213;
assign var395 = var207 | var394;
assign var396 = var208 & var214;
assign var397 = var211 & var216;
assign var398 = var210 | var397;
assign var399 = var211 & var217;
assign var400 = var214 & var219;
assign var401 = var213 | var400;
assign var402 = var214 & var220;
assign var403 = var217 & var222;
assign var404 = var216 | var403;
assign var405 = var217 & var223;
assign var406 = var220 & var225;
assign var407 = var219 | var406;
assign var408 = var220 & var226;
assign var409 = var223 & var228;
assign var410 = var222 | var409;
assign var411 = var223 & var229;
assign var412 = var226 & var231;
assign var413 = var225 | var412;
assign var414 = var226 & var232;
assign var415 = var229 & var234;
assign var416 = var228 | var415;
assign var417 = var229 & var235;
assign var418 = var232 & var237;
assign var419 = var231 | var418;
assign var420 = var232 & var238;
assign var421 = var235 & var240;
assign var422 = var234 | var421;
assign var423 = var235 & var241;
assign var424 = var238 & var243;
assign var425 = var237 | var424;
assign var426 = var238 & var244;
assign var427 = var241 & var246;
assign var428 = var240 | var427;
assign var429 = var241 & var247;
assign var430 = var244 & var249;
assign var431 = var243 | var430;
assign var432 = var244 & var250;
assign var433 = var247 & var252;
assign var434 = var246 | var433;
assign var435 = var247 & var253;
assign var436 = var250 & var255;
assign var437 = var249 | var436;
assign var438 = var250 & var256;
assign var439 = var253 & var258;
assign var440 = var252 | var439;
assign var441 = var253 & var259;
assign var442 = var256 & var261;
assign var443 = var255 | var442;
assign var444 = var256 & var262;
assign var445 = var259 & var264;
assign var446 = var258 | var445;
assign var447 = var259 & var265;
assign var448 = var262 & var267;
assign var449 = var261 | var448;
assign var450 = var262 & var268;
assign var451 = var265 & var270;
assign var452 = var264 | var451;
assign var453 = var265 & var271;
assign var454 = var268 & var273;
assign var455 = var267 | var454;
assign var456 = var268 & var274;
assign var457 = var271 & var276;
assign var458 = var270 | var457;
assign var459 = var271 & var277;
assign var460 = var274 & var279;
assign var461 = var273 | var460;
assign var462 = var274 & var280;
assign var463 = var277 & var282;
assign var464 = var276 | var463;
assign var465 = var277 & var283;
assign var466 = var280 & var285;
assign var467 = var279 | var466;
assign var468 = var280 & var286;
assign var469 = var283 & var288;
assign var470 = var282 | var469;
assign var471 = var283 & var289;
assign var472 = var286 & var291;
assign var473 = var285 | var472;
assign var474 = var286 & var292;
assign var475 = var289 & var294;
assign var476 = var288 | var475;
assign var477 = var289 & var295;
assign var478 = var292 & var297;
assign var479 = var291 | var478;
assign var480 = var292 & var298;
assign var481 = var295 & var300;
assign var482 = var294 | var481;
assign var483 = var295 & var301;
assign var484 = var298 & var303;
assign var485 = var297 | var484;
assign var486 = var298 & var304;
assign var487 = var301 & var306;
assign var488 = var300 | var487;
assign var489 = var301 & var307;
assign var490 = var304 & var309;
assign var491 = var303 | var490;
assign var492 = var304 & var310;
assign var493 = var307 & var312;
assign var494 = var306 | var493;
assign var495 = var307 & var313;
assign var496 = var310 & var315;
assign var497 = var309 | var496;
assign var498 = var313 & var0;
assign var499 = var312 | var498;
assign var500 = var318 & var329;
assign var501 = var317 | var500;
assign var502 = var318 & var330;
assign var503 = var321 & var332;
assign var504 = var320 | var503;
assign var505 = var321 & var333;
assign var506 = var324 & var335;
assign var507 = var323 | var506;
assign var508 = var324 & var336;
assign var509 = var327 & var338;
assign var510 = var326 | var509;
assign var511 = var327 & var339;
assign var512 = var330 & var341;
assign var513 = var329 | var512;
assign var514 = var330 & var342;
assign var515 = var333 & var344;
assign var516 = var332 | var515;
assign var517 = var333 & var345;
assign var518 = var336 & var347;
assign var519 = var335 | var518;
assign var520 = var336 & var348;
assign var521 = var339 & var350;
assign var522 = var338 | var521;
assign var523 = var339 & var351;
assign var524 = var342 & var353;
assign var525 = var341 | var524;
assign var526 = var342 & var354;
assign var527 = var345 & var356;
assign var528 = var344 | var527;
assign var529 = var345 & var357;
assign var530 = var348 & var359;
assign var531 = var347 | var530;
assign var532 = var348 & var360;
assign var533 = var351 & var362;
assign var534 = var350 | var533;
assign var535 = var351 & var363;
assign var536 = var354 & var365;
assign var537 = var353 | var536;
assign var538 = var354 & var366;
assign var539 = var357 & var368;
assign var540 = var356 | var539;
assign var541 = var357 & var369;
assign var542 = var360 & var371;
assign var543 = var359 | var542;
assign var544 = var360 & var372;
assign var545 = var363 & var374;
assign var546 = var362 | var545;
assign var547 = var363 & var375;
assign var548 = var366 & var377;
assign var549 = var365 | var548;
assign var550 = var366 & var378;
assign var551 = var369 & var380;
assign var552 = var368 | var551;
assign var553 = var369 & var381;
assign var554 = var372 & var383;
assign var555 = var371 | var554;
assign var556 = var372 & var384;
assign var557 = var375 & var386;
assign var558 = var374 | var557;
assign var559 = var375 & var387;
assign var560 = var378 & var389;
assign var561 = var377 | var560;
assign var562 = var378 & var390;
assign var563 = var381 & var392;
assign var564 = var380 | var563;
assign var565 = var381 & var393;
assign var566 = var384 & var395;
assign var567 = var383 | var566;
assign var568 = var384 & var396;
assign var569 = var387 & var398;
assign var570 = var386 | var569;
assign var571 = var387 & var399;
assign var572 = var390 & var401;
assign var573 = var389 | var572;
assign var574 = var390 & var402;
assign var575 = var393 & var404;
assign var576 = var392 | var575;
assign var577 = var393 & var405;
assign var578 = var396 & var407;
assign var579 = var395 | var578;
assign var580 = var396 & var408;
assign var581 = var399 & var410;
assign var582 = var398 | var581;
assign var583 = var399 & var411;
assign var584 = var402 & var413;
assign var585 = var401 | var584;
assign var586 = var402 & var414;
assign var587 = var405 & var416;
assign var588 = var404 | var587;
assign var589 = var405 & var417;
assign var590 = var408 & var419;
assign var591 = var407 | var590;
assign var592 = var408 & var420;
assign var593 = var411 & var422;
assign var594 = var410 | var593;
assign var595 = var411 & var423;
assign var596 = var414 & var425;
assign var597 = var413 | var596;
assign var598 = var414 & var426;
assign var599 = var417 & var428;
assign var600 = var416 | var599;
assign var601 = var417 & var429;
assign var602 = var420 & var431;
assign var603 = var419 | var602;
assign var604 = var420 & var432;
assign var605 = var423 & var434;
assign var606 = var422 | var605;
assign var607 = var423 & var435;
assign var608 = var426 & var437;
assign var609 = var425 | var608;
assign var610 = var426 & var438;
assign var611 = var429 & var440;
assign var612 = var428 | var611;
assign var613 = var429 & var441;
assign var614 = var432 & var443;
assign var615 = var431 | var614;
assign var616 = var432 & var444;
assign var617 = var435 & var446;
assign var618 = var434 | var617;
assign var619 = var435 & var447;
assign var620 = var438 & var449;
assign var621 = var437 | var620;
assign var622 = var438 & var450;
assign var623 = var441 & var452;
assign var624 = var440 | var623;
assign var625 = var441 & var453;
assign var626 = var444 & var455;
assign var627 = var443 | var626;
assign var628 = var444 & var456;
assign var629 = var447 & var458;
assign var630 = var446 | var629;
assign var631 = var447 & var459;
assign var632 = var450 & var461;
assign var633 = var449 | var632;
assign var634 = var450 & var462;
assign var635 = var453 & var464;
assign var636 = var452 | var635;
assign var637 = var453 & var465;
assign var638 = var456 & var467;
assign var639 = var455 | var638;
assign var640 = var456 & var468;
assign var641 = var459 & var470;
assign var642 = var458 | var641;
assign var643 = var459 & var471;
assign var644 = var462 & var473;
assign var645 = var461 | var644;
assign var646 = var462 & var474;
assign var647 = var465 & var476;
assign var648 = var464 | var647;
assign var649 = var465 & var477;
assign var650 = var468 & var479;
assign var651 = var467 | var650;
assign var652 = var468 & var480;
assign var653 = var471 & var482;
assign var654 = var470 | var653;
assign var655 = var471 & var483;
assign var656 = var474 & var485;
assign var657 = var473 | var656;
assign var658 = var474 & var486;
assign var659 = var477 & var488;
assign var660 = var476 | var659;
assign var661 = var477 & var489;
assign var662 = var480 & var491;
assign var663 = var479 | var662;
assign var664 = var480 & var492;
assign var665 = var483 & var494;
assign var666 = var482 | var665;
assign var667 = var483 & var495;
assign var668 = var486 & var497;
assign var669 = var485 | var668;
assign var670 = var489 & var499;
assign var671 = var488 | var670;
assign var672 = var492 & var315;
assign var673 = var491 | var672;
assign var674 = var495 & var0;
assign var675 = var494 | var674;
assign var676 = var502 & var525;
assign var677 = var501 | var676;
assign var678 = var502 & var526;
assign var679 = var505 & var528;
assign var680 = var504 | var679;
assign var681 = var505 & var529;
assign var682 = var508 & var531;
assign var683 = var507 | var682;
assign var684 = var508 & var532;
assign var685 = var511 & var534;
assign var686 = var510 | var685;
assign var687 = var511 & var535;
assign var688 = var514 & var537;
assign var689 = var513 | var688;
assign var690 = var514 & var538;
assign var691 = var517 & var540;
assign var692 = var516 | var691;
assign var693 = var517 & var541;
assign var694 = var520 & var543;
assign var695 = var519 | var694;
assign var696 = var520 & var544;
assign var697 = var523 & var546;
assign var698 = var522 | var697;
assign var699 = var523 & var547;
assign var700 = var526 & var549;
assign var701 = var525 | var700;
assign var702 = var526 & var550;
assign var703 = var529 & var552;
assign var704 = var528 | var703;
assign var705 = var529 & var553;
assign var706 = var532 & var555;
assign var707 = var531 | var706;
assign var708 = var532 & var556;
assign var709 = var535 & var558;
assign var710 = var534 | var709;
assign var711 = var535 & var559;
assign var712 = var538 & var561;
assign var713 = var537 | var712;
assign var714 = var538 & var562;
assign var715 = var541 & var564;
assign var716 = var540 | var715;
assign var717 = var541 & var565;
assign var718 = var544 & var567;
assign var719 = var543 | var718;
assign var720 = var544 & var568;
assign var721 = var547 & var570;
assign var722 = var546 | var721;
assign var723 = var547 & var571;
assign var724 = var550 & var573;
assign var725 = var549 | var724;
assign var726 = var550 & var574;
assign var727 = var553 & var576;
assign var728 = var552 | var727;
assign var729 = var553 & var577;
assign var730 = var556 & var579;
assign var731 = var555 | var730;
assign var732 = var556 & var580;
assign var733 = var559 & var582;
assign var734 = var558 | var733;
assign var735 = var559 & var583;
assign var736 = var562 & var585;
assign var737 = var561 | var736;
assign var738 = var562 & var586;
assign var739 = var565 & var588;
assign var740 = var564 | var739;
assign var741 = var565 & var589;
assign var742 = var568 & var591;
assign var743 = var567 | var742;
assign var744 = var568 & var592;
assign var745 = var571 & var594;
assign var746 = var570 | var745;
assign var747 = var571 & var595;
assign var748 = var574 & var597;
assign var749 = var573 | var748;
assign var750 = var574 & var598;
assign var751 = var577 & var600;
assign var752 = var576 | var751;
assign var753 = var577 & var601;
assign var754 = var580 & var603;
assign var755 = var579 | var754;
assign var756 = var580 & var604;
assign var757 = var583 & var606;
assign var758 = var582 | var757;
assign var759 = var583 & var607;
assign var760 = var586 & var609;
assign var761 = var585 | var760;
assign var762 = var586 & var610;
assign var763 = var589 & var612;
assign var764 = var588 | var763;
assign var765 = var589 & var613;
assign var766 = var592 & var615;
assign var767 = var591 | var766;
assign var768 = var592 & var616;
assign var769 = var595 & var618;
assign var770 = var594 | var769;
assign var771 = var595 & var619;
assign var772 = var598 & var621;
assign var773 = var597 | var772;
assign var774 = var598 & var622;
assign var775 = var601 & var624;
assign var776 = var600 | var775;
assign var777 = var601 & var625;
assign var778 = var604 & var627;
assign var779 = var603 | var778;
assign var780 = var604 & var628;
assign var781 = var607 & var630;
assign var782 = var606 | var781;
assign var783 = var607 & var631;
assign var784 = var610 & var633;
assign var785 = var609 | var784;
assign var786 = var610 & var634;
assign var787 = var613 & var636;
assign var788 = var612 | var787;
assign var789 = var613 & var637;
assign var790 = var616 & var639;
assign var791 = var615 | var790;
assign var792 = var616 & var640;
assign var793 = var619 & var642;
assign var794 = var618 | var793;
assign var795 = var619 & var643;
assign var796 = var622 & var645;
assign var797 = var621 | var796;
assign var798 = var622 & var646;
assign var799 = var625 & var648;
assign var800 = var624 | var799;
assign var801 = var625 & var649;
assign var802 = var628 & var651;
assign var803 = var627 | var802;
assign var804 = var628 & var652;
assign var805 = var631 & var654;
assign var806 = var630 | var805;
assign var807 = var631 & var655;
assign var808 = var634 & var657;
assign var809 = var633 | var808;
assign var810 = var634 & var658;
assign var811 = var637 & var660;
assign var812 = var636 | var811;
assign var813 = var637 & var661;
assign var814 = var640 & var663;
assign var815 = var639 | var814;
assign var816 = var640 & var664;
assign var817 = var643 & var666;
assign var818 = var642 | var817;
assign var819 = var643 & var667;
assign var820 = var646 & var669;
assign var821 = var645 | var820;
assign var822 = var649 & var671;
assign var823 = var648 | var822;
assign var824 = var652 & var673;
assign var825 = var651 | var824;
assign var826 = var655 & var675;
assign var827 = var654 | var826;
assign var828 = var658 & var497;
assign var829 = var657 | var828;
assign var830 = var661 & var499;
assign var831 = var660 | var830;
assign var832 = var664 & var315;
assign var833 = var663 | var832;
assign var834 = var667 & var0;
assign var835 = var666 | var834;
assign var836 = var678 & var725;
assign var837 = var677 | var836;
assign var838 = var678 & var726;
assign var839 = var681 & var728;
assign var840 = var680 | var839;
assign var841 = var681 & var729;
assign var842 = var684 & var731;
assign var843 = var683 | var842;
assign var844 = var684 & var732;
assign var845 = var687 & var734;
assign var846 = var686 | var845;
assign var847 = var687 & var735;
assign var848 = var690 & var737;
assign var849 = var689 | var848;
assign var850 = var690 & var738;
assign var851 = var693 & var740;
assign var852 = var692 | var851;
assign var853 = var693 & var741;
assign var854 = var696 & var743;
assign var855 = var695 | var854;
assign var856 = var696 & var744;
assign var857 = var699 & var746;
assign var858 = var698 | var857;
assign var859 = var699 & var747;
assign var860 = var702 & var749;
assign var861 = var701 | var860;
assign var862 = var702 & var750;
assign var863 = var705 & var752;
assign var864 = var704 | var863;
assign var865 = var705 & var753;
assign var866 = var708 & var755;
assign var867 = var707 | var866;
assign var868 = var708 & var756;
assign var869 = var711 & var758;
assign var870 = var710 | var869;
assign var871 = var711 & var759;
assign var872 = var714 & var761;
assign var873 = var713 | var872;
assign var874 = var714 & var762;
assign var875 = var717 & var764;
assign var876 = var716 | var875;
assign var877 = var717 & var765;
assign var878 = var720 & var767;
assign var879 = var719 | var878;
assign var880 = var720 & var768;
assign var881 = var723 & var770;
assign var882 = var722 | var881;
assign var883 = var723 & var771;
assign var884 = var726 & var773;
assign var885 = var725 | var884;
assign var886 = var726 & var774;
assign var887 = var729 & var776;
assign var888 = var728 | var887;
assign var889 = var729 & var777;
assign var890 = var732 & var779;
assign var891 = var731 | var890;
assign var892 = var732 & var780;
assign var893 = var735 & var782;
assign var894 = var734 | var893;
assign var895 = var735 & var783;
assign var896 = var738 & var785;
assign var897 = var737 | var896;
assign var898 = var738 & var786;
assign var899 = var741 & var788;
assign var900 = var740 | var899;
assign var901 = var741 & var789;
assign var902 = var744 & var791;
assign var903 = var743 | var902;
assign var904 = var744 & var792;
assign var905 = var747 & var794;
assign var906 = var746 | var905;
assign var907 = var747 & var795;
assign var908 = var750 & var797;
assign var909 = var749 | var908;
assign var910 = var750 & var798;
assign var911 = var753 & var800;
assign var912 = var752 | var911;
assign var913 = var753 & var801;
assign var914 = var756 & var803;
assign var915 = var755 | var914;
assign var916 = var756 & var804;
assign var917 = var759 & var806;
assign var918 = var758 | var917;
assign var919 = var759 & var807;
assign var920 = var762 & var809;
assign var921 = var761 | var920;
assign var922 = var762 & var810;
assign var923 = var765 & var812;
assign var924 = var764 | var923;
assign var925 = var765 & var813;
assign var926 = var768 & var815;
assign var927 = var767 | var926;
assign var928 = var768 & var816;
assign var929 = var771 & var818;
assign var930 = var770 | var929;
assign var931 = var771 & var819;
assign var932 = var774 & var821;
assign var933 = var773 | var932;
assign var934 = var777 & var823;
assign var935 = var776 | var934;
assign var936 = var780 & var825;
assign var937 = var779 | var936;
assign var938 = var783 & var827;
assign var939 = var782 | var938;
assign var940 = var786 & var829;
assign var941 = var785 | var940;
assign var942 = var789 & var831;
assign var943 = var788 | var942;
assign var944 = var792 & var833;
assign var945 = var791 | var944;
assign var946 = var795 & var835;
assign var947 = var794 | var946;
assign var948 = var798 & var669;
assign var949 = var797 | var948;
assign var950 = var801 & var671;
assign var951 = var800 | var950;
assign var952 = var804 & var673;
assign var953 = var803 | var952;
assign var954 = var807 & var675;
assign var955 = var806 | var954;
assign var956 = var810 & var497;
assign var957 = var809 | var956;
assign var958 = var813 & var499;
assign var959 = var812 | var958;
assign var960 = var816 & var315;
assign var961 = var815 | var960;
assign var962 = var819 & var0;
assign var963 = var818 | var962;
assign var964 = var838 & var933;
assign var965 = var837 | var964;
assign var966 = var841 & var935;
assign var967 = var840 | var966;
assign var968 = var844 & var937;
assign var969 = var843 | var968;
assign var970 = var847 & var939;
assign var971 = var846 | var970;
assign var972 = var850 & var941;
assign var973 = var849 | var972;
assign var974 = var853 & var943;
assign var975 = var852 | var974;
assign var976 = var856 & var945;
assign var977 = var855 | var976;
assign var978 = var859 & var947;
assign var979 = var858 | var978;
assign var980 = var862 & var949;
assign var981 = var861 | var980;
assign var982 = var865 & var951;
assign var983 = var864 | var982;
assign var984 = var868 & var953;
assign var985 = var867 | var984;
assign var986 = var871 & var955;
assign var987 = var870 | var986;
assign var988 = var874 & var957;
assign var989 = var873 | var988;
assign var990 = var877 & var959;
assign var991 = var876 | var990;
assign var992 = var880 & var961;
assign var993 = var879 | var992;
assign var994 = var883 & var963;
assign var995 = var882 | var994;
assign var996 = var886 & var821;
assign var997 = var885 | var996;
assign var998 = var889 & var823;
assign var999 = var888 | var998;
assign var1000 = var892 & var825;
assign var1001 = var891 | var1000;
assign var1002 = var895 & var827;
assign var1003 = var894 | var1002;
assign var1004 = var898 & var829;
assign var1005 = var897 | var1004;
assign var1006 = var901 & var831;
assign var1007 = var900 | var1006;
assign var1008 = var904 & var833;
assign var1009 = var903 | var1008;
assign var1010 = var907 & var835;
assign var1011 = var906 | var1010;
assign var1012 = var910 & var669;
assign var1013 = var909 | var1012;
assign var1014 = var913 & var671;
assign var1015 = var912 | var1014;
assign var1016 = var916 & var673;
assign var1017 = var915 | var1016;
assign var1018 = var919 & var675;
assign var1019 = var918 | var1018;
assign var1020 = var922 & var497;
assign var1021 = var921 | var1020;
assign var1022 = var925 & var499;
assign var1023 = var924 | var1022;
assign var1024 = var928 & var315;
assign var1025 = var927 | var1024;
assign var1026 = var931 & var0;
assign var1027 = var930 | var1026;
assign var1028 = var65 ^ var0;
assign var1029 = var66 ^ var315;
assign var1030 = var67 ^ var499;
assign var1031 = var68 ^ var497;
assign var1032 = var69 ^ var675;
assign var1033 = var70 ^ var673;
assign var1034 = var71 ^ var671;
assign var1035 = var72 ^ var669;
assign var1036 = var73 ^ var835;
assign var1037 = var74 ^ var833;
assign var1038 = var75 ^ var831;
assign var1039 = var76 ^ var829;
assign var1040 = var77 ^ var827;
assign var1041 = var78 ^ var825;
assign var1042 = var79 ^ var823;
assign var1043 = var80 ^ var821;
assign var1044 = var81 ^ var963;
assign var1045 = var82 ^ var961;
assign var1046 = var83 ^ var959;
assign var1047 = var84 ^ var957;
assign var1048 = var85 ^ var955;
assign var1049 = var86 ^ var953;
assign var1050 = var87 ^ var951;
assign var1051 = var88 ^ var949;
assign var1052 = var89 ^ var947;
assign var1053 = var90 ^ var945;
assign var1054 = var91 ^ var943;
assign var1055 = var92 ^ var941;
assign var1056 = var93 ^ var939;
assign var1057 = var94 ^ var937;
assign var1058 = var95 ^ var935;
assign var1059 = var96 ^ var933;
assign var1060 = var97 ^ var1027;
assign var1061 = var98 ^ var1025;
assign var1062 = var99 ^ var1023;
assign var1063 = var100 ^ var1021;
assign var1064 = var101 ^ var1019;
assign var1065 = var102 ^ var1017;
assign var1066 = var103 ^ var1015;
assign var1067 = var104 ^ var1013;
assign var1068 = var105 ^ var1011;
assign var1069 = var106 ^ var1009;
assign var1070 = var107 ^ var1007;
assign var1071 = var108 ^ var1005;
assign var1072 = var109 ^ var1003;
assign var1073 = var110 ^ var1001;
assign var1074 = var111 ^ var999;
assign var1075 = var112 ^ var997;
assign var1076 = var113 ^ var995;
assign var1077 = var114 ^ var993;
assign var1078 = var115 ^ var991;
assign var1079 = var116 ^ var989;
assign var1080 = var117 ^ var987;
assign var1081 = var118 ^ var985;
assign var1082 = var119 ^ var983;
assign var1083 = var120 ^ var981;
assign var1084 = var121 ^ var979;
assign var1085 = var122 ^ var977;
assign var1086 = var123 ^ var975;
assign var1087 = var124 ^ var973;
assign var1088 = var125 ^ var971;
assign var1089 = var126 ^ var969;
assign var1090 = var127 ^ var967;
assign out0 = var965;
assign out1 = var1090;
assign out2 = var1089;
assign out3 = var1088;
assign out4 = var1087;
assign out5 = var1086;
assign out6 = var1085;
assign out7 = var1084;
assign out8 = var1083;
assign out9 = var1082;
assign out10 = var1081;
assign out11 = var1080;
assign out12 = var1079;
assign out13 = var1078;
assign out14 = var1077;
assign out15 = var1076;
assign out16 = var1075;
assign out17 = var1074;
assign out18 = var1073;
assign out19 = var1072;
assign out20 = var1071;
assign out21 = var1070;
assign out22 = var1069;
assign out23 = var1068;
assign out24 = var1067;
assign out25 = var1066;
assign out26 = var1065;
assign out27 = var1064;
assign out28 = var1063;
assign out29 = var1062;
assign out30 = var1061;
assign out31 = var1060;
assign out32 = var1059;
assign out33 = var1058;
assign out34 = var1057;
assign out35 = var1056;
assign out36 = var1055;
assign out37 = var1054;
assign out38 = var1053;
assign out39 = var1052;
assign out40 = var1051;
assign out41 = var1050;
assign out42 = var1049;
assign out43 = var1048;
assign out44 = var1047;
assign out45 = var1046;
assign out46 = var1045;
assign out47 = var1044;
assign out48 = var1043;
assign out49 = var1042;
assign out50 = var1041;
assign out51 = var1040;
assign out52 = var1039;
assign out53 = var1038;
assign out54 = var1037;
assign out55 = var1036;
assign out56 = var1035;
assign out57 = var1034;
assign out58 = var1033;
assign out59 = var1032;
assign out60 = var1031;
assign out61 = var1030;
assign out62 = var1029;
assign out63 = var1028;
assign out64 = var64;
endmodule 
