module sk64 (in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, in100, in101, in102, in103, in104, in105, in106, in107, in108, in109, in110, in111, in112, in113, in114, in115, in116, in117, in118, in119, in120, in121, in122, in123, in124, in125, in126, in127, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, out30, out31, out32, out33, out34, out35, out36, out37, out38, out39, out40, out41, out42, out43, out44, out45, out46, out47, out48, out49, out50, out51, out52, out53, out54, out55, out56, out57, out58, out59, out60, out61, out62, out63, out64, );
input in0;
input in1;
input in2;
input in3;
input in4;
input in5;
input in6;
input in7;
input in8;
input in9;
input in10;
input in11;
input in12;
input in13;
input in14;
input in15;
input in16;
input in17;
input in18;
input in19;
input in20;
input in21;
input in22;
input in23;
input in24;
input in25;
input in26;
input in27;
input in28;
input in29;
input in30;
input in31;
input in32;
input in33;
input in34;
input in35;
input in36;
input in37;
input in38;
input in39;
input in40;
input in41;
input in42;
input in43;
input in44;
input in45;
input in46;
input in47;
input in48;
input in49;
input in50;
input in51;
input in52;
input in53;
input in54;
input in55;
input in56;
input in57;
input in58;
input in59;
input in60;
input in61;
input in62;
input in63;
input in64;
input in65;
input in66;
input in67;
input in68;
input in69;
input in70;
input in71;
input in72;
input in73;
input in74;
input in75;
input in76;
input in77;
input in78;
input in79;
input in80;
input in81;
input in82;
input in83;
input in84;
input in85;
input in86;
input in87;
input in88;
input in89;
input in90;
input in91;
input in92;
input in93;
input in94;
input in95;
input in96;
input in97;
input in98;
input in99;
input in100;
input in101;
input in102;
input in103;
input in104;
input in105;
input in106;
input in107;
input in108;
input in109;
input in110;
input in111;
input in112;
input in113;
input in114;
input in115;
input in116;
input in117;
input in118;
input in119;
input in120;
input in121;
input in122;
input in123;
input in124;
input in125;
input in126;
input in127;
output out0;
output out1;
output out2;
output out3;
output out4;
output out5;
output out6;
output out7;
output out8;
output out9;
output out10;
output out11;
output out12;
output out13;
output out14;
output out15;
output out16;
output out17;
output out18;
output out19;
output out20;
output out21;
output out22;
output out23;
output out24;
output out25;
output out26;
output out27;
output out28;
output out29;
output out30;
output out31;
output out32;
output out33;
output out34;
output out35;
output out36;
output out37;
output out38;
output out39;
output out40;
output out41;
output out42;
output out43;
output out44;
output out45;
output out46;
output out47;
output out48;
output out49;
output out50;
output out51;
output out52;
output out53;
output out54;
output out55;
output out56;
output out57;
output out58;
output out59;
output out60;
output out61;
output out62;
output out63;
output out64;
wire var0;
wire var1;
wire var2;
wire var3;
wire var4;
wire var5;
wire var6;
wire var7;
wire var8;
wire var9;
wire var10;
wire var11;
wire var12;
wire var13;
wire var14;
wire var15;
wire var16;
wire var17;
wire var18;
wire var19;
wire var20;
wire var21;
wire var22;
wire var23;
wire var24;
wire var25;
wire var26;
wire var27;
wire var28;
wire var29;
wire var30;
wire var31;
wire var32;
wire var33;
wire var34;
wire var35;
wire var36;
wire var37;
wire var38;
wire var39;
wire var40;
wire var41;
wire var42;
wire var43;
wire var44;
wire var45;
wire var46;
wire var47;
wire var48;
wire var49;
wire var50;
wire var51;
wire var52;
wire var53;
wire var54;
wire var55;
wire var56;
wire var57;
wire var58;
wire var59;
wire var60;
wire var61;
wire var62;
wire var63;
wire var64;
wire var65;
wire var66;
wire var67;
wire var68;
wire var69;
wire var70;
wire var71;
wire var72;
wire var73;
wire var74;
wire var75;
wire var76;
wire var77;
wire var78;
wire var79;
wire var80;
wire var81;
wire var82;
wire var83;
wire var84;
wire var85;
wire var86;
wire var87;
wire var88;
wire var89;
wire var90;
wire var91;
wire var92;
wire var93;
wire var94;
wire var95;
wire var96;
wire var97;
wire var98;
wire var99;
wire var100;
wire var101;
wire var102;
wire var103;
wire var104;
wire var105;
wire var106;
wire var107;
wire var108;
wire var109;
wire var110;
wire var111;
wire var112;
wire var113;
wire var114;
wire var115;
wire var116;
wire var117;
wire var118;
wire var119;
wire var120;
wire var121;
wire var122;
wire var123;
wire var124;
wire var125;
wire var126;
wire var127;
wire var128;
wire var129;
wire var130;
wire var131;
wire var132;
wire var133;
wire var134;
wire var135;
wire var136;
wire var137;
wire var138;
wire var139;
wire var140;
wire var141;
wire var142;
wire var143;
wire var144;
wire var145;
wire var146;
wire var147;
wire var148;
wire var149;
wire var150;
wire var151;
wire var152;
wire var153;
wire var154;
wire var155;
wire var156;
wire var157;
wire var158;
wire var159;
wire var160;
wire var161;
wire var162;
wire var163;
wire var164;
wire var165;
wire var166;
wire var167;
wire var168;
wire var169;
wire var170;
wire var171;
wire var172;
wire var173;
wire var174;
wire var175;
wire var176;
wire var177;
wire var178;
wire var179;
wire var180;
wire var181;
wire var182;
wire var183;
wire var184;
wire var185;
wire var186;
wire var187;
wire var188;
wire var189;
wire var190;
wire var191;
wire var192;
wire var193;
wire var194;
wire var195;
wire var196;
wire var197;
wire var198;
wire var199;
wire var200;
wire var201;
wire var202;
wire var203;
wire var204;
wire var205;
wire var206;
wire var207;
wire var208;
wire var209;
wire var210;
wire var211;
wire var212;
wire var213;
wire var214;
wire var215;
wire var216;
wire var217;
wire var218;
wire var219;
wire var220;
wire var221;
wire var222;
wire var223;
wire var224;
wire var225;
wire var226;
wire var227;
wire var228;
wire var229;
wire var230;
wire var231;
wire var232;
wire var233;
wire var234;
wire var235;
wire var236;
wire var237;
wire var238;
wire var239;
wire var240;
wire var241;
wire var242;
wire var243;
wire var244;
wire var245;
wire var246;
wire var247;
wire var248;
wire var249;
wire var250;
wire var251;
wire var252;
wire var253;
wire var254;
wire var255;
wire var256;
wire var257;
wire var258;
wire var259;
wire var260;
wire var261;
wire var262;
wire var263;
wire var264;
wire var265;
wire var266;
wire var267;
wire var268;
wire var269;
wire var270;
wire var271;
wire var272;
wire var273;
wire var274;
wire var275;
wire var276;
wire var277;
wire var278;
wire var279;
wire var280;
wire var281;
wire var282;
wire var283;
wire var284;
wire var285;
wire var286;
wire var287;
wire var288;
wire var289;
wire var290;
wire var291;
wire var292;
wire var293;
wire var294;
wire var295;
wire var296;
wire var297;
wire var298;
wire var299;
wire var300;
wire var301;
wire var302;
wire var303;
wire var304;
wire var305;
wire var306;
wire var307;
wire var308;
wire var309;
wire var310;
wire var311;
wire var312;
wire var313;
wire var314;
wire var315;
wire var316;
wire var317;
wire var318;
wire var319;
wire var320;
wire var321;
wire var322;
wire var323;
wire var324;
wire var325;
wire var326;
wire var327;
wire var328;
wire var329;
wire var330;
wire var331;
wire var332;
wire var333;
wire var334;
wire var335;
wire var336;
wire var337;
wire var338;
wire var339;
wire var340;
wire var341;
wire var342;
wire var343;
wire var344;
wire var345;
wire var346;
wire var347;
wire var348;
wire var349;
wire var350;
wire var351;
wire var352;
wire var353;
wire var354;
wire var355;
wire var356;
wire var357;
wire var358;
wire var359;
wire var360;
wire var361;
wire var362;
wire var363;
wire var364;
wire var365;
wire var366;
wire var367;
wire var368;
wire var369;
wire var370;
wire var371;
wire var372;
wire var373;
wire var374;
wire var375;
wire var376;
wire var377;
wire var378;
wire var379;
wire var380;
wire var381;
wire var382;
wire var383;
wire var384;
wire var385;
wire var386;
wire var387;
wire var388;
wire var389;
wire var390;
wire var391;
wire var392;
wire var393;
wire var394;
wire var395;
wire var396;
wire var397;
wire var398;
wire var399;
wire var400;
wire var401;
wire var402;
wire var403;
wire var404;
wire var405;
wire var406;
wire var407;
wire var408;
wire var409;
wire var410;
wire var411;
wire var412;
wire var413;
wire var414;
wire var415;
wire var416;
wire var417;
wire var418;
wire var419;
wire var420;
wire var421;
wire var422;
wire var423;
wire var424;
wire var425;
wire var426;
wire var427;
wire var428;
wire var429;
wire var430;
wire var431;
wire var432;
wire var433;
wire var434;
wire var435;
wire var436;
wire var437;
wire var438;
wire var439;
wire var440;
wire var441;
wire var442;
wire var443;
wire var444;
wire var445;
wire var446;
wire var447;
wire var448;
wire var449;
wire var450;
wire var451;
wire var452;
wire var453;
wire var454;
wire var455;
wire var456;
wire var457;
wire var458;
wire var459;
wire var460;
wire var461;
wire var462;
wire var463;
wire var464;
wire var465;
wire var466;
wire var467;
wire var468;
wire var469;
wire var470;
wire var471;
wire var472;
wire var473;
wire var474;
wire var475;
wire var476;
wire var477;
wire var478;
wire var479;
wire var480;
wire var481;
wire var482;
wire var483;
wire var484;
wire var485;
wire var486;
wire var487;
wire var488;
wire var489;
wire var490;
wire var491;
wire var492;
wire var493;
wire var494;
wire var495;
wire var496;
wire var497;
wire var498;
wire var499;
wire var500;
wire var501;
wire var502;
wire var503;
wire var504;
wire var505;
wire var506;
wire var507;
wire var508;
wire var509;
wire var510;
wire var511;
wire var512;
wire var513;
wire var514;
wire var515;
wire var516;
wire var517;
wire var518;
wire var519;
wire var520;
wire var521;
wire var522;
wire var523;
wire var524;
wire var525;
wire var526;
wire var527;
wire var528;
wire var529;
wire var530;
wire var531;
wire var532;
wire var533;
wire var534;
wire var535;
wire var536;
wire var537;
wire var538;
wire var539;
wire var540;
wire var541;
wire var542;
wire var543;
wire var544;
wire var545;
wire var546;
wire var547;
wire var548;
wire var549;
wire var550;
wire var551;
wire var552;
wire var553;
wire var554;
wire var555;
wire var556;
wire var557;
wire var558;
wire var559;
wire var560;
wire var561;
wire var562;
wire var563;
wire var564;
wire var565;
wire var566;
wire var567;
wire var568;
wire var569;
wire var570;
wire var571;
wire var572;
wire var573;
wire var574;
wire var575;
wire var576;
wire var577;
wire var578;
wire var579;
wire var580;
wire var581;
wire var582;
wire var583;
wire var584;
wire var585;
wire var586;
wire var587;
wire var588;
wire var589;
wire var590;
wire var591;
wire var592;
wire var593;
wire var594;
wire var595;
wire var596;
wire var597;
wire var598;
wire var599;
wire var600;
wire var601;
wire var602;
wire var603;
wire var604;
wire var605;
wire var606;
wire var607;
wire var608;
wire var609;
wire var610;
wire var611;
wire var612;
wire var613;
wire var614;
wire var615;
wire var616;
wire var617;
wire var618;
wire var619;
wire var620;
wire var621;
wire var622;
wire var623;
wire var624;
wire var625;
wire var626;
wire var627;
wire var628;
wire var629;
wire var630;
wire var631;
wire var632;
wire var633;
wire var634;
wire var635;
wire var636;
wire var637;
wire var638;
wire var639;
wire var640;
wire var641;
wire var642;
wire var643;
wire var644;
wire var645;
wire var646;
wire var647;
wire var648;
wire var649;
wire var650;
wire var651;
wire var652;
wire var653;
wire var654;
wire var655;
wire var656;
wire var657;
wire var658;
wire var659;
wire var660;
wire var661;
wire var662;
wire var663;
wire var664;
wire var665;
wire var666;
wire var667;
wire var668;
wire var669;
wire var670;
wire var671;
wire var672;
wire var673;
wire var674;
wire var675;
wire var676;
wire var677;
wire var678;
wire var679;
wire var680;
wire var681;
wire var682;
wire var683;
wire var684;
wire var685;
wire var686;
wire var687;
wire var688;
wire var689;
wire var690;
wire var691;
wire var692;
wire var693;
wire var694;
wire var695;
wire var696;
wire var697;
wire var698;
wire var699;
wire var700;
wire var701;
wire var702;
wire var703;
assign var0 = in127 & in63;
assign var1 = in126 & in62;
assign var2 = in125 & in61;
assign var3 = in124 & in60;
assign var4 = in123 & in59;
assign var5 = in122 & in58;
assign var6 = in121 & in57;
assign var7 = in120 & in56;
assign var8 = in119 & in55;
assign var9 = in118 & in54;
assign var10 = in117 & in53;
assign var11 = in116 & in52;
assign var12 = in115 & in51;
assign var13 = in114 & in50;
assign var14 = in113 & in49;
assign var15 = in112 & in48;
assign var16 = in111 & in47;
assign var17 = in110 & in46;
assign var18 = in109 & in45;
assign var19 = in108 & in44;
assign var20 = in107 & in43;
assign var21 = in106 & in42;
assign var22 = in105 & in41;
assign var23 = in104 & in40;
assign var24 = in103 & in39;
assign var25 = in102 & in38;
assign var26 = in101 & in37;
assign var27 = in100 & in36;
assign var28 = in99 & in35;
assign var29 = in98 & in34;
assign var30 = in97 & in33;
assign var31 = in96 & in32;
assign var32 = in95 & in31;
assign var33 = in94 & in30;
assign var34 = in93 & in29;
assign var35 = in92 & in28;
assign var36 = in91 & in27;
assign var37 = in90 & in26;
assign var38 = in89 & in25;
assign var39 = in88 & in24;
assign var40 = in87 & in23;
assign var41 = in86 & in22;
assign var42 = in85 & in21;
assign var43 = in84 & in20;
assign var44 = in83 & in19;
assign var45 = in82 & in18;
assign var46 = in81 & in17;
assign var47 = in80 & in16;
assign var48 = in79 & in15;
assign var49 = in78 & in14;
assign var50 = in77 & in13;
assign var51 = in76 & in12;
assign var52 = in75 & in11;
assign var53 = in74 & in10;
assign var54 = in73 & in9;
assign var55 = in72 & in8;
assign var56 = in71 & in7;
assign var57 = in70 & in6;
assign var58 = in69 & in5;
assign var59 = in68 & in4;
assign var60 = in67 & in3;
assign var61 = in66 & in2;
assign var62 = in65 & in1;
assign var63 = in64 & in0;
assign var64 = in127 ^ in63;
assign var65 = in126 ^ in62;
assign var66 = in125 ^ in61;
assign var67 = in124 ^ in60;
assign var68 = in123 ^ in59;
assign var69 = in122 ^ in58;
assign var70 = in121 ^ in57;
assign var71 = in120 ^ in56;
assign var72 = in119 ^ in55;
assign var73 = in118 ^ in54;
assign var74 = in117 ^ in53;
assign var75 = in116 ^ in52;
assign var76 = in115 ^ in51;
assign var77 = in114 ^ in50;
assign var78 = in113 ^ in49;
assign var79 = in112 ^ in48;
assign var80 = in111 ^ in47;
assign var81 = in110 ^ in46;
assign var82 = in109 ^ in45;
assign var83 = in108 ^ in44;
assign var84 = in107 ^ in43;
assign var85 = in106 ^ in42;
assign var86 = in105 ^ in41;
assign var87 = in104 ^ in40;
assign var88 = in103 ^ in39;
assign var89 = in102 ^ in38;
assign var90 = in101 ^ in37;
assign var91 = in100 ^ in36;
assign var92 = in99 ^ in35;
assign var93 = in98 ^ in34;
assign var94 = in97 ^ in33;
assign var95 = in96 ^ in32;
assign var96 = in95 ^ in31;
assign var97 = in94 ^ in30;
assign var98 = in93 ^ in29;
assign var99 = in92 ^ in28;
assign var100 = in91 ^ in27;
assign var101 = in90 ^ in26;
assign var102 = in89 ^ in25;
assign var103 = in88 ^ in24;
assign var104 = in87 ^ in23;
assign var105 = in86 ^ in22;
assign var106 = in85 ^ in21;
assign var107 = in84 ^ in20;
assign var108 = in83 ^ in19;
assign var109 = in82 ^ in18;
assign var110 = in81 ^ in17;
assign var111 = in80 ^ in16;
assign var112 = in79 ^ in15;
assign var113 = in78 ^ in14;
assign var114 = in77 ^ in13;
assign var115 = in76 ^ in12;
assign var116 = in75 ^ in11;
assign var117 = in74 ^ in10;
assign var118 = in73 ^ in9;
assign var119 = in72 ^ in8;
assign var120 = in71 ^ in7;
assign var121 = in70 ^ in6;
assign var122 = in69 ^ in5;
assign var123 = in68 ^ in4;
assign var124 = in67 ^ in3;
assign var125 = in66 ^ in2;
assign var126 = in65 ^ in1;
assign var127 = in64 ^ in0;
assign var128 = var127 & var62;
assign var129 = var63 | var128;
assign var130 = var127 & var126;
assign var131 = var125 & var60;
assign var132 = var61 | var131;
assign var133 = var125 & var124;
assign var134 = var123 & var58;
assign var135 = var59 | var134;
assign var136 = var123 & var122;
assign var137 = var121 & var56;
assign var138 = var57 | var137;
assign var139 = var121 & var120;
assign var140 = var119 & var54;
assign var141 = var55 | var140;
assign var142 = var119 & var118;
assign var143 = var117 & var52;
assign var144 = var53 | var143;
assign var145 = var117 & var116;
assign var146 = var115 & var50;
assign var147 = var51 | var146;
assign var148 = var115 & var114;
assign var149 = var113 & var48;
assign var150 = var49 | var149;
assign var151 = var113 & var112;
assign var152 = var111 & var46;
assign var153 = var47 | var152;
assign var154 = var111 & var110;
assign var155 = var109 & var44;
assign var156 = var45 | var155;
assign var157 = var109 & var108;
assign var158 = var107 & var42;
assign var159 = var43 | var158;
assign var160 = var107 & var106;
assign var161 = var105 & var40;
assign var162 = var41 | var161;
assign var163 = var105 & var104;
assign var164 = var103 & var38;
assign var165 = var39 | var164;
assign var166 = var103 & var102;
assign var167 = var101 & var36;
assign var168 = var37 | var167;
assign var169 = var101 & var100;
assign var170 = var99 & var34;
assign var171 = var35 | var170;
assign var172 = var99 & var98;
assign var173 = var97 & var32;
assign var174 = var33 | var173;
assign var175 = var97 & var96;
assign var176 = var95 & var30;
assign var177 = var31 | var176;
assign var178 = var95 & var94;
assign var179 = var93 & var28;
assign var180 = var29 | var179;
assign var181 = var93 & var92;
assign var182 = var91 & var26;
assign var183 = var27 | var182;
assign var184 = var91 & var90;
assign var185 = var89 & var24;
assign var186 = var25 | var185;
assign var187 = var89 & var88;
assign var188 = var87 & var22;
assign var189 = var23 | var188;
assign var190 = var87 & var86;
assign var191 = var85 & var20;
assign var192 = var21 | var191;
assign var193 = var85 & var84;
assign var194 = var83 & var18;
assign var195 = var19 | var194;
assign var196 = var83 & var82;
assign var197 = var81 & var16;
assign var198 = var17 | var197;
assign var199 = var81 & var80;
assign var200 = var79 & var14;
assign var201 = var15 | var200;
assign var202 = var79 & var78;
assign var203 = var77 & var12;
assign var204 = var13 | var203;
assign var205 = var77 & var76;
assign var206 = var75 & var10;
assign var207 = var11 | var206;
assign var208 = var75 & var74;
assign var209 = var73 & var8;
assign var210 = var9 | var209;
assign var211 = var73 & var72;
assign var212 = var71 & var6;
assign var213 = var7 | var212;
assign var214 = var71 & var70;
assign var215 = var69 & var4;
assign var216 = var5 | var215;
assign var217 = var69 & var68;
assign var218 = var67 & var2;
assign var219 = var3 | var218;
assign var220 = var67 & var66;
assign var221 = var65 & var0;
assign var222 = var1 | var221;
assign var223 = var130 & var132;
assign var224 = var129 | var223;
assign var225 = var130 & var133;
assign var226 = var126 & var132;
assign var227 = var62 | var226;
assign var228 = var126 & var133;
assign var229 = var136 & var138;
assign var230 = var135 | var229;
assign var231 = var136 & var139;
assign var232 = var122 & var138;
assign var233 = var58 | var232;
assign var234 = var122 & var139;
assign var235 = var142 & var144;
assign var236 = var141 | var235;
assign var237 = var142 & var145;
assign var238 = var118 & var144;
assign var239 = var54 | var238;
assign var240 = var118 & var145;
assign var241 = var148 & var150;
assign var242 = var147 | var241;
assign var243 = var148 & var151;
assign var244 = var114 & var150;
assign var245 = var50 | var244;
assign var246 = var114 & var151;
assign var247 = var154 & var156;
assign var248 = var153 | var247;
assign var249 = var154 & var157;
assign var250 = var110 & var156;
assign var251 = var46 | var250;
assign var252 = var110 & var157;
assign var253 = var160 & var162;
assign var254 = var159 | var253;
assign var255 = var160 & var163;
assign var256 = var106 & var162;
assign var257 = var42 | var256;
assign var258 = var106 & var163;
assign var259 = var166 & var168;
assign var260 = var165 | var259;
assign var261 = var166 & var169;
assign var262 = var102 & var168;
assign var263 = var38 | var262;
assign var264 = var102 & var169;
assign var265 = var172 & var174;
assign var266 = var171 | var265;
assign var267 = var172 & var175;
assign var268 = var98 & var174;
assign var269 = var34 | var268;
assign var270 = var98 & var175;
assign var271 = var178 & var180;
assign var272 = var177 | var271;
assign var273 = var178 & var181;
assign var274 = var94 & var180;
assign var275 = var30 | var274;
assign var276 = var94 & var181;
assign var277 = var184 & var186;
assign var278 = var183 | var277;
assign var279 = var184 & var187;
assign var280 = var90 & var186;
assign var281 = var26 | var280;
assign var282 = var90 & var187;
assign var283 = var190 & var192;
assign var284 = var189 | var283;
assign var285 = var190 & var193;
assign var286 = var86 & var192;
assign var287 = var22 | var286;
assign var288 = var86 & var193;
assign var289 = var196 & var198;
assign var290 = var195 | var289;
assign var291 = var196 & var199;
assign var292 = var82 & var198;
assign var293 = var18 | var292;
assign var294 = var82 & var199;
assign var295 = var202 & var204;
assign var296 = var201 | var295;
assign var297 = var202 & var205;
assign var298 = var78 & var204;
assign var299 = var14 | var298;
assign var300 = var78 & var205;
assign var301 = var208 & var210;
assign var302 = var207 | var301;
assign var303 = var208 & var211;
assign var304 = var74 & var210;
assign var305 = var10 | var304;
assign var306 = var74 & var211;
assign var307 = var214 & var216;
assign var308 = var213 | var307;
assign var309 = var214 & var217;
assign var310 = var70 & var216;
assign var311 = var6 | var310;
assign var312 = var70 & var217;
assign var313 = var220 & var222;
assign var314 = var219 | var313;
assign var315 = var66 & var222;
assign var316 = var2 | var315;
assign var317 = var225 & var230;
assign var318 = var224 | var317;
assign var319 = var225 & var231;
assign var320 = var228 & var230;
assign var321 = var227 | var320;
assign var322 = var228 & var231;
assign var323 = var133 & var230;
assign var324 = var132 | var323;
assign var325 = var133 & var231;
assign var326 = var124 & var230;
assign var327 = var60 | var326;
assign var328 = var124 & var231;
assign var329 = var237 & var242;
assign var330 = var236 | var329;
assign var331 = var237 & var243;
assign var332 = var240 & var242;
assign var333 = var239 | var332;
assign var334 = var240 & var243;
assign var335 = var145 & var242;
assign var336 = var144 | var335;
assign var337 = var145 & var243;
assign var338 = var116 & var242;
assign var339 = var52 | var338;
assign var340 = var116 & var243;
assign var341 = var249 & var254;
assign var342 = var248 | var341;
assign var343 = var249 & var255;
assign var344 = var252 & var254;
assign var345 = var251 | var344;
assign var346 = var252 & var255;
assign var347 = var157 & var254;
assign var348 = var156 | var347;
assign var349 = var157 & var255;
assign var350 = var108 & var254;
assign var351 = var44 | var350;
assign var352 = var108 & var255;
assign var353 = var261 & var266;
assign var354 = var260 | var353;
assign var355 = var261 & var267;
assign var356 = var264 & var266;
assign var357 = var263 | var356;
assign var358 = var264 & var267;
assign var359 = var169 & var266;
assign var360 = var168 | var359;
assign var361 = var169 & var267;
assign var362 = var100 & var266;
assign var363 = var36 | var362;
assign var364 = var100 & var267;
assign var365 = var273 & var278;
assign var366 = var272 | var365;
assign var367 = var273 & var279;
assign var368 = var276 & var278;
assign var369 = var275 | var368;
assign var370 = var276 & var279;
assign var371 = var181 & var278;
assign var372 = var180 | var371;
assign var373 = var181 & var279;
assign var374 = var92 & var278;
assign var375 = var28 | var374;
assign var376 = var92 & var279;
assign var377 = var285 & var290;
assign var378 = var284 | var377;
assign var379 = var285 & var291;
assign var380 = var288 & var290;
assign var381 = var287 | var380;
assign var382 = var288 & var291;
assign var383 = var193 & var290;
assign var384 = var192 | var383;
assign var385 = var193 & var291;
assign var386 = var84 & var290;
assign var387 = var20 | var386;
assign var388 = var84 & var291;
assign var389 = var297 & var302;
assign var390 = var296 | var389;
assign var391 = var297 & var303;
assign var392 = var300 & var302;
assign var393 = var299 | var392;
assign var394 = var300 & var303;
assign var395 = var205 & var302;
assign var396 = var204 | var395;
assign var397 = var205 & var303;
assign var398 = var76 & var302;
assign var399 = var12 | var398;
assign var400 = var76 & var303;
assign var401 = var309 & var314;
assign var402 = var308 | var401;
assign var403 = var312 & var314;
assign var404 = var311 | var403;
assign var405 = var217 & var314;
assign var406 = var216 | var405;
assign var407 = var68 & var314;
assign var408 = var4 | var407;
assign var409 = var319 & var330;
assign var410 = var318 | var409;
assign var411 = var319 & var331;
assign var412 = var322 & var330;
assign var413 = var321 | var412;
assign var414 = var322 & var331;
assign var415 = var325 & var330;
assign var416 = var324 | var415;
assign var417 = var325 & var331;
assign var418 = var328 & var330;
assign var419 = var327 | var418;
assign var420 = var328 & var331;
assign var421 = var231 & var330;
assign var422 = var230 | var421;
assign var423 = var231 & var331;
assign var424 = var234 & var330;
assign var425 = var233 | var424;
assign var426 = var234 & var331;
assign var427 = var139 & var330;
assign var428 = var138 | var427;
assign var429 = var139 & var331;
assign var430 = var120 & var330;
assign var431 = var56 | var430;
assign var432 = var120 & var331;
assign var433 = var343 & var354;
assign var434 = var342 | var433;
assign var435 = var343 & var355;
assign var436 = var346 & var354;
assign var437 = var345 | var436;
assign var438 = var346 & var355;
assign var439 = var349 & var354;
assign var440 = var348 | var439;
assign var441 = var349 & var355;
assign var442 = var352 & var354;
assign var443 = var351 | var442;
assign var444 = var352 & var355;
assign var445 = var255 & var354;
assign var446 = var254 | var445;
assign var447 = var255 & var355;
assign var448 = var258 & var354;
assign var449 = var257 | var448;
assign var450 = var258 & var355;
assign var451 = var163 & var354;
assign var452 = var162 | var451;
assign var453 = var163 & var355;
assign var454 = var104 & var354;
assign var455 = var40 | var454;
assign var456 = var104 & var355;
assign var457 = var367 & var378;
assign var458 = var366 | var457;
assign var459 = var367 & var379;
assign var460 = var370 & var378;
assign var461 = var369 | var460;
assign var462 = var370 & var379;
assign var463 = var373 & var378;
assign var464 = var372 | var463;
assign var465 = var373 & var379;
assign var466 = var376 & var378;
assign var467 = var375 | var466;
assign var468 = var376 & var379;
assign var469 = var279 & var378;
assign var470 = var278 | var469;
assign var471 = var279 & var379;
assign var472 = var282 & var378;
assign var473 = var281 | var472;
assign var474 = var282 & var379;
assign var475 = var187 & var378;
assign var476 = var186 | var475;
assign var477 = var187 & var379;
assign var478 = var88 & var378;
assign var479 = var24 | var478;
assign var480 = var88 & var379;
assign var481 = var391 & var402;
assign var482 = var390 | var481;
assign var483 = var394 & var402;
assign var484 = var393 | var483;
assign var485 = var397 & var402;
assign var486 = var396 | var485;
assign var487 = var400 & var402;
assign var488 = var399 | var487;
assign var489 = var303 & var402;
assign var490 = var302 | var489;
assign var491 = var306 & var402;
assign var492 = var305 | var491;
assign var493 = var211 & var402;
assign var494 = var210 | var493;
assign var495 = var72 & var402;
assign var496 = var8 | var495;
assign var497 = var411 & var434;
assign var498 = var410 | var497;
assign var499 = var411 & var435;
assign var500 = var414 & var434;
assign var501 = var413 | var500;
assign var502 = var414 & var435;
assign var503 = var417 & var434;
assign var504 = var416 | var503;
assign var505 = var417 & var435;
assign var506 = var420 & var434;
assign var507 = var419 | var506;
assign var508 = var420 & var435;
assign var509 = var423 & var434;
assign var510 = var422 | var509;
assign var511 = var423 & var435;
assign var512 = var426 & var434;
assign var513 = var425 | var512;
assign var514 = var426 & var435;
assign var515 = var429 & var434;
assign var516 = var428 | var515;
assign var517 = var429 & var435;
assign var518 = var432 & var434;
assign var519 = var431 | var518;
assign var520 = var432 & var435;
assign var521 = var331 & var434;
assign var522 = var330 | var521;
assign var523 = var331 & var435;
assign var524 = var334 & var434;
assign var525 = var333 | var524;
assign var526 = var334 & var435;
assign var527 = var337 & var434;
assign var528 = var336 | var527;
assign var529 = var337 & var435;
assign var530 = var340 & var434;
assign var531 = var339 | var530;
assign var532 = var340 & var435;
assign var533 = var243 & var434;
assign var534 = var242 | var533;
assign var535 = var243 & var435;
assign var536 = var246 & var434;
assign var537 = var245 | var536;
assign var538 = var246 & var435;
assign var539 = var151 & var434;
assign var540 = var150 | var539;
assign var541 = var151 & var435;
assign var542 = var112 & var434;
assign var543 = var48 | var542;
assign var544 = var112 & var435;
assign var545 = var459 & var482;
assign var546 = var458 | var545;
assign var547 = var462 & var482;
assign var548 = var461 | var547;
assign var549 = var465 & var482;
assign var550 = var464 | var549;
assign var551 = var468 & var482;
assign var552 = var467 | var551;
assign var553 = var471 & var482;
assign var554 = var470 | var553;
assign var555 = var474 & var482;
assign var556 = var473 | var555;
assign var557 = var477 & var482;
assign var558 = var476 | var557;
assign var559 = var480 & var482;
assign var560 = var479 | var559;
assign var561 = var379 & var482;
assign var562 = var378 | var561;
assign var563 = var382 & var482;
assign var564 = var381 | var563;
assign var565 = var385 & var482;
assign var566 = var384 | var565;
assign var567 = var388 & var482;
assign var568 = var387 | var567;
assign var569 = var291 & var482;
assign var570 = var290 | var569;
assign var571 = var294 & var482;
assign var572 = var293 | var571;
assign var573 = var199 & var482;
assign var574 = var198 | var573;
assign var575 = var80 & var482;
assign var576 = var16 | var575;
assign var577 = var499 & var546;
assign var578 = var498 | var577;
assign var579 = var502 & var546;
assign var580 = var501 | var579;
assign var581 = var505 & var546;
assign var582 = var504 | var581;
assign var583 = var508 & var546;
assign var584 = var507 | var583;
assign var585 = var511 & var546;
assign var586 = var510 | var585;
assign var587 = var514 & var546;
assign var588 = var513 | var587;
assign var589 = var517 & var546;
assign var590 = var516 | var589;
assign var591 = var520 & var546;
assign var592 = var519 | var591;
assign var593 = var523 & var546;
assign var594 = var522 | var593;
assign var595 = var526 & var546;
assign var596 = var525 | var595;
assign var597 = var529 & var546;
assign var598 = var528 | var597;
assign var599 = var532 & var546;
assign var600 = var531 | var599;
assign var601 = var535 & var546;
assign var602 = var534 | var601;
assign var603 = var538 & var546;
assign var604 = var537 | var603;
assign var605 = var541 & var546;
assign var606 = var540 | var605;
assign var607 = var544 & var546;
assign var608 = var543 | var607;
assign var609 = var435 & var546;
assign var610 = var434 | var609;
assign var611 = var438 & var546;
assign var612 = var437 | var611;
assign var613 = var441 & var546;
assign var614 = var440 | var613;
assign var615 = var444 & var546;
assign var616 = var443 | var615;
assign var617 = var447 & var546;
assign var618 = var446 | var617;
assign var619 = var450 & var546;
assign var620 = var449 | var619;
assign var621 = var453 & var546;
assign var622 = var452 | var621;
assign var623 = var456 & var546;
assign var624 = var455 | var623;
assign var625 = var355 & var546;
assign var626 = var354 | var625;
assign var627 = var358 & var546;
assign var628 = var357 | var627;
assign var629 = var361 & var546;
assign var630 = var360 | var629;
assign var631 = var364 & var546;
assign var632 = var363 | var631;
assign var633 = var267 & var546;
assign var634 = var266 | var633;
assign var635 = var270 & var546;
assign var636 = var269 | var635;
assign var637 = var175 & var546;
assign var638 = var174 | var637;
assign var639 = var96 & var546;
assign var640 = var32 | var639;
assign var641 = var65 ^ var0;
assign var642 = var66 ^ var222;
assign var643 = var67 ^ var316;
assign var644 = var68 ^ var314;
assign var645 = var69 ^ var408;
assign var646 = var70 ^ var406;
assign var647 = var71 ^ var404;
assign var648 = var72 ^ var402;
assign var649 = var73 ^ var496;
assign var650 = var74 ^ var494;
assign var651 = var75 ^ var492;
assign var652 = var76 ^ var490;
assign var653 = var77 ^ var488;
assign var654 = var78 ^ var486;
assign var655 = var79 ^ var484;
assign var656 = var80 ^ var482;
assign var657 = var81 ^ var576;
assign var658 = var82 ^ var574;
assign var659 = var83 ^ var572;
assign var660 = var84 ^ var570;
assign var661 = var85 ^ var568;
assign var662 = var86 ^ var566;
assign var663 = var87 ^ var564;
assign var664 = var88 ^ var562;
assign var665 = var89 ^ var560;
assign var666 = var90 ^ var558;
assign var667 = var91 ^ var556;
assign var668 = var92 ^ var554;
assign var669 = var93 ^ var552;
assign var670 = var94 ^ var550;
assign var671 = var95 ^ var548;
assign var672 = var96 ^ var546;
assign var673 = var97 ^ var640;
assign var674 = var98 ^ var638;
assign var675 = var99 ^ var636;
assign var676 = var100 ^ var634;
assign var677 = var101 ^ var632;
assign var678 = var102 ^ var630;
assign var679 = var103 ^ var628;
assign var680 = var104 ^ var626;
assign var681 = var105 ^ var624;
assign var682 = var106 ^ var622;
assign var683 = var107 ^ var620;
assign var684 = var108 ^ var618;
assign var685 = var109 ^ var616;
assign var686 = var110 ^ var614;
assign var687 = var111 ^ var612;
assign var688 = var112 ^ var610;
assign var689 = var113 ^ var608;
assign var690 = var114 ^ var606;
assign var691 = var115 ^ var604;
assign var692 = var116 ^ var602;
assign var693 = var117 ^ var600;
assign var694 = var118 ^ var598;
assign var695 = var119 ^ var596;
assign var696 = var120 ^ var594;
assign var697 = var121 ^ var592;
assign var698 = var122 ^ var590;
assign var699 = var123 ^ var588;
assign var700 = var124 ^ var586;
assign var701 = var125 ^ var584;
assign var702 = var126 ^ var582;
assign var703 = var127 ^ var580;
assign out0 = var578;
assign out1 = var703;
assign out2 = var702;
assign out3 = var701;
assign out4 = var700;
assign out5 = var699;
assign out6 = var698;
assign out7 = var697;
assign out8 = var696;
assign out9 = var695;
assign out10 = var694;
assign out11 = var693;
assign out12 = var692;
assign out13 = var691;
assign out14 = var690;
assign out15 = var689;
assign out16 = var688;
assign out17 = var687;
assign out18 = var686;
assign out19 = var685;
assign out20 = var684;
assign out21 = var683;
assign out22 = var682;
assign out23 = var681;
assign out24 = var680;
assign out25 = var679;
assign out26 = var678;
assign out27 = var677;
assign out28 = var676;
assign out29 = var675;
assign out30 = var674;
assign out31 = var673;
assign out32 = var672;
assign out33 = var671;
assign out34 = var670;
assign out35 = var669;
assign out36 = var668;
assign out37 = var667;
assign out38 = var666;
assign out39 = var665;
assign out40 = var664;
assign out41 = var663;
assign out42 = var662;
assign out43 = var661;
assign out44 = var660;
assign out45 = var659;
assign out46 = var658;
assign out47 = var657;
assign out48 = var656;
assign out49 = var655;
assign out50 = var654;
assign out51 = var653;
assign out52 = var652;
assign out53 = var651;
assign out54 = var650;
assign out55 = var649;
assign out56 = var648;
assign out57 = var647;
assign out58 = var646;
assign out59 = var645;
assign out60 = var644;
assign out61 = var643;
assign out62 = var642;
assign out63 = var641;
assign out64 = var64;
endmodule 
