module lf128 (in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, in100, in101, in102, in103, in104, in105, in106, in107, in108, in109, in110, in111, in112, in113, in114, in115, in116, in117, in118, in119, in120, in121, in122, in123, in124, in125, in126, in127, in128, in129, in130, in131, in132, in133, in134, in135, in136, in137, in138, in139, in140, in141, in142, in143, in144, in145, in146, in147, in148, in149, in150, in151, in152, in153, in154, in155, in156, in157, in158, in159, in160, in161, in162, in163, in164, in165, in166, in167, in168, in169, in170, in171, in172, in173, in174, in175, in176, in177, in178, in179, in180, in181, in182, in183, in184, in185, in186, in187, in188, in189, in190, in191, in192, in193, in194, in195, in196, in197, in198, in199, in200, in201, in202, in203, in204, in205, in206, in207, in208, in209, in210, in211, in212, in213, in214, in215, in216, in217, in218, in219, in220, in221, in222, in223, in224, in225, in226, in227, in228, in229, in230, in231, in232, in233, in234, in235, in236, in237, in238, in239, in240, in241, in242, in243, in244, in245, in246, in247, in248, in249, in250, in251, in252, in253, in254, in255, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, out30, out31, out32, out33, out34, out35, out36, out37, out38, out39, out40, out41, out42, out43, out44, out45, out46, out47, out48, out49, out50, out51, out52, out53, out54, out55, out56, out57, out58, out59, out60, out61, out62, out63, out64, out65, out66, out67, out68, out69, out70, out71, out72, out73, out74, out75, out76, out77, out78, out79, out80, out81, out82, out83, out84, out85, out86, out87, out88, out89, out90, out91, out92, out93, out94, out95, out96, out97, out98, out99, out100, out101, out102, out103, out104, out105, out106, out107, out108, out109, out110, out111, out112, out113, out114, out115, out116, out117, out118, out119, out120, out121, out122, out123, out124, out125, out126, out127, out128, );
input in0;
input in1;
input in2;
input in3;
input in4;
input in5;
input in6;
input in7;
input in8;
input in9;
input in10;
input in11;
input in12;
input in13;
input in14;
input in15;
input in16;
input in17;
input in18;
input in19;
input in20;
input in21;
input in22;
input in23;
input in24;
input in25;
input in26;
input in27;
input in28;
input in29;
input in30;
input in31;
input in32;
input in33;
input in34;
input in35;
input in36;
input in37;
input in38;
input in39;
input in40;
input in41;
input in42;
input in43;
input in44;
input in45;
input in46;
input in47;
input in48;
input in49;
input in50;
input in51;
input in52;
input in53;
input in54;
input in55;
input in56;
input in57;
input in58;
input in59;
input in60;
input in61;
input in62;
input in63;
input in64;
input in65;
input in66;
input in67;
input in68;
input in69;
input in70;
input in71;
input in72;
input in73;
input in74;
input in75;
input in76;
input in77;
input in78;
input in79;
input in80;
input in81;
input in82;
input in83;
input in84;
input in85;
input in86;
input in87;
input in88;
input in89;
input in90;
input in91;
input in92;
input in93;
input in94;
input in95;
input in96;
input in97;
input in98;
input in99;
input in100;
input in101;
input in102;
input in103;
input in104;
input in105;
input in106;
input in107;
input in108;
input in109;
input in110;
input in111;
input in112;
input in113;
input in114;
input in115;
input in116;
input in117;
input in118;
input in119;
input in120;
input in121;
input in122;
input in123;
input in124;
input in125;
input in126;
input in127;
input in128;
input in129;
input in130;
input in131;
input in132;
input in133;
input in134;
input in135;
input in136;
input in137;
input in138;
input in139;
input in140;
input in141;
input in142;
input in143;
input in144;
input in145;
input in146;
input in147;
input in148;
input in149;
input in150;
input in151;
input in152;
input in153;
input in154;
input in155;
input in156;
input in157;
input in158;
input in159;
input in160;
input in161;
input in162;
input in163;
input in164;
input in165;
input in166;
input in167;
input in168;
input in169;
input in170;
input in171;
input in172;
input in173;
input in174;
input in175;
input in176;
input in177;
input in178;
input in179;
input in180;
input in181;
input in182;
input in183;
input in184;
input in185;
input in186;
input in187;
input in188;
input in189;
input in190;
input in191;
input in192;
input in193;
input in194;
input in195;
input in196;
input in197;
input in198;
input in199;
input in200;
input in201;
input in202;
input in203;
input in204;
input in205;
input in206;
input in207;
input in208;
input in209;
input in210;
input in211;
input in212;
input in213;
input in214;
input in215;
input in216;
input in217;
input in218;
input in219;
input in220;
input in221;
input in222;
input in223;
input in224;
input in225;
input in226;
input in227;
input in228;
input in229;
input in230;
input in231;
input in232;
input in233;
input in234;
input in235;
input in236;
input in237;
input in238;
input in239;
input in240;
input in241;
input in242;
input in243;
input in244;
input in245;
input in246;
input in247;
input in248;
input in249;
input in250;
input in251;
input in252;
input in253;
input in254;
input in255;
output out0;
output out1;
output out2;
output out3;
output out4;
output out5;
output out6;
output out7;
output out8;
output out9;
output out10;
output out11;
output out12;
output out13;
output out14;
output out15;
output out16;
output out17;
output out18;
output out19;
output out20;
output out21;
output out22;
output out23;
output out24;
output out25;
output out26;
output out27;
output out28;
output out29;
output out30;
output out31;
output out32;
output out33;
output out34;
output out35;
output out36;
output out37;
output out38;
output out39;
output out40;
output out41;
output out42;
output out43;
output out44;
output out45;
output out46;
output out47;
output out48;
output out49;
output out50;
output out51;
output out52;
output out53;
output out54;
output out55;
output out56;
output out57;
output out58;
output out59;
output out60;
output out61;
output out62;
output out63;
output out64;
output out65;
output out66;
output out67;
output out68;
output out69;
output out70;
output out71;
output out72;
output out73;
output out74;
output out75;
output out76;
output out77;
output out78;
output out79;
output out80;
output out81;
output out82;
output out83;
output out84;
output out85;
output out86;
output out87;
output out88;
output out89;
output out90;
output out91;
output out92;
output out93;
output out94;
output out95;
output out96;
output out97;
output out98;
output out99;
output out100;
output out101;
output out102;
output out103;
output out104;
output out105;
output out106;
output out107;
output out108;
output out109;
output out110;
output out111;
output out112;
output out113;
output out114;
output out115;
output out116;
output out117;
output out118;
output out119;
output out120;
output out121;
output out122;
output out123;
output out124;
output out125;
output out126;
output out127;
output out128;
wire var0;
wire var1;
wire var2;
wire var3;
wire var4;
wire var5;
wire var6;
wire var7;
wire var8;
wire var9;
wire var10;
wire var11;
wire var12;
wire var13;
wire var14;
wire var15;
wire var16;
wire var17;
wire var18;
wire var19;
wire var20;
wire var21;
wire var22;
wire var23;
wire var24;
wire var25;
wire var26;
wire var27;
wire var28;
wire var29;
wire var30;
wire var31;
wire var32;
wire var33;
wire var34;
wire var35;
wire var36;
wire var37;
wire var38;
wire var39;
wire var40;
wire var41;
wire var42;
wire var43;
wire var44;
wire var45;
wire var46;
wire var47;
wire var48;
wire var49;
wire var50;
wire var51;
wire var52;
wire var53;
wire var54;
wire var55;
wire var56;
wire var57;
wire var58;
wire var59;
wire var60;
wire var61;
wire var62;
wire var63;
wire var64;
wire var65;
wire var66;
wire var67;
wire var68;
wire var69;
wire var70;
wire var71;
wire var72;
wire var73;
wire var74;
wire var75;
wire var76;
wire var77;
wire var78;
wire var79;
wire var80;
wire var81;
wire var82;
wire var83;
wire var84;
wire var85;
wire var86;
wire var87;
wire var88;
wire var89;
wire var90;
wire var91;
wire var92;
wire var93;
wire var94;
wire var95;
wire var96;
wire var97;
wire var98;
wire var99;
wire var100;
wire var101;
wire var102;
wire var103;
wire var104;
wire var105;
wire var106;
wire var107;
wire var108;
wire var109;
wire var110;
wire var111;
wire var112;
wire var113;
wire var114;
wire var115;
wire var116;
wire var117;
wire var118;
wire var119;
wire var120;
wire var121;
wire var122;
wire var123;
wire var124;
wire var125;
wire var126;
wire var127;
wire var128;
wire var129;
wire var130;
wire var131;
wire var132;
wire var133;
wire var134;
wire var135;
wire var136;
wire var137;
wire var138;
wire var139;
wire var140;
wire var141;
wire var142;
wire var143;
wire var144;
wire var145;
wire var146;
wire var147;
wire var148;
wire var149;
wire var150;
wire var151;
wire var152;
wire var153;
wire var154;
wire var155;
wire var156;
wire var157;
wire var158;
wire var159;
wire var160;
wire var161;
wire var162;
wire var163;
wire var164;
wire var165;
wire var166;
wire var167;
wire var168;
wire var169;
wire var170;
wire var171;
wire var172;
wire var173;
wire var174;
wire var175;
wire var176;
wire var177;
wire var178;
wire var179;
wire var180;
wire var181;
wire var182;
wire var183;
wire var184;
wire var185;
wire var186;
wire var187;
wire var188;
wire var189;
wire var190;
wire var191;
wire var192;
wire var193;
wire var194;
wire var195;
wire var196;
wire var197;
wire var198;
wire var199;
wire var200;
wire var201;
wire var202;
wire var203;
wire var204;
wire var205;
wire var206;
wire var207;
wire var208;
wire var209;
wire var210;
wire var211;
wire var212;
wire var213;
wire var214;
wire var215;
wire var216;
wire var217;
wire var218;
wire var219;
wire var220;
wire var221;
wire var222;
wire var223;
wire var224;
wire var225;
wire var226;
wire var227;
wire var228;
wire var229;
wire var230;
wire var231;
wire var232;
wire var233;
wire var234;
wire var235;
wire var236;
wire var237;
wire var238;
wire var239;
wire var240;
wire var241;
wire var242;
wire var243;
wire var244;
wire var245;
wire var246;
wire var247;
wire var248;
wire var249;
wire var250;
wire var251;
wire var252;
wire var253;
wire var254;
wire var255;
wire var256;
wire var257;
wire var258;
wire var259;
wire var260;
wire var261;
wire var262;
wire var263;
wire var264;
wire var265;
wire var266;
wire var267;
wire var268;
wire var269;
wire var270;
wire var271;
wire var272;
wire var273;
wire var274;
wire var275;
wire var276;
wire var277;
wire var278;
wire var279;
wire var280;
wire var281;
wire var282;
wire var283;
wire var284;
wire var285;
wire var286;
wire var287;
wire var288;
wire var289;
wire var290;
wire var291;
wire var292;
wire var293;
wire var294;
wire var295;
wire var296;
wire var297;
wire var298;
wire var299;
wire var300;
wire var301;
wire var302;
wire var303;
wire var304;
wire var305;
wire var306;
wire var307;
wire var308;
wire var309;
wire var310;
wire var311;
wire var312;
wire var313;
wire var314;
wire var315;
wire var316;
wire var317;
wire var318;
wire var319;
wire var320;
wire var321;
wire var322;
wire var323;
wire var324;
wire var325;
wire var326;
wire var327;
wire var328;
wire var329;
wire var330;
wire var331;
wire var332;
wire var333;
wire var334;
wire var335;
wire var336;
wire var337;
wire var338;
wire var339;
wire var340;
wire var341;
wire var342;
wire var343;
wire var344;
wire var345;
wire var346;
wire var347;
wire var348;
wire var349;
wire var350;
wire var351;
wire var352;
wire var353;
wire var354;
wire var355;
wire var356;
wire var357;
wire var358;
wire var359;
wire var360;
wire var361;
wire var362;
wire var363;
wire var364;
wire var365;
wire var366;
wire var367;
wire var368;
wire var369;
wire var370;
wire var371;
wire var372;
wire var373;
wire var374;
wire var375;
wire var376;
wire var377;
wire var378;
wire var379;
wire var380;
wire var381;
wire var382;
wire var383;
wire var384;
wire var385;
wire var386;
wire var387;
wire var388;
wire var389;
wire var390;
wire var391;
wire var392;
wire var393;
wire var394;
wire var395;
wire var396;
wire var397;
wire var398;
wire var399;
wire var400;
wire var401;
wire var402;
wire var403;
wire var404;
wire var405;
wire var406;
wire var407;
wire var408;
wire var409;
wire var410;
wire var411;
wire var412;
wire var413;
wire var414;
wire var415;
wire var416;
wire var417;
wire var418;
wire var419;
wire var420;
wire var421;
wire var422;
wire var423;
wire var424;
wire var425;
wire var426;
wire var427;
wire var428;
wire var429;
wire var430;
wire var431;
wire var432;
wire var433;
wire var434;
wire var435;
wire var436;
wire var437;
wire var438;
wire var439;
wire var440;
wire var441;
wire var442;
wire var443;
wire var444;
wire var445;
wire var446;
wire var447;
wire var448;
wire var449;
wire var450;
wire var451;
wire var452;
wire var453;
wire var454;
wire var455;
wire var456;
wire var457;
wire var458;
wire var459;
wire var460;
wire var461;
wire var462;
wire var463;
wire var464;
wire var465;
wire var466;
wire var467;
wire var468;
wire var469;
wire var470;
wire var471;
wire var472;
wire var473;
wire var474;
wire var475;
wire var476;
wire var477;
wire var478;
wire var479;
wire var480;
wire var481;
wire var482;
wire var483;
wire var484;
wire var485;
wire var486;
wire var487;
wire var488;
wire var489;
wire var490;
wire var491;
wire var492;
wire var493;
wire var494;
wire var495;
wire var496;
wire var497;
wire var498;
wire var499;
wire var500;
wire var501;
wire var502;
wire var503;
wire var504;
wire var505;
wire var506;
wire var507;
wire var508;
wire var509;
wire var510;
wire var511;
wire var512;
wire var513;
wire var514;
wire var515;
wire var516;
wire var517;
wire var518;
wire var519;
wire var520;
wire var521;
wire var522;
wire var523;
wire var524;
wire var525;
wire var526;
wire var527;
wire var528;
wire var529;
wire var530;
wire var531;
wire var532;
wire var533;
wire var534;
wire var535;
wire var536;
wire var537;
wire var538;
wire var539;
wire var540;
wire var541;
wire var542;
wire var543;
wire var544;
wire var545;
wire var546;
wire var547;
wire var548;
wire var549;
wire var550;
wire var551;
wire var552;
wire var553;
wire var554;
wire var555;
wire var556;
wire var557;
wire var558;
wire var559;
wire var560;
wire var561;
wire var562;
wire var563;
wire var564;
wire var565;
wire var566;
wire var567;
wire var568;
wire var569;
wire var570;
wire var571;
wire var572;
wire var573;
wire var574;
wire var575;
wire var576;
wire var577;
wire var578;
wire var579;
wire var580;
wire var581;
wire var582;
wire var583;
wire var584;
wire var585;
wire var586;
wire var587;
wire var588;
wire var589;
wire var590;
wire var591;
wire var592;
wire var593;
wire var594;
wire var595;
wire var596;
wire var597;
wire var598;
wire var599;
wire var600;
wire var601;
wire var602;
wire var603;
wire var604;
wire var605;
wire var606;
wire var607;
wire var608;
wire var609;
wire var610;
wire var611;
wire var612;
wire var613;
wire var614;
wire var615;
wire var616;
wire var617;
wire var618;
wire var619;
wire var620;
wire var621;
wire var622;
wire var623;
wire var624;
wire var625;
wire var626;
wire var627;
wire var628;
wire var629;
wire var630;
wire var631;
wire var632;
wire var633;
wire var634;
wire var635;
wire var636;
wire var637;
wire var638;
wire var639;
wire var640;
wire var641;
wire var642;
wire var643;
wire var644;
wire var645;
wire var646;
wire var647;
wire var648;
wire var649;
wire var650;
wire var651;
wire var652;
wire var653;
wire var654;
wire var655;
wire var656;
wire var657;
wire var658;
wire var659;
wire var660;
wire var661;
wire var662;
wire var663;
wire var664;
wire var665;
wire var666;
wire var667;
wire var668;
wire var669;
wire var670;
wire var671;
wire var672;
wire var673;
wire var674;
wire var675;
wire var676;
wire var677;
wire var678;
wire var679;
wire var680;
wire var681;
wire var682;
wire var683;
wire var684;
wire var685;
wire var686;
wire var687;
wire var688;
wire var689;
wire var690;
wire var691;
wire var692;
wire var693;
wire var694;
wire var695;
wire var696;
wire var697;
wire var698;
wire var699;
wire var700;
wire var701;
wire var702;
wire var703;
wire var704;
wire var705;
wire var706;
wire var707;
wire var708;
wire var709;
wire var710;
wire var711;
wire var712;
wire var713;
wire var714;
wire var715;
wire var716;
wire var717;
wire var718;
wire var719;
wire var720;
wire var721;
wire var722;
wire var723;
wire var724;
wire var725;
wire var726;
wire var727;
wire var728;
wire var729;
wire var730;
wire var731;
wire var732;
wire var733;
wire var734;
wire var735;
wire var736;
wire var737;
wire var738;
wire var739;
wire var740;
wire var741;
wire var742;
wire var743;
wire var744;
wire var745;
wire var746;
wire var747;
wire var748;
wire var749;
wire var750;
wire var751;
wire var752;
wire var753;
wire var754;
wire var755;
wire var756;
wire var757;
wire var758;
wire var759;
wire var760;
wire var761;
wire var762;
wire var763;
wire var764;
wire var765;
wire var766;
wire var767;
wire var768;
wire var769;
wire var770;
wire var771;
wire var772;
wire var773;
wire var774;
wire var775;
wire var776;
wire var777;
wire var778;
wire var779;
wire var780;
wire var781;
wire var782;
wire var783;
wire var784;
wire var785;
wire var786;
wire var787;
wire var788;
wire var789;
wire var790;
wire var791;
wire var792;
wire var793;
wire var794;
wire var795;
wire var796;
wire var797;
wire var798;
wire var799;
wire var800;
wire var801;
wire var802;
wire var803;
wire var804;
wire var805;
wire var806;
wire var807;
wire var808;
wire var809;
wire var810;
wire var811;
wire var812;
wire var813;
wire var814;
wire var815;
wire var816;
wire var817;
wire var818;
wire var819;
wire var820;
wire var821;
wire var822;
wire var823;
wire var824;
wire var825;
wire var826;
wire var827;
wire var828;
wire var829;
wire var830;
wire var831;
wire var832;
wire var833;
wire var834;
wire var835;
wire var836;
wire var837;
wire var838;
wire var839;
wire var840;
wire var841;
wire var842;
wire var843;
wire var844;
wire var845;
wire var846;
wire var847;
wire var848;
wire var849;
wire var850;
wire var851;
wire var852;
wire var853;
wire var854;
wire var855;
wire var856;
wire var857;
wire var858;
wire var859;
wire var860;
wire var861;
wire var862;
wire var863;
wire var864;
wire var865;
wire var866;
wire var867;
wire var868;
wire var869;
wire var870;
wire var871;
wire var872;
wire var873;
wire var874;
wire var875;
wire var876;
wire var877;
wire var878;
wire var879;
wire var880;
wire var881;
wire var882;
wire var883;
wire var884;
wire var885;
wire var886;
wire var887;
wire var888;
wire var889;
wire var890;
wire var891;
wire var892;
wire var893;
wire var894;
wire var895;
wire var896;
wire var897;
wire var898;
wire var899;
wire var900;
wire var901;
wire var902;
wire var903;
wire var904;
wire var905;
wire var906;
wire var907;
wire var908;
wire var909;
wire var910;
wire var911;
wire var912;
wire var913;
wire var914;
wire var915;
wire var916;
wire var917;
wire var918;
wire var919;
wire var920;
wire var921;
wire var922;
wire var923;
wire var924;
wire var925;
wire var926;
wire var927;
wire var928;
wire var929;
wire var930;
wire var931;
wire var932;
wire var933;
wire var934;
wire var935;
wire var936;
wire var937;
wire var938;
wire var939;
wire var940;
wire var941;
wire var942;
wire var943;
wire var944;
wire var945;
wire var946;
wire var947;
wire var948;
wire var949;
wire var950;
wire var951;
wire var952;
wire var953;
wire var954;
wire var955;
wire var956;
wire var957;
wire var958;
wire var959;
wire var960;
wire var961;
wire var962;
wire var963;
wire var964;
wire var965;
wire var966;
wire var967;
wire var968;
wire var969;
wire var970;
wire var971;
wire var972;
wire var973;
wire var974;
wire var975;
wire var976;
wire var977;
wire var978;
wire var979;
wire var980;
wire var981;
wire var982;
wire var983;
wire var984;
wire var985;
wire var986;
wire var987;
wire var988;
wire var989;
wire var990;
wire var991;
wire var992;
wire var993;
wire var994;
wire var995;
wire var996;
wire var997;
wire var998;
wire var999;
wire var1000;
wire var1001;
wire var1002;
wire var1003;
wire var1004;
wire var1005;
wire var1006;
wire var1007;
wire var1008;
wire var1009;
wire var1010;
wire var1011;
wire var1012;
wire var1013;
wire var1014;
wire var1015;
wire var1016;
wire var1017;
wire var1018;
wire var1019;
wire var1020;
wire var1021;
wire var1022;
wire var1023;
wire var1024;
wire var1025;
wire var1026;
wire var1027;
wire var1028;
wire var1029;
wire var1030;
wire var1031;
wire var1032;
wire var1033;
wire var1034;
wire var1035;
wire var1036;
wire var1037;
wire var1038;
wire var1039;
wire var1040;
wire var1041;
wire var1042;
wire var1043;
wire var1044;
wire var1045;
wire var1046;
wire var1047;
wire var1048;
wire var1049;
wire var1050;
wire var1051;
wire var1052;
wire var1053;
wire var1054;
wire var1055;
wire var1056;
wire var1057;
wire var1058;
wire var1059;
wire var1060;
wire var1061;
wire var1062;
wire var1063;
wire var1064;
wire var1065;
wire var1066;
wire var1067;
wire var1068;
wire var1069;
wire var1070;
wire var1071;
wire var1072;
wire var1073;
wire var1074;
wire var1075;
wire var1076;
wire var1077;
wire var1078;
wire var1079;
wire var1080;
wire var1081;
wire var1082;
wire var1083;
wire var1084;
wire var1085;
wire var1086;
wire var1087;
wire var1088;
wire var1089;
wire var1090;
wire var1091;
wire var1092;
wire var1093;
wire var1094;
wire var1095;
wire var1096;
wire var1097;
wire var1098;
wire var1099;
wire var1100;
wire var1101;
wire var1102;
wire var1103;
wire var1104;
wire var1105;
wire var1106;
wire var1107;
wire var1108;
wire var1109;
wire var1110;
wire var1111;
wire var1112;
wire var1113;
wire var1114;
wire var1115;
wire var1116;
wire var1117;
wire var1118;
wire var1119;
wire var1120;
wire var1121;
wire var1122;
wire var1123;
wire var1124;
wire var1125;
wire var1126;
wire var1127;
wire var1128;
wire var1129;
wire var1130;
wire var1131;
wire var1132;
wire var1133;
wire var1134;
wire var1135;
wire var1136;
wire var1137;
wire var1138;
wire var1139;
wire var1140;
wire var1141;
wire var1142;
wire var1143;
wire var1144;
wire var1145;
wire var1146;
wire var1147;
wire var1148;
wire var1149;
wire var1150;
wire var1151;
wire var1152;
wire var1153;
wire var1154;
wire var1155;
wire var1156;
wire var1157;
wire var1158;
wire var1159;
wire var1160;
wire var1161;
wire var1162;
wire var1163;
wire var1164;
wire var1165;
wire var1166;
wire var1167;
wire var1168;
wire var1169;
wire var1170;
wire var1171;
wire var1172;
wire var1173;
wire var1174;
wire var1175;
wire var1176;
wire var1177;
wire var1178;
wire var1179;
wire var1180;
wire var1181;
wire var1182;
wire var1183;
wire var1184;
wire var1185;
wire var1186;
wire var1187;
wire var1188;
wire var1189;
wire var1190;
wire var1191;
wire var1192;
wire var1193;
wire var1194;
wire var1195;
wire var1196;
wire var1197;
wire var1198;
wire var1199;
wire var1200;
wire var1201;
wire var1202;
wire var1203;
wire var1204;
wire var1205;
wire var1206;
wire var1207;
wire var1208;
wire var1209;
wire var1210;
wire var1211;
wire var1212;
wire var1213;
wire var1214;
wire var1215;
wire var1216;
wire var1217;
wire var1218;
wire var1219;
wire var1220;
wire var1221;
wire var1222;
wire var1223;
wire var1224;
wire var1225;
wire var1226;
wire var1227;
wire var1228;
wire var1229;
wire var1230;
wire var1231;
wire var1232;
wire var1233;
wire var1234;
wire var1235;
wire var1236;
wire var1237;
wire var1238;
wire var1239;
wire var1240;
wire var1241;
wire var1242;
wire var1243;
wire var1244;
wire var1245;
wire var1246;
wire var1247;
wire var1248;
wire var1249;
wire var1250;
wire var1251;
wire var1252;
wire var1253;
wire var1254;
wire var1255;
wire var1256;
wire var1257;
wire var1258;
wire var1259;
wire var1260;
wire var1261;
wire var1262;
wire var1263;
wire var1264;
wire var1265;
wire var1266;
wire var1267;
wire var1268;
wire var1269;
wire var1270;
wire var1271;
wire var1272;
wire var1273;
wire var1274;
wire var1275;
assign var0 = in255 & in127;
assign var1 = in254 & in126;
assign var2 = in253 & in125;
assign var3 = in252 & in124;
assign var4 = in251 & in123;
assign var5 = in250 & in122;
assign var6 = in249 & in121;
assign var7 = in248 & in120;
assign var8 = in247 & in119;
assign var9 = in246 & in118;
assign var10 = in245 & in117;
assign var11 = in244 & in116;
assign var12 = in243 & in115;
assign var13 = in242 & in114;
assign var14 = in241 & in113;
assign var15 = in240 & in112;
assign var16 = in239 & in111;
assign var17 = in238 & in110;
assign var18 = in237 & in109;
assign var19 = in236 & in108;
assign var20 = in235 & in107;
assign var21 = in234 & in106;
assign var22 = in233 & in105;
assign var23 = in232 & in104;
assign var24 = in231 & in103;
assign var25 = in230 & in102;
assign var26 = in229 & in101;
assign var27 = in228 & in100;
assign var28 = in227 & in99;
assign var29 = in226 & in98;
assign var30 = in225 & in97;
assign var31 = in224 & in96;
assign var32 = in223 & in95;
assign var33 = in222 & in94;
assign var34 = in221 & in93;
assign var35 = in220 & in92;
assign var36 = in219 & in91;
assign var37 = in218 & in90;
assign var38 = in217 & in89;
assign var39 = in216 & in88;
assign var40 = in215 & in87;
assign var41 = in214 & in86;
assign var42 = in213 & in85;
assign var43 = in212 & in84;
assign var44 = in211 & in83;
assign var45 = in210 & in82;
assign var46 = in209 & in81;
assign var47 = in208 & in80;
assign var48 = in207 & in79;
assign var49 = in206 & in78;
assign var50 = in205 & in77;
assign var51 = in204 & in76;
assign var52 = in203 & in75;
assign var53 = in202 & in74;
assign var54 = in201 & in73;
assign var55 = in200 & in72;
assign var56 = in199 & in71;
assign var57 = in198 & in70;
assign var58 = in197 & in69;
assign var59 = in196 & in68;
assign var60 = in195 & in67;
assign var61 = in194 & in66;
assign var62 = in193 & in65;
assign var63 = in192 & in64;
assign var64 = in191 & in63;
assign var65 = in190 & in62;
assign var66 = in189 & in61;
assign var67 = in188 & in60;
assign var68 = in187 & in59;
assign var69 = in186 & in58;
assign var70 = in185 & in57;
assign var71 = in184 & in56;
assign var72 = in183 & in55;
assign var73 = in182 & in54;
assign var74 = in181 & in53;
assign var75 = in180 & in52;
assign var76 = in179 & in51;
assign var77 = in178 & in50;
assign var78 = in177 & in49;
assign var79 = in176 & in48;
assign var80 = in175 & in47;
assign var81 = in174 & in46;
assign var82 = in173 & in45;
assign var83 = in172 & in44;
assign var84 = in171 & in43;
assign var85 = in170 & in42;
assign var86 = in169 & in41;
assign var87 = in168 & in40;
assign var88 = in167 & in39;
assign var89 = in166 & in38;
assign var90 = in165 & in37;
assign var91 = in164 & in36;
assign var92 = in163 & in35;
assign var93 = in162 & in34;
assign var94 = in161 & in33;
assign var95 = in160 & in32;
assign var96 = in159 & in31;
assign var97 = in158 & in30;
assign var98 = in157 & in29;
assign var99 = in156 & in28;
assign var100 = in155 & in27;
assign var101 = in154 & in26;
assign var102 = in153 & in25;
assign var103 = in152 & in24;
assign var104 = in151 & in23;
assign var105 = in150 & in22;
assign var106 = in149 & in21;
assign var107 = in148 & in20;
assign var108 = in147 & in19;
assign var109 = in146 & in18;
assign var110 = in145 & in17;
assign var111 = in144 & in16;
assign var112 = in143 & in15;
assign var113 = in142 & in14;
assign var114 = in141 & in13;
assign var115 = in140 & in12;
assign var116 = in139 & in11;
assign var117 = in138 & in10;
assign var118 = in137 & in9;
assign var119 = in136 & in8;
assign var120 = in135 & in7;
assign var121 = in134 & in6;
assign var122 = in133 & in5;
assign var123 = in132 & in4;
assign var124 = in131 & in3;
assign var125 = in130 & in2;
assign var126 = in129 & in1;
assign var127 = in128 & in0;
assign var128 = in255 ^ in127;
assign var129 = in254 ^ in126;
assign var130 = in253 ^ in125;
assign var131 = in252 ^ in124;
assign var132 = in251 ^ in123;
assign var133 = in250 ^ in122;
assign var134 = in249 ^ in121;
assign var135 = in248 ^ in120;
assign var136 = in247 ^ in119;
assign var137 = in246 ^ in118;
assign var138 = in245 ^ in117;
assign var139 = in244 ^ in116;
assign var140 = in243 ^ in115;
assign var141 = in242 ^ in114;
assign var142 = in241 ^ in113;
assign var143 = in240 ^ in112;
assign var144 = in239 ^ in111;
assign var145 = in238 ^ in110;
assign var146 = in237 ^ in109;
assign var147 = in236 ^ in108;
assign var148 = in235 ^ in107;
assign var149 = in234 ^ in106;
assign var150 = in233 ^ in105;
assign var151 = in232 ^ in104;
assign var152 = in231 ^ in103;
assign var153 = in230 ^ in102;
assign var154 = in229 ^ in101;
assign var155 = in228 ^ in100;
assign var156 = in227 ^ in99;
assign var157 = in226 ^ in98;
assign var158 = in225 ^ in97;
assign var159 = in224 ^ in96;
assign var160 = in223 ^ in95;
assign var161 = in222 ^ in94;
assign var162 = in221 ^ in93;
assign var163 = in220 ^ in92;
assign var164 = in219 ^ in91;
assign var165 = in218 ^ in90;
assign var166 = in217 ^ in89;
assign var167 = in216 ^ in88;
assign var168 = in215 ^ in87;
assign var169 = in214 ^ in86;
assign var170 = in213 ^ in85;
assign var171 = in212 ^ in84;
assign var172 = in211 ^ in83;
assign var173 = in210 ^ in82;
assign var174 = in209 ^ in81;
assign var175 = in208 ^ in80;
assign var176 = in207 ^ in79;
assign var177 = in206 ^ in78;
assign var178 = in205 ^ in77;
assign var179 = in204 ^ in76;
assign var180 = in203 ^ in75;
assign var181 = in202 ^ in74;
assign var182 = in201 ^ in73;
assign var183 = in200 ^ in72;
assign var184 = in199 ^ in71;
assign var185 = in198 ^ in70;
assign var186 = in197 ^ in69;
assign var187 = in196 ^ in68;
assign var188 = in195 ^ in67;
assign var189 = in194 ^ in66;
assign var190 = in193 ^ in65;
assign var191 = in192 ^ in64;
assign var192 = in191 ^ in63;
assign var193 = in190 ^ in62;
assign var194 = in189 ^ in61;
assign var195 = in188 ^ in60;
assign var196 = in187 ^ in59;
assign var197 = in186 ^ in58;
assign var198 = in185 ^ in57;
assign var199 = in184 ^ in56;
assign var200 = in183 ^ in55;
assign var201 = in182 ^ in54;
assign var202 = in181 ^ in53;
assign var203 = in180 ^ in52;
assign var204 = in179 ^ in51;
assign var205 = in178 ^ in50;
assign var206 = in177 ^ in49;
assign var207 = in176 ^ in48;
assign var208 = in175 ^ in47;
assign var209 = in174 ^ in46;
assign var210 = in173 ^ in45;
assign var211 = in172 ^ in44;
assign var212 = in171 ^ in43;
assign var213 = in170 ^ in42;
assign var214 = in169 ^ in41;
assign var215 = in168 ^ in40;
assign var216 = in167 ^ in39;
assign var217 = in166 ^ in38;
assign var218 = in165 ^ in37;
assign var219 = in164 ^ in36;
assign var220 = in163 ^ in35;
assign var221 = in162 ^ in34;
assign var222 = in161 ^ in33;
assign var223 = in160 ^ in32;
assign var224 = in159 ^ in31;
assign var225 = in158 ^ in30;
assign var226 = in157 ^ in29;
assign var227 = in156 ^ in28;
assign var228 = in155 ^ in27;
assign var229 = in154 ^ in26;
assign var230 = in153 ^ in25;
assign var231 = in152 ^ in24;
assign var232 = in151 ^ in23;
assign var233 = in150 ^ in22;
assign var234 = in149 ^ in21;
assign var235 = in148 ^ in20;
assign var236 = in147 ^ in19;
assign var237 = in146 ^ in18;
assign var238 = in145 ^ in17;
assign var239 = in144 ^ in16;
assign var240 = in143 ^ in15;
assign var241 = in142 ^ in14;
assign var242 = in141 ^ in13;
assign var243 = in140 ^ in12;
assign var244 = in139 ^ in11;
assign var245 = in138 ^ in10;
assign var246 = in137 ^ in9;
assign var247 = in136 ^ in8;
assign var248 = in135 ^ in7;
assign var249 = in134 ^ in6;
assign var250 = in133 ^ in5;
assign var251 = in132 ^ in4;
assign var252 = in131 ^ in3;
assign var253 = in130 ^ in2;
assign var254 = in129 ^ in1;
assign var255 = in128 ^ in0;
assign var256 = var255 & var126;
assign var257 = var127 | var256;
assign var258 = var255 & var254;
assign var259 = var253 & var124;
assign var260 = var125 | var259;
assign var261 = var253 & var252;
assign var262 = var251 & var122;
assign var263 = var123 | var262;
assign var264 = var251 & var250;
assign var265 = var249 & var120;
assign var266 = var121 | var265;
assign var267 = var249 & var248;
assign var268 = var247 & var118;
assign var269 = var119 | var268;
assign var270 = var247 & var246;
assign var271 = var245 & var116;
assign var272 = var117 | var271;
assign var273 = var245 & var244;
assign var274 = var243 & var114;
assign var275 = var115 | var274;
assign var276 = var243 & var242;
assign var277 = var241 & var112;
assign var278 = var113 | var277;
assign var279 = var241 & var240;
assign var280 = var239 & var110;
assign var281 = var111 | var280;
assign var282 = var239 & var238;
assign var283 = var237 & var108;
assign var284 = var109 | var283;
assign var285 = var237 & var236;
assign var286 = var235 & var106;
assign var287 = var107 | var286;
assign var288 = var235 & var234;
assign var289 = var233 & var104;
assign var290 = var105 | var289;
assign var291 = var233 & var232;
assign var292 = var231 & var102;
assign var293 = var103 | var292;
assign var294 = var231 & var230;
assign var295 = var229 & var100;
assign var296 = var101 | var295;
assign var297 = var229 & var228;
assign var298 = var227 & var98;
assign var299 = var99 | var298;
assign var300 = var227 & var226;
assign var301 = var225 & var96;
assign var302 = var97 | var301;
assign var303 = var225 & var224;
assign var304 = var223 & var94;
assign var305 = var95 | var304;
assign var306 = var223 & var222;
assign var307 = var221 & var92;
assign var308 = var93 | var307;
assign var309 = var221 & var220;
assign var310 = var219 & var90;
assign var311 = var91 | var310;
assign var312 = var219 & var218;
assign var313 = var217 & var88;
assign var314 = var89 | var313;
assign var315 = var217 & var216;
assign var316 = var215 & var86;
assign var317 = var87 | var316;
assign var318 = var215 & var214;
assign var319 = var213 & var84;
assign var320 = var85 | var319;
assign var321 = var213 & var212;
assign var322 = var211 & var82;
assign var323 = var83 | var322;
assign var324 = var211 & var210;
assign var325 = var209 & var80;
assign var326 = var81 | var325;
assign var327 = var209 & var208;
assign var328 = var207 & var78;
assign var329 = var79 | var328;
assign var330 = var207 & var206;
assign var331 = var205 & var76;
assign var332 = var77 | var331;
assign var333 = var205 & var204;
assign var334 = var203 & var74;
assign var335 = var75 | var334;
assign var336 = var203 & var202;
assign var337 = var201 & var72;
assign var338 = var73 | var337;
assign var339 = var201 & var200;
assign var340 = var199 & var70;
assign var341 = var71 | var340;
assign var342 = var199 & var198;
assign var343 = var197 & var68;
assign var344 = var69 | var343;
assign var345 = var197 & var196;
assign var346 = var195 & var66;
assign var347 = var67 | var346;
assign var348 = var195 & var194;
assign var349 = var193 & var64;
assign var350 = var65 | var349;
assign var351 = var193 & var192;
assign var352 = var191 & var62;
assign var353 = var63 | var352;
assign var354 = var191 & var190;
assign var355 = var189 & var60;
assign var356 = var61 | var355;
assign var357 = var189 & var188;
assign var358 = var187 & var58;
assign var359 = var59 | var358;
assign var360 = var187 & var186;
assign var361 = var185 & var56;
assign var362 = var57 | var361;
assign var363 = var185 & var184;
assign var364 = var183 & var54;
assign var365 = var55 | var364;
assign var366 = var183 & var182;
assign var367 = var181 & var52;
assign var368 = var53 | var367;
assign var369 = var181 & var180;
assign var370 = var179 & var50;
assign var371 = var51 | var370;
assign var372 = var179 & var178;
assign var373 = var177 & var48;
assign var374 = var49 | var373;
assign var375 = var177 & var176;
assign var376 = var175 & var46;
assign var377 = var47 | var376;
assign var378 = var175 & var174;
assign var379 = var173 & var44;
assign var380 = var45 | var379;
assign var381 = var173 & var172;
assign var382 = var171 & var42;
assign var383 = var43 | var382;
assign var384 = var171 & var170;
assign var385 = var169 & var40;
assign var386 = var41 | var385;
assign var387 = var169 & var168;
assign var388 = var167 & var38;
assign var389 = var39 | var388;
assign var390 = var167 & var166;
assign var391 = var165 & var36;
assign var392 = var37 | var391;
assign var393 = var165 & var164;
assign var394 = var163 & var34;
assign var395 = var35 | var394;
assign var396 = var163 & var162;
assign var397 = var161 & var32;
assign var398 = var33 | var397;
assign var399 = var161 & var160;
assign var400 = var159 & var30;
assign var401 = var31 | var400;
assign var402 = var159 & var158;
assign var403 = var157 & var28;
assign var404 = var29 | var403;
assign var405 = var157 & var156;
assign var406 = var155 & var26;
assign var407 = var27 | var406;
assign var408 = var155 & var154;
assign var409 = var153 & var24;
assign var410 = var25 | var409;
assign var411 = var153 & var152;
assign var412 = var151 & var22;
assign var413 = var23 | var412;
assign var414 = var151 & var150;
assign var415 = var149 & var20;
assign var416 = var21 | var415;
assign var417 = var149 & var148;
assign var418 = var147 & var18;
assign var419 = var19 | var418;
assign var420 = var147 & var146;
assign var421 = var145 & var16;
assign var422 = var17 | var421;
assign var423 = var145 & var144;
assign var424 = var143 & var14;
assign var425 = var15 | var424;
assign var426 = var143 & var142;
assign var427 = var141 & var12;
assign var428 = var13 | var427;
assign var429 = var141 & var140;
assign var430 = var139 & var10;
assign var431 = var11 | var430;
assign var432 = var139 & var138;
assign var433 = var137 & var8;
assign var434 = var9 | var433;
assign var435 = var137 & var136;
assign var436 = var135 & var6;
assign var437 = var7 | var436;
assign var438 = var135 & var134;
assign var439 = var133 & var4;
assign var440 = var5 | var439;
assign var441 = var133 & var132;
assign var442 = var131 & var2;
assign var443 = var3 | var442;
assign var444 = var131 & var130;
assign var445 = var129 & var0;
assign var446 = var1 | var445;
assign var447 = var258 & var260;
assign var448 = var257 | var447;
assign var449 = var258 & var261;
assign var450 = var264 & var266;
assign var451 = var263 | var450;
assign var452 = var264 & var267;
assign var453 = var270 & var272;
assign var454 = var269 | var453;
assign var455 = var270 & var273;
assign var456 = var276 & var278;
assign var457 = var275 | var456;
assign var458 = var276 & var279;
assign var459 = var282 & var284;
assign var460 = var281 | var459;
assign var461 = var282 & var285;
assign var462 = var288 & var290;
assign var463 = var287 | var462;
assign var464 = var288 & var291;
assign var465 = var294 & var296;
assign var466 = var293 | var465;
assign var467 = var294 & var297;
assign var468 = var300 & var302;
assign var469 = var299 | var468;
assign var470 = var300 & var303;
assign var471 = var306 & var308;
assign var472 = var305 | var471;
assign var473 = var306 & var309;
assign var474 = var312 & var314;
assign var475 = var311 | var474;
assign var476 = var312 & var315;
assign var477 = var318 & var320;
assign var478 = var317 | var477;
assign var479 = var318 & var321;
assign var480 = var324 & var326;
assign var481 = var323 | var480;
assign var482 = var324 & var327;
assign var483 = var330 & var332;
assign var484 = var329 | var483;
assign var485 = var330 & var333;
assign var486 = var336 & var338;
assign var487 = var335 | var486;
assign var488 = var336 & var339;
assign var489 = var342 & var344;
assign var490 = var341 | var489;
assign var491 = var342 & var345;
assign var492 = var348 & var350;
assign var493 = var347 | var492;
assign var494 = var348 & var351;
assign var495 = var354 & var356;
assign var496 = var353 | var495;
assign var497 = var354 & var357;
assign var498 = var360 & var362;
assign var499 = var359 | var498;
assign var500 = var360 & var363;
assign var501 = var366 & var368;
assign var502 = var365 | var501;
assign var503 = var366 & var369;
assign var504 = var372 & var374;
assign var505 = var371 | var504;
assign var506 = var372 & var375;
assign var507 = var378 & var380;
assign var508 = var377 | var507;
assign var509 = var378 & var381;
assign var510 = var384 & var386;
assign var511 = var383 | var510;
assign var512 = var384 & var387;
assign var513 = var390 & var392;
assign var514 = var389 | var513;
assign var515 = var390 & var393;
assign var516 = var396 & var398;
assign var517 = var395 | var516;
assign var518 = var396 & var399;
assign var519 = var402 & var404;
assign var520 = var401 | var519;
assign var521 = var402 & var405;
assign var522 = var408 & var410;
assign var523 = var407 | var522;
assign var524 = var408 & var411;
assign var525 = var414 & var416;
assign var526 = var413 | var525;
assign var527 = var414 & var417;
assign var528 = var420 & var422;
assign var529 = var419 | var528;
assign var530 = var420 & var423;
assign var531 = var426 & var428;
assign var532 = var425 | var531;
assign var533 = var426 & var429;
assign var534 = var432 & var434;
assign var535 = var431 | var534;
assign var536 = var432 & var435;
assign var537 = var438 & var440;
assign var538 = var437 | var537;
assign var539 = var438 & var441;
assign var540 = var444 & var446;
assign var541 = var443 | var540;
assign var542 = var449 & var451;
assign var543 = var448 | var542;
assign var544 = var449 & var452;
assign var545 = var261 & var451;
assign var546 = var260 | var545;
assign var547 = var261 & var452;
assign var548 = var455 & var457;
assign var549 = var454 | var548;
assign var550 = var455 & var458;
assign var551 = var273 & var457;
assign var552 = var272 | var551;
assign var553 = var273 & var458;
assign var554 = var461 & var463;
assign var555 = var460 | var554;
assign var556 = var461 & var464;
assign var557 = var285 & var463;
assign var558 = var284 | var557;
assign var559 = var285 & var464;
assign var560 = var467 & var469;
assign var561 = var466 | var560;
assign var562 = var467 & var470;
assign var563 = var297 & var469;
assign var564 = var296 | var563;
assign var565 = var297 & var470;
assign var566 = var473 & var475;
assign var567 = var472 | var566;
assign var568 = var473 & var476;
assign var569 = var309 & var475;
assign var570 = var308 | var569;
assign var571 = var309 & var476;
assign var572 = var479 & var481;
assign var573 = var478 | var572;
assign var574 = var479 & var482;
assign var575 = var321 & var481;
assign var576 = var320 | var575;
assign var577 = var321 & var482;
assign var578 = var485 & var487;
assign var579 = var484 | var578;
assign var580 = var485 & var488;
assign var581 = var333 & var487;
assign var582 = var332 | var581;
assign var583 = var333 & var488;
assign var584 = var491 & var493;
assign var585 = var490 | var584;
assign var586 = var491 & var494;
assign var587 = var345 & var493;
assign var588 = var344 | var587;
assign var589 = var345 & var494;
assign var590 = var497 & var499;
assign var591 = var496 | var590;
assign var592 = var497 & var500;
assign var593 = var357 & var499;
assign var594 = var356 | var593;
assign var595 = var357 & var500;
assign var596 = var503 & var505;
assign var597 = var502 | var596;
assign var598 = var503 & var506;
assign var599 = var369 & var505;
assign var600 = var368 | var599;
assign var601 = var369 & var506;
assign var602 = var509 & var511;
assign var603 = var508 | var602;
assign var604 = var509 & var512;
assign var605 = var381 & var511;
assign var606 = var380 | var605;
assign var607 = var381 & var512;
assign var608 = var515 & var517;
assign var609 = var514 | var608;
assign var610 = var515 & var518;
assign var611 = var393 & var517;
assign var612 = var392 | var611;
assign var613 = var393 & var518;
assign var614 = var521 & var523;
assign var615 = var520 | var614;
assign var616 = var521 & var524;
assign var617 = var405 & var523;
assign var618 = var404 | var617;
assign var619 = var405 & var524;
assign var620 = var527 & var529;
assign var621 = var526 | var620;
assign var622 = var527 & var530;
assign var623 = var417 & var529;
assign var624 = var416 | var623;
assign var625 = var417 & var530;
assign var626 = var533 & var535;
assign var627 = var532 | var626;
assign var628 = var533 & var536;
assign var629 = var429 & var535;
assign var630 = var428 | var629;
assign var631 = var429 & var536;
assign var632 = var539 & var541;
assign var633 = var538 | var632;
assign var634 = var441 & var541;
assign var635 = var440 | var634;
assign var636 = var544 & var549;
assign var637 = var543 | var636;
assign var638 = var544 & var550;
assign var639 = var547 & var549;
assign var640 = var546 | var639;
assign var641 = var547 & var550;
assign var642 = var452 & var549;
assign var643 = var451 | var642;
assign var644 = var452 & var550;
assign var645 = var267 & var549;
assign var646 = var266 | var645;
assign var647 = var267 & var550;
assign var648 = var556 & var561;
assign var649 = var555 | var648;
assign var650 = var556 & var562;
assign var651 = var559 & var561;
assign var652 = var558 | var651;
assign var653 = var559 & var562;
assign var654 = var464 & var561;
assign var655 = var463 | var654;
assign var656 = var464 & var562;
assign var657 = var291 & var561;
assign var658 = var290 | var657;
assign var659 = var291 & var562;
assign var660 = var568 & var573;
assign var661 = var567 | var660;
assign var662 = var568 & var574;
assign var663 = var571 & var573;
assign var664 = var570 | var663;
assign var665 = var571 & var574;
assign var666 = var476 & var573;
assign var667 = var475 | var666;
assign var668 = var476 & var574;
assign var669 = var315 & var573;
assign var670 = var314 | var669;
assign var671 = var315 & var574;
assign var672 = var580 & var585;
assign var673 = var579 | var672;
assign var674 = var580 & var586;
assign var675 = var583 & var585;
assign var676 = var582 | var675;
assign var677 = var583 & var586;
assign var678 = var488 & var585;
assign var679 = var487 | var678;
assign var680 = var488 & var586;
assign var681 = var339 & var585;
assign var682 = var338 | var681;
assign var683 = var339 & var586;
assign var684 = var592 & var597;
assign var685 = var591 | var684;
assign var686 = var592 & var598;
assign var687 = var595 & var597;
assign var688 = var594 | var687;
assign var689 = var595 & var598;
assign var690 = var500 & var597;
assign var691 = var499 | var690;
assign var692 = var500 & var598;
assign var693 = var363 & var597;
assign var694 = var362 | var693;
assign var695 = var363 & var598;
assign var696 = var604 & var609;
assign var697 = var603 | var696;
assign var698 = var604 & var610;
assign var699 = var607 & var609;
assign var700 = var606 | var699;
assign var701 = var607 & var610;
assign var702 = var512 & var609;
assign var703 = var511 | var702;
assign var704 = var512 & var610;
assign var705 = var387 & var609;
assign var706 = var386 | var705;
assign var707 = var387 & var610;
assign var708 = var616 & var621;
assign var709 = var615 | var708;
assign var710 = var616 & var622;
assign var711 = var619 & var621;
assign var712 = var618 | var711;
assign var713 = var619 & var622;
assign var714 = var524 & var621;
assign var715 = var523 | var714;
assign var716 = var524 & var622;
assign var717 = var411 & var621;
assign var718 = var410 | var717;
assign var719 = var411 & var622;
assign var720 = var628 & var633;
assign var721 = var627 | var720;
assign var722 = var631 & var633;
assign var723 = var630 | var722;
assign var724 = var536 & var633;
assign var725 = var535 | var724;
assign var726 = var435 & var633;
assign var727 = var434 | var726;
assign var728 = var638 & var649;
assign var729 = var637 | var728;
assign var730 = var638 & var650;
assign var731 = var641 & var649;
assign var732 = var640 | var731;
assign var733 = var641 & var650;
assign var734 = var644 & var649;
assign var735 = var643 | var734;
assign var736 = var644 & var650;
assign var737 = var647 & var649;
assign var738 = var646 | var737;
assign var739 = var647 & var650;
assign var740 = var550 & var649;
assign var741 = var549 | var740;
assign var742 = var550 & var650;
assign var743 = var553 & var649;
assign var744 = var552 | var743;
assign var745 = var553 & var650;
assign var746 = var458 & var649;
assign var747 = var457 | var746;
assign var748 = var458 & var650;
assign var749 = var279 & var649;
assign var750 = var278 | var749;
assign var751 = var279 & var650;
assign var752 = var662 & var673;
assign var753 = var661 | var752;
assign var754 = var662 & var674;
assign var755 = var665 & var673;
assign var756 = var664 | var755;
assign var757 = var665 & var674;
assign var758 = var668 & var673;
assign var759 = var667 | var758;
assign var760 = var668 & var674;
assign var761 = var671 & var673;
assign var762 = var670 | var761;
assign var763 = var671 & var674;
assign var764 = var574 & var673;
assign var765 = var573 | var764;
assign var766 = var574 & var674;
assign var767 = var577 & var673;
assign var768 = var576 | var767;
assign var769 = var577 & var674;
assign var770 = var482 & var673;
assign var771 = var481 | var770;
assign var772 = var482 & var674;
assign var773 = var327 & var673;
assign var774 = var326 | var773;
assign var775 = var327 & var674;
assign var776 = var686 & var697;
assign var777 = var685 | var776;
assign var778 = var686 & var698;
assign var779 = var689 & var697;
assign var780 = var688 | var779;
assign var781 = var689 & var698;
assign var782 = var692 & var697;
assign var783 = var691 | var782;
assign var784 = var692 & var698;
assign var785 = var695 & var697;
assign var786 = var694 | var785;
assign var787 = var695 & var698;
assign var788 = var598 & var697;
assign var789 = var597 | var788;
assign var790 = var598 & var698;
assign var791 = var601 & var697;
assign var792 = var600 | var791;
assign var793 = var601 & var698;
assign var794 = var506 & var697;
assign var795 = var505 | var794;
assign var796 = var506 & var698;
assign var797 = var375 & var697;
assign var798 = var374 | var797;
assign var799 = var375 & var698;
assign var800 = var710 & var721;
assign var801 = var709 | var800;
assign var802 = var713 & var721;
assign var803 = var712 | var802;
assign var804 = var716 & var721;
assign var805 = var715 | var804;
assign var806 = var719 & var721;
assign var807 = var718 | var806;
assign var808 = var622 & var721;
assign var809 = var621 | var808;
assign var810 = var625 & var721;
assign var811 = var624 | var810;
assign var812 = var530 & var721;
assign var813 = var529 | var812;
assign var814 = var423 & var721;
assign var815 = var422 | var814;
assign var816 = var730 & var753;
assign var817 = var729 | var816;
assign var818 = var730 & var754;
assign var819 = var733 & var753;
assign var820 = var732 | var819;
assign var821 = var733 & var754;
assign var822 = var736 & var753;
assign var823 = var735 | var822;
assign var824 = var736 & var754;
assign var825 = var739 & var753;
assign var826 = var738 | var825;
assign var827 = var739 & var754;
assign var828 = var742 & var753;
assign var829 = var741 | var828;
assign var830 = var742 & var754;
assign var831 = var745 & var753;
assign var832 = var744 | var831;
assign var833 = var745 & var754;
assign var834 = var748 & var753;
assign var835 = var747 | var834;
assign var836 = var748 & var754;
assign var837 = var751 & var753;
assign var838 = var750 | var837;
assign var839 = var751 & var754;
assign var840 = var650 & var753;
assign var841 = var649 | var840;
assign var842 = var650 & var754;
assign var843 = var653 & var753;
assign var844 = var652 | var843;
assign var845 = var653 & var754;
assign var846 = var656 & var753;
assign var847 = var655 | var846;
assign var848 = var656 & var754;
assign var849 = var659 & var753;
assign var850 = var658 | var849;
assign var851 = var659 & var754;
assign var852 = var562 & var753;
assign var853 = var561 | var852;
assign var854 = var562 & var754;
assign var855 = var565 & var753;
assign var856 = var564 | var855;
assign var857 = var565 & var754;
assign var858 = var470 & var753;
assign var859 = var469 | var858;
assign var860 = var470 & var754;
assign var861 = var303 & var753;
assign var862 = var302 | var861;
assign var863 = var303 & var754;
assign var864 = var778 & var801;
assign var865 = var777 | var864;
assign var866 = var781 & var801;
assign var867 = var780 | var866;
assign var868 = var784 & var801;
assign var869 = var783 | var868;
assign var870 = var787 & var801;
assign var871 = var786 | var870;
assign var872 = var790 & var801;
assign var873 = var789 | var872;
assign var874 = var793 & var801;
assign var875 = var792 | var874;
assign var876 = var796 & var801;
assign var877 = var795 | var876;
assign var878 = var799 & var801;
assign var879 = var798 | var878;
assign var880 = var698 & var801;
assign var881 = var697 | var880;
assign var882 = var701 & var801;
assign var883 = var700 | var882;
assign var884 = var704 & var801;
assign var885 = var703 | var884;
assign var886 = var707 & var801;
assign var887 = var706 | var886;
assign var888 = var610 & var801;
assign var889 = var609 | var888;
assign var890 = var613 & var801;
assign var891 = var612 | var890;
assign var892 = var518 & var801;
assign var893 = var517 | var892;
assign var894 = var399 & var801;
assign var895 = var398 | var894;
assign var896 = var818 & var865;
assign var897 = var817 | var896;
assign var898 = var821 & var865;
assign var899 = var820 | var898;
assign var900 = var824 & var865;
assign var901 = var823 | var900;
assign var902 = var827 & var865;
assign var903 = var826 | var902;
assign var904 = var830 & var865;
assign var905 = var829 | var904;
assign var906 = var833 & var865;
assign var907 = var832 | var906;
assign var908 = var836 & var865;
assign var909 = var835 | var908;
assign var910 = var839 & var865;
assign var911 = var838 | var910;
assign var912 = var842 & var865;
assign var913 = var841 | var912;
assign var914 = var845 & var865;
assign var915 = var844 | var914;
assign var916 = var848 & var865;
assign var917 = var847 | var916;
assign var918 = var851 & var865;
assign var919 = var850 | var918;
assign var920 = var854 & var865;
assign var921 = var853 | var920;
assign var922 = var857 & var865;
assign var923 = var856 | var922;
assign var924 = var860 & var865;
assign var925 = var859 | var924;
assign var926 = var863 & var865;
assign var927 = var862 | var926;
assign var928 = var754 & var865;
assign var929 = var753 | var928;
assign var930 = var757 & var865;
assign var931 = var756 | var930;
assign var932 = var760 & var865;
assign var933 = var759 | var932;
assign var934 = var763 & var865;
assign var935 = var762 | var934;
assign var936 = var766 & var865;
assign var937 = var765 | var936;
assign var938 = var769 & var865;
assign var939 = var768 | var938;
assign var940 = var772 & var865;
assign var941 = var771 | var940;
assign var942 = var775 & var865;
assign var943 = var774 | var942;
assign var944 = var674 & var865;
assign var945 = var673 | var944;
assign var946 = var677 & var865;
assign var947 = var676 | var946;
assign var948 = var680 & var865;
assign var949 = var679 | var948;
assign var950 = var683 & var865;
assign var951 = var682 | var950;
assign var952 = var586 & var865;
assign var953 = var585 | var952;
assign var954 = var589 & var865;
assign var955 = var588 | var954;
assign var956 = var494 & var865;
assign var957 = var493 | var956;
assign var958 = var351 & var865;
assign var959 = var350 | var958;
assign var960 = var254 & var899;
assign var961 = var126 | var960;
assign var962 = var254 & var821;
assign var963 = var252 & var901;
assign var964 = var124 | var963;
assign var965 = var252 & var824;
assign var966 = var250 & var903;
assign var967 = var122 | var966;
assign var968 = var250 & var827;
assign var969 = var248 & var905;
assign var970 = var120 | var969;
assign var971 = var248 & var830;
assign var972 = var246 & var907;
assign var973 = var118 | var972;
assign var974 = var246 & var833;
assign var975 = var244 & var909;
assign var976 = var116 | var975;
assign var977 = var244 & var836;
assign var978 = var242 & var911;
assign var979 = var114 | var978;
assign var980 = var242 & var839;
assign var981 = var240 & var913;
assign var982 = var112 | var981;
assign var983 = var240 & var842;
assign var984 = var238 & var915;
assign var985 = var110 | var984;
assign var986 = var238 & var845;
assign var987 = var236 & var917;
assign var988 = var108 | var987;
assign var989 = var236 & var848;
assign var990 = var234 & var919;
assign var991 = var106 | var990;
assign var992 = var234 & var851;
assign var993 = var232 & var921;
assign var994 = var104 | var993;
assign var995 = var232 & var854;
assign var996 = var230 & var923;
assign var997 = var102 | var996;
assign var998 = var230 & var857;
assign var999 = var228 & var925;
assign var1000 = var100 | var999;
assign var1001 = var228 & var860;
assign var1002 = var226 & var927;
assign var1003 = var98 | var1002;
assign var1004 = var226 & var863;
assign var1005 = var224 & var929;
assign var1006 = var96 | var1005;
assign var1007 = var224 & var754;
assign var1008 = var222 & var931;
assign var1009 = var94 | var1008;
assign var1010 = var222 & var757;
assign var1011 = var220 & var933;
assign var1012 = var92 | var1011;
assign var1013 = var220 & var760;
assign var1014 = var218 & var935;
assign var1015 = var90 | var1014;
assign var1016 = var218 & var763;
assign var1017 = var216 & var937;
assign var1018 = var88 | var1017;
assign var1019 = var216 & var766;
assign var1020 = var214 & var939;
assign var1021 = var86 | var1020;
assign var1022 = var214 & var769;
assign var1023 = var212 & var941;
assign var1024 = var84 | var1023;
assign var1025 = var212 & var772;
assign var1026 = var210 & var943;
assign var1027 = var82 | var1026;
assign var1028 = var210 & var775;
assign var1029 = var208 & var945;
assign var1030 = var80 | var1029;
assign var1031 = var208 & var674;
assign var1032 = var206 & var947;
assign var1033 = var78 | var1032;
assign var1034 = var206 & var677;
assign var1035 = var204 & var949;
assign var1036 = var76 | var1035;
assign var1037 = var204 & var680;
assign var1038 = var202 & var951;
assign var1039 = var74 | var1038;
assign var1040 = var202 & var683;
assign var1041 = var200 & var953;
assign var1042 = var72 | var1041;
assign var1043 = var200 & var586;
assign var1044 = var198 & var955;
assign var1045 = var70 | var1044;
assign var1046 = var198 & var589;
assign var1047 = var196 & var957;
assign var1048 = var68 | var1047;
assign var1049 = var196 & var494;
assign var1050 = var194 & var959;
assign var1051 = var66 | var1050;
assign var1052 = var194 & var351;
assign var1053 = var192 & var865;
assign var1054 = var64 | var1053;
assign var1055 = var192 & var778;
assign var1056 = var190 & var867;
assign var1057 = var62 | var1056;
assign var1058 = var190 & var781;
assign var1059 = var188 & var869;
assign var1060 = var60 | var1059;
assign var1061 = var188 & var784;
assign var1062 = var186 & var871;
assign var1063 = var58 | var1062;
assign var1064 = var186 & var787;
assign var1065 = var184 & var873;
assign var1066 = var56 | var1065;
assign var1067 = var184 & var790;
assign var1068 = var182 & var875;
assign var1069 = var54 | var1068;
assign var1070 = var182 & var793;
assign var1071 = var180 & var877;
assign var1072 = var52 | var1071;
assign var1073 = var180 & var796;
assign var1074 = var178 & var879;
assign var1075 = var50 | var1074;
assign var1076 = var178 & var799;
assign var1077 = var176 & var881;
assign var1078 = var48 | var1077;
assign var1079 = var176 & var698;
assign var1080 = var174 & var883;
assign var1081 = var46 | var1080;
assign var1082 = var174 & var701;
assign var1083 = var172 & var885;
assign var1084 = var44 | var1083;
assign var1085 = var172 & var704;
assign var1086 = var170 & var887;
assign var1087 = var42 | var1086;
assign var1088 = var170 & var707;
assign var1089 = var168 & var889;
assign var1090 = var40 | var1089;
assign var1091 = var168 & var610;
assign var1092 = var166 & var891;
assign var1093 = var38 | var1092;
assign var1094 = var166 & var613;
assign var1095 = var164 & var893;
assign var1096 = var36 | var1095;
assign var1097 = var164 & var518;
assign var1098 = var162 & var895;
assign var1099 = var34 | var1098;
assign var1100 = var162 & var399;
assign var1101 = var160 & var801;
assign var1102 = var32 | var1101;
assign var1103 = var160 & var710;
assign var1104 = var158 & var803;
assign var1105 = var30 | var1104;
assign var1106 = var158 & var713;
assign var1107 = var156 & var805;
assign var1108 = var28 | var1107;
assign var1109 = var156 & var716;
assign var1110 = var154 & var807;
assign var1111 = var26 | var1110;
assign var1112 = var154 & var719;
assign var1113 = var152 & var809;
assign var1114 = var24 | var1113;
assign var1115 = var152 & var622;
assign var1116 = var150 & var811;
assign var1117 = var22 | var1116;
assign var1118 = var150 & var625;
assign var1119 = var148 & var813;
assign var1120 = var20 | var1119;
assign var1121 = var148 & var530;
assign var1122 = var146 & var815;
assign var1123 = var18 | var1122;
assign var1124 = var146 & var423;
assign var1125 = var144 & var721;
assign var1126 = var16 | var1125;
assign var1127 = var144 & var628;
assign var1128 = var142 & var723;
assign var1129 = var14 | var1128;
assign var1130 = var142 & var631;
assign var1131 = var140 & var725;
assign var1132 = var12 | var1131;
assign var1133 = var140 & var536;
assign var1134 = var138 & var727;
assign var1135 = var10 | var1134;
assign var1136 = var138 & var435;
assign var1137 = var136 & var633;
assign var1138 = var8 | var1137;
assign var1139 = var136 & var539;
assign var1140 = var134 & var635;
assign var1141 = var6 | var1140;
assign var1142 = var134 & var441;
assign var1143 = var132 & var541;
assign var1144 = var4 | var1143;
assign var1145 = var132 & var444;
assign var1146 = var130 & var446;
assign var1147 = var2 | var1146;
assign var1148 = var130 & var129;
assign var1149 = var129 ^ var0;
assign var1150 = var130 ^ var446;
assign var1151 = var131 ^ var1147;
assign var1152 = var132 ^ var541;
assign var1153 = var133 ^ var1144;
assign var1154 = var134 ^ var635;
assign var1155 = var135 ^ var1141;
assign var1156 = var136 ^ var633;
assign var1157 = var137 ^ var1138;
assign var1158 = var138 ^ var727;
assign var1159 = var139 ^ var1135;
assign var1160 = var140 ^ var725;
assign var1161 = var141 ^ var1132;
assign var1162 = var142 ^ var723;
assign var1163 = var143 ^ var1129;
assign var1164 = var144 ^ var721;
assign var1165 = var145 ^ var1126;
assign var1166 = var146 ^ var815;
assign var1167 = var147 ^ var1123;
assign var1168 = var148 ^ var813;
assign var1169 = var149 ^ var1120;
assign var1170 = var150 ^ var811;
assign var1171 = var151 ^ var1117;
assign var1172 = var152 ^ var809;
assign var1173 = var153 ^ var1114;
assign var1174 = var154 ^ var807;
assign var1175 = var155 ^ var1111;
assign var1176 = var156 ^ var805;
assign var1177 = var157 ^ var1108;
assign var1178 = var158 ^ var803;
assign var1179 = var159 ^ var1105;
assign var1180 = var160 ^ var801;
assign var1181 = var161 ^ var1102;
assign var1182 = var162 ^ var895;
assign var1183 = var163 ^ var1099;
assign var1184 = var164 ^ var893;
assign var1185 = var165 ^ var1096;
assign var1186 = var166 ^ var891;
assign var1187 = var167 ^ var1093;
assign var1188 = var168 ^ var889;
assign var1189 = var169 ^ var1090;
assign var1190 = var170 ^ var887;
assign var1191 = var171 ^ var1087;
assign var1192 = var172 ^ var885;
assign var1193 = var173 ^ var1084;
assign var1194 = var174 ^ var883;
assign var1195 = var175 ^ var1081;
assign var1196 = var176 ^ var881;
assign var1197 = var177 ^ var1078;
assign var1198 = var178 ^ var879;
assign var1199 = var179 ^ var1075;
assign var1200 = var180 ^ var877;
assign var1201 = var181 ^ var1072;
assign var1202 = var182 ^ var875;
assign var1203 = var183 ^ var1069;
assign var1204 = var184 ^ var873;
assign var1205 = var185 ^ var1066;
assign var1206 = var186 ^ var871;
assign var1207 = var187 ^ var1063;
assign var1208 = var188 ^ var869;
assign var1209 = var189 ^ var1060;
assign var1210 = var190 ^ var867;
assign var1211 = var191 ^ var1057;
assign var1212 = var192 ^ var865;
assign var1213 = var193 ^ var1054;
assign var1214 = var194 ^ var959;
assign var1215 = var195 ^ var1051;
assign var1216 = var196 ^ var957;
assign var1217 = var197 ^ var1048;
assign var1218 = var198 ^ var955;
assign var1219 = var199 ^ var1045;
assign var1220 = var200 ^ var953;
assign var1221 = var201 ^ var1042;
assign var1222 = var202 ^ var951;
assign var1223 = var203 ^ var1039;
assign var1224 = var204 ^ var949;
assign var1225 = var205 ^ var1036;
assign var1226 = var206 ^ var947;
assign var1227 = var207 ^ var1033;
assign var1228 = var208 ^ var945;
assign var1229 = var209 ^ var1030;
assign var1230 = var210 ^ var943;
assign var1231 = var211 ^ var1027;
assign var1232 = var212 ^ var941;
assign var1233 = var213 ^ var1024;
assign var1234 = var214 ^ var939;
assign var1235 = var215 ^ var1021;
assign var1236 = var216 ^ var937;
assign var1237 = var217 ^ var1018;
assign var1238 = var218 ^ var935;
assign var1239 = var219 ^ var1015;
assign var1240 = var220 ^ var933;
assign var1241 = var221 ^ var1012;
assign var1242 = var222 ^ var931;
assign var1243 = var223 ^ var1009;
assign var1244 = var224 ^ var929;
assign var1245 = var225 ^ var1006;
assign var1246 = var226 ^ var927;
assign var1247 = var227 ^ var1003;
assign var1248 = var228 ^ var925;
assign var1249 = var229 ^ var1000;
assign var1250 = var230 ^ var923;
assign var1251 = var231 ^ var997;
assign var1252 = var232 ^ var921;
assign var1253 = var233 ^ var994;
assign var1254 = var234 ^ var919;
assign var1255 = var235 ^ var991;
assign var1256 = var236 ^ var917;
assign var1257 = var237 ^ var988;
assign var1258 = var238 ^ var915;
assign var1259 = var239 ^ var985;
assign var1260 = var240 ^ var913;
assign var1261 = var241 ^ var982;
assign var1262 = var242 ^ var911;
assign var1263 = var243 ^ var979;
assign var1264 = var244 ^ var909;
assign var1265 = var245 ^ var976;
assign var1266 = var246 ^ var907;
assign var1267 = var247 ^ var973;
assign var1268 = var248 ^ var905;
assign var1269 = var249 ^ var970;
assign var1270 = var250 ^ var903;
assign var1271 = var251 ^ var967;
assign var1272 = var252 ^ var901;
assign var1273 = var253 ^ var964;
assign var1274 = var254 ^ var899;
assign var1275 = var255 ^ var961;
assign out0 = var897;
assign out1 = var1275;
assign out2 = var1274;
assign out3 = var1273;
assign out4 = var1272;
assign out5 = var1271;
assign out6 = var1270;
assign out7 = var1269;
assign out8 = var1268;
assign out9 = var1267;
assign out10 = var1266;
assign out11 = var1265;
assign out12 = var1264;
assign out13 = var1263;
assign out14 = var1262;
assign out15 = var1261;
assign out16 = var1260;
assign out17 = var1259;
assign out18 = var1258;
assign out19 = var1257;
assign out20 = var1256;
assign out21 = var1255;
assign out22 = var1254;
assign out23 = var1253;
assign out24 = var1252;
assign out25 = var1251;
assign out26 = var1250;
assign out27 = var1249;
assign out28 = var1248;
assign out29 = var1247;
assign out30 = var1246;
assign out31 = var1245;
assign out32 = var1244;
assign out33 = var1243;
assign out34 = var1242;
assign out35 = var1241;
assign out36 = var1240;
assign out37 = var1239;
assign out38 = var1238;
assign out39 = var1237;
assign out40 = var1236;
assign out41 = var1235;
assign out42 = var1234;
assign out43 = var1233;
assign out44 = var1232;
assign out45 = var1231;
assign out46 = var1230;
assign out47 = var1229;
assign out48 = var1228;
assign out49 = var1227;
assign out50 = var1226;
assign out51 = var1225;
assign out52 = var1224;
assign out53 = var1223;
assign out54 = var1222;
assign out55 = var1221;
assign out56 = var1220;
assign out57 = var1219;
assign out58 = var1218;
assign out59 = var1217;
assign out60 = var1216;
assign out61 = var1215;
assign out62 = var1214;
assign out63 = var1213;
assign out64 = var1212;
assign out65 = var1211;
assign out66 = var1210;
assign out67 = var1209;
assign out68 = var1208;
assign out69 = var1207;
assign out70 = var1206;
assign out71 = var1205;
assign out72 = var1204;
assign out73 = var1203;
assign out74 = var1202;
assign out75 = var1201;
assign out76 = var1200;
assign out77 = var1199;
assign out78 = var1198;
assign out79 = var1197;
assign out80 = var1196;
assign out81 = var1195;
assign out82 = var1194;
assign out83 = var1193;
assign out84 = var1192;
assign out85 = var1191;
assign out86 = var1190;
assign out87 = var1189;
assign out88 = var1188;
assign out89 = var1187;
assign out90 = var1186;
assign out91 = var1185;
assign out92 = var1184;
assign out93 = var1183;
assign out94 = var1182;
assign out95 = var1181;
assign out96 = var1180;
assign out97 = var1179;
assign out98 = var1178;
assign out99 = var1177;
assign out100 = var1176;
assign out101 = var1175;
assign out102 = var1174;
assign out103 = var1173;
assign out104 = var1172;
assign out105 = var1171;
assign out106 = var1170;
assign out107 = var1169;
assign out108 = var1168;
assign out109 = var1167;
assign out110 = var1166;
assign out111 = var1165;
assign out112 = var1164;
assign out113 = var1163;
assign out114 = var1162;
assign out115 = var1161;
assign out116 = var1160;
assign out117 = var1159;
assign out118 = var1158;
assign out119 = var1157;
assign out120 = var1156;
assign out121 = var1155;
assign out122 = var1154;
assign out123 = var1153;
assign out124 = var1152;
assign out125 = var1151;
assign out126 = var1150;
assign out127 = var1149;
assign out128 = var128;
endmodule 
