module bk8 (in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, out0, out1, out2, out3, out4, out5, out6, out7, out8, );
input in0;
input in1;
input in2;
input in3;
input in4;
input in5;
input in6;
input in7;
input in8;
input in9;
input in10;
input in11;
input in12;
input in13;
input in14;
input in15;
output out0;
output out1;
output out2;
output out3;
output out4;
output out5;
output out6;
output out7;
output out8;
wire var0;
wire var1;
wire var2;
wire var3;
wire var4;
wire var5;
wire var6;
wire var7;
wire var8;
wire var9;
wire var10;
wire var11;
wire var12;
wire var13;
wire var14;
wire var15;
wire var16;
wire var17;
wire var18;
wire var19;
wire var20;
wire var21;
wire var22;
wire var23;
wire var24;
wire var25;
wire var26;
wire var27;
wire var28;
wire var29;
wire var30;
wire var31;
wire var32;
wire var33;
wire var34;
wire var35;
wire var36;
wire var37;
wire var38;
wire var39;
wire var40;
wire var41;
wire var42;
wire var43;
wire var44;
wire var45;
wire var46;
wire var47;
wire var48;
wire var49;
wire var50;
wire var51;
assign var0 = in15 & in7;
assign var1 = in14 & in6;
assign var2 = in13 & in5;
assign var3 = in12 & in4;
assign var4 = in11 & in3;
assign var5 = in10 & in2;
assign var6 = in9 & in1;
assign var7 = in8 & in0;
assign var8 = in15 ^ in7;
assign var9 = in14 ^ in6;
assign var10 = in13 ^ in5;
assign var11 = in12 ^ in4;
assign var12 = in11 ^ in3;
assign var13 = in10 ^ in2;
assign var14 = in9 ^ in1;
assign var15 = in8 ^ in0;
assign var16 = var15 & var6;
assign var17 = var7 | var16;
assign var18 = var15 & var14;
assign var19 = var13 & var4;
assign var20 = var5 | var19;
assign var21 = var13 & var12;
assign var22 = var11 & var2;
assign var23 = var3 | var22;
assign var24 = var11 & var10;
assign var25 = var9 & var0;
assign var26 = var1 | var25;
assign var27 = var18 & var20;
assign var28 = var17 | var27;
assign var29 = var18 & var21;
assign var30 = var24 & var26;
assign var31 = var23 | var30;
assign var32 = var29 & var31;
assign var33 = var28 | var32;
assign var34 = var21 & var31;
assign var35 = var20 | var34;
assign var36 = var14 & var35;
assign var37 = var6 | var36;
assign var38 = var14 & var21;
assign var39 = var12 & var31;
assign var40 = var4 | var39;
assign var41 = var12 & var24;
assign var42 = var10 & var26;
assign var43 = var2 | var42;
assign var44 = var10 & var9;
assign var45 = var9 ^ var0;
assign var46 = var10 ^ var26;
assign var47 = var11 ^ var43;
assign var48 = var12 ^ var31;
assign var49 = var13 ^ var40;
assign var50 = var14 ^ var35;
assign var51 = var15 ^ var37;
assign out0 = var33;
assign out1 = var51;
assign out2 = var50;
assign out3 = var49;
assign out4 = var48;
assign out5 = var47;
assign out6 = var46;
assign out7 = var45;
assign out8 = var8;
endmodule 
