module ks16 (in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, );
input in0;
input in1;
input in2;
input in3;
input in4;
input in5;
input in6;
input in7;
input in8;
input in9;
input in10;
input in11;
input in12;
input in13;
input in14;
input in15;
input in16;
input in17;
input in18;
input in19;
input in20;
input in21;
input in22;
input in23;
input in24;
input in25;
input in26;
input in27;
input in28;
input in29;
input in30;
input in31;
output out0;
output out1;
output out2;
output out3;
output out4;
output out5;
output out6;
output out7;
output out8;
output out9;
output out10;
output out11;
output out12;
output out13;
output out14;
output out15;
output out16;
wire var0;
wire var1;
wire var2;
wire var3;
wire var4;
wire var5;
wire var6;
wire var7;
wire var8;
wire var9;
wire var10;
wire var11;
wire var12;
wire var13;
wire var14;
wire var15;
wire var16;
wire var17;
wire var18;
wire var19;
wire var20;
wire var21;
wire var22;
wire var23;
wire var24;
wire var25;
wire var26;
wire var27;
wire var28;
wire var29;
wire var30;
wire var31;
wire var32;
wire var33;
wire var34;
wire var35;
wire var36;
wire var37;
wire var38;
wire var39;
wire var40;
wire var41;
wire var42;
wire var43;
wire var44;
wire var45;
wire var46;
wire var47;
wire var48;
wire var49;
wire var50;
wire var51;
wire var52;
wire var53;
wire var54;
wire var55;
wire var56;
wire var57;
wire var58;
wire var59;
wire var60;
wire var61;
wire var62;
wire var63;
wire var64;
wire var65;
wire var66;
wire var67;
wire var68;
wire var69;
wire var70;
wire var71;
wire var72;
wire var73;
wire var74;
wire var75;
wire var76;
wire var77;
wire var78;
wire var79;
wire var80;
wire var81;
wire var82;
wire var83;
wire var84;
wire var85;
wire var86;
wire var87;
wire var88;
wire var89;
wire var90;
wire var91;
wire var92;
wire var93;
wire var94;
wire var95;
wire var96;
wire var97;
wire var98;
wire var99;
wire var100;
wire var101;
wire var102;
wire var103;
wire var104;
wire var105;
wire var106;
wire var107;
wire var108;
wire var109;
wire var110;
wire var111;
wire var112;
wire var113;
wire var114;
wire var115;
wire var116;
wire var117;
wire var118;
wire var119;
wire var120;
wire var121;
wire var122;
wire var123;
wire var124;
wire var125;
wire var126;
wire var127;
wire var128;
wire var129;
wire var130;
wire var131;
wire var132;
wire var133;
wire var134;
wire var135;
wire var136;
wire var137;
wire var138;
wire var139;
wire var140;
wire var141;
wire var142;
wire var143;
wire var144;
wire var145;
wire var146;
wire var147;
wire var148;
wire var149;
wire var150;
wire var151;
wire var152;
wire var153;
wire var154;
wire var155;
wire var156;
wire var157;
wire var158;
wire var159;
wire var160;
wire var161;
wire var162;
wire var163;
wire var164;
wire var165;
wire var166;
wire var167;
wire var168;
wire var169;
wire var170;
wire var171;
wire var172;
wire var173;
wire var174;
wire var175;
wire var176;
wire var177;
wire var178;
assign var0 = in31 & in15;
assign var1 = in30 & in14;
assign var2 = in29 & in13;
assign var3 = in28 & in12;
assign var4 = in27 & in11;
assign var5 = in26 & in10;
assign var6 = in25 & in9;
assign var7 = in24 & in8;
assign var8 = in23 & in7;
assign var9 = in22 & in6;
assign var10 = in21 & in5;
assign var11 = in20 & in4;
assign var12 = in19 & in3;
assign var13 = in18 & in2;
assign var14 = in17 & in1;
assign var15 = in16 & in0;
assign var16 = in31 ^ in15;
assign var17 = in30 ^ in14;
assign var18 = in29 ^ in13;
assign var19 = in28 ^ in12;
assign var20 = in27 ^ in11;
assign var21 = in26 ^ in10;
assign var22 = in25 ^ in9;
assign var23 = in24 ^ in8;
assign var24 = in23 ^ in7;
assign var25 = in22 ^ in6;
assign var26 = in21 ^ in5;
assign var27 = in20 ^ in4;
assign var28 = in19 ^ in3;
assign var29 = in18 ^ in2;
assign var30 = in17 ^ in1;
assign var31 = in16 ^ in0;
assign var32 = var31 & var14;
assign var33 = var15 | var32;
assign var34 = var31 & var30;
assign var35 = var30 & var13;
assign var36 = var14 | var35;
assign var37 = var30 & var29;
assign var38 = var29 & var12;
assign var39 = var13 | var38;
assign var40 = var29 & var28;
assign var41 = var28 & var11;
assign var42 = var12 | var41;
assign var43 = var28 & var27;
assign var44 = var27 & var10;
assign var45 = var11 | var44;
assign var46 = var27 & var26;
assign var47 = var26 & var9;
assign var48 = var10 | var47;
assign var49 = var26 & var25;
assign var50 = var25 & var8;
assign var51 = var9 | var50;
assign var52 = var25 & var24;
assign var53 = var24 & var7;
assign var54 = var8 | var53;
assign var55 = var24 & var23;
assign var56 = var23 & var6;
assign var57 = var7 | var56;
assign var58 = var23 & var22;
assign var59 = var22 & var5;
assign var60 = var6 | var59;
assign var61 = var22 & var21;
assign var62 = var21 & var4;
assign var63 = var5 | var62;
assign var64 = var21 & var20;
assign var65 = var20 & var3;
assign var66 = var4 | var65;
assign var67 = var20 & var19;
assign var68 = var19 & var2;
assign var69 = var3 | var68;
assign var70 = var19 & var18;
assign var71 = var18 & var1;
assign var72 = var2 | var71;
assign var73 = var18 & var17;
assign var74 = var17 & var0;
assign var75 = var1 | var74;
assign var76 = var34 & var39;
assign var77 = var33 | var76;
assign var78 = var34 & var40;
assign var79 = var37 & var42;
assign var80 = var36 | var79;
assign var81 = var37 & var43;
assign var82 = var40 & var45;
assign var83 = var39 | var82;
assign var84 = var40 & var46;
assign var85 = var43 & var48;
assign var86 = var42 | var85;
assign var87 = var43 & var49;
assign var88 = var46 & var51;
assign var89 = var45 | var88;
assign var90 = var46 & var52;
assign var91 = var49 & var54;
assign var92 = var48 | var91;
assign var93 = var49 & var55;
assign var94 = var52 & var57;
assign var95 = var51 | var94;
assign var96 = var52 & var58;
assign var97 = var55 & var60;
assign var98 = var54 | var97;
assign var99 = var55 & var61;
assign var100 = var58 & var63;
assign var101 = var57 | var100;
assign var102 = var58 & var64;
assign var103 = var61 & var66;
assign var104 = var60 | var103;
assign var105 = var61 & var67;
assign var106 = var64 & var69;
assign var107 = var63 | var106;
assign var108 = var64 & var70;
assign var109 = var67 & var72;
assign var110 = var66 | var109;
assign var111 = var67 & var73;
assign var112 = var70 & var75;
assign var113 = var69 | var112;
assign var114 = var73 & var0;
assign var115 = var72 | var114;
assign var116 = var78 & var89;
assign var117 = var77 | var116;
assign var118 = var78 & var90;
assign var119 = var81 & var92;
assign var120 = var80 | var119;
assign var121 = var81 & var93;
assign var122 = var84 & var95;
assign var123 = var83 | var122;
assign var124 = var84 & var96;
assign var125 = var87 & var98;
assign var126 = var86 | var125;
assign var127 = var87 & var99;
assign var128 = var90 & var101;
assign var129 = var89 | var128;
assign var130 = var90 & var102;
assign var131 = var93 & var104;
assign var132 = var92 | var131;
assign var133 = var93 & var105;
assign var134 = var96 & var107;
assign var135 = var95 | var134;
assign var136 = var96 & var108;
assign var137 = var99 & var110;
assign var138 = var98 | var137;
assign var139 = var99 & var111;
assign var140 = var102 & var113;
assign var141 = var101 | var140;
assign var142 = var105 & var115;
assign var143 = var104 | var142;
assign var144 = var108 & var75;
assign var145 = var107 | var144;
assign var146 = var111 & var0;
assign var147 = var110 | var146;
assign var148 = var118 & var141;
assign var149 = var117 | var148;
assign var150 = var121 & var143;
assign var151 = var120 | var150;
assign var152 = var124 & var145;
assign var153 = var123 | var152;
assign var154 = var127 & var147;
assign var155 = var126 | var154;
assign var156 = var130 & var113;
assign var157 = var129 | var156;
assign var158 = var133 & var115;
assign var159 = var132 | var158;
assign var160 = var136 & var75;
assign var161 = var135 | var160;
assign var162 = var139 & var0;
assign var163 = var138 | var162;
assign var164 = var17 ^ var0;
assign var165 = var18 ^ var75;
assign var166 = var19 ^ var115;
assign var167 = var20 ^ var113;
assign var168 = var21 ^ var147;
assign var169 = var22 ^ var145;
assign var170 = var23 ^ var143;
assign var171 = var24 ^ var141;
assign var172 = var25 ^ var163;
assign var173 = var26 ^ var161;
assign var174 = var27 ^ var159;
assign var175 = var28 ^ var157;
assign var176 = var29 ^ var155;
assign var177 = var30 ^ var153;
assign var178 = var31 ^ var151;
assign out0 = var149;
assign out1 = var178;
assign out2 = var177;
assign out3 = var176;
assign out4 = var175;
assign out5 = var174;
assign out6 = var173;
assign out7 = var172;
assign out8 = var171;
assign out9 = var170;
assign out10 = var169;
assign out11 = var168;
assign out12 = var167;
assign out13 = var166;
assign out14 = var165;
assign out15 = var164;
assign out16 = var16;
endmodule 
