module kn128 (in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, in100, in101, in102, in103, in104, in105, in106, in107, in108, in109, in110, in111, in112, in113, in114, in115, in116, in117, in118, in119, in120, in121, in122, in123, in124, in125, in126, in127, in128, in129, in130, in131, in132, in133, in134, in135, in136, in137, in138, in139, in140, in141, in142, in143, in144, in145, in146, in147, in148, in149, in150, in151, in152, in153, in154, in155, in156, in157, in158, in159, in160, in161, in162, in163, in164, in165, in166, in167, in168, in169, in170, in171, in172, in173, in174, in175, in176, in177, in178, in179, in180, in181, in182, in183, in184, in185, in186, in187, in188, in189, in190, in191, in192, in193, in194, in195, in196, in197, in198, in199, in200, in201, in202, in203, in204, in205, in206, in207, in208, in209, in210, in211, in212, in213, in214, in215, in216, in217, in218, in219, in220, in221, in222, in223, in224, in225, in226, in227, in228, in229, in230, in231, in232, in233, in234, in235, in236, in237, in238, in239, in240, in241, in242, in243, in244, in245, in246, in247, in248, in249, in250, in251, in252, in253, in254, in255, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, out30, out31, out32, out33, out34, out35, out36, out37, out38, out39, out40, out41, out42, out43, out44, out45, out46, out47, out48, out49, out50, out51, out52, out53, out54, out55, out56, out57, out58, out59, out60, out61, out62, out63, out64, out65, out66, out67, out68, out69, out70, out71, out72, out73, out74, out75, out76, out77, out78, out79, out80, out81, out82, out83, out84, out85, out86, out87, out88, out89, out90, out91, out92, out93, out94, out95, out96, out97, out98, out99, out100, out101, out102, out103, out104, out105, out106, out107, out108, out109, out110, out111, out112, out113, out114, out115, out116, out117, out118, out119, out120, out121, out122, out123, out124, out125, out126, out127, out128, );
input in0;
input in1;
input in2;
input in3;
input in4;
input in5;
input in6;
input in7;
input in8;
input in9;
input in10;
input in11;
input in12;
input in13;
input in14;
input in15;
input in16;
input in17;
input in18;
input in19;
input in20;
input in21;
input in22;
input in23;
input in24;
input in25;
input in26;
input in27;
input in28;
input in29;
input in30;
input in31;
input in32;
input in33;
input in34;
input in35;
input in36;
input in37;
input in38;
input in39;
input in40;
input in41;
input in42;
input in43;
input in44;
input in45;
input in46;
input in47;
input in48;
input in49;
input in50;
input in51;
input in52;
input in53;
input in54;
input in55;
input in56;
input in57;
input in58;
input in59;
input in60;
input in61;
input in62;
input in63;
input in64;
input in65;
input in66;
input in67;
input in68;
input in69;
input in70;
input in71;
input in72;
input in73;
input in74;
input in75;
input in76;
input in77;
input in78;
input in79;
input in80;
input in81;
input in82;
input in83;
input in84;
input in85;
input in86;
input in87;
input in88;
input in89;
input in90;
input in91;
input in92;
input in93;
input in94;
input in95;
input in96;
input in97;
input in98;
input in99;
input in100;
input in101;
input in102;
input in103;
input in104;
input in105;
input in106;
input in107;
input in108;
input in109;
input in110;
input in111;
input in112;
input in113;
input in114;
input in115;
input in116;
input in117;
input in118;
input in119;
input in120;
input in121;
input in122;
input in123;
input in124;
input in125;
input in126;
input in127;
input in128;
input in129;
input in130;
input in131;
input in132;
input in133;
input in134;
input in135;
input in136;
input in137;
input in138;
input in139;
input in140;
input in141;
input in142;
input in143;
input in144;
input in145;
input in146;
input in147;
input in148;
input in149;
input in150;
input in151;
input in152;
input in153;
input in154;
input in155;
input in156;
input in157;
input in158;
input in159;
input in160;
input in161;
input in162;
input in163;
input in164;
input in165;
input in166;
input in167;
input in168;
input in169;
input in170;
input in171;
input in172;
input in173;
input in174;
input in175;
input in176;
input in177;
input in178;
input in179;
input in180;
input in181;
input in182;
input in183;
input in184;
input in185;
input in186;
input in187;
input in188;
input in189;
input in190;
input in191;
input in192;
input in193;
input in194;
input in195;
input in196;
input in197;
input in198;
input in199;
input in200;
input in201;
input in202;
input in203;
input in204;
input in205;
input in206;
input in207;
input in208;
input in209;
input in210;
input in211;
input in212;
input in213;
input in214;
input in215;
input in216;
input in217;
input in218;
input in219;
input in220;
input in221;
input in222;
input in223;
input in224;
input in225;
input in226;
input in227;
input in228;
input in229;
input in230;
input in231;
input in232;
input in233;
input in234;
input in235;
input in236;
input in237;
input in238;
input in239;
input in240;
input in241;
input in242;
input in243;
input in244;
input in245;
input in246;
input in247;
input in248;
input in249;
input in250;
input in251;
input in252;
input in253;
input in254;
input in255;
output out0;
output out1;
output out2;
output out3;
output out4;
output out5;
output out6;
output out7;
output out8;
output out9;
output out10;
output out11;
output out12;
output out13;
output out14;
output out15;
output out16;
output out17;
output out18;
output out19;
output out20;
output out21;
output out22;
output out23;
output out24;
output out25;
output out26;
output out27;
output out28;
output out29;
output out30;
output out31;
output out32;
output out33;
output out34;
output out35;
output out36;
output out37;
output out38;
output out39;
output out40;
output out41;
output out42;
output out43;
output out44;
output out45;
output out46;
output out47;
output out48;
output out49;
output out50;
output out51;
output out52;
output out53;
output out54;
output out55;
output out56;
output out57;
output out58;
output out59;
output out60;
output out61;
output out62;
output out63;
output out64;
output out65;
output out66;
output out67;
output out68;
output out69;
output out70;
output out71;
output out72;
output out73;
output out74;
output out75;
output out76;
output out77;
output out78;
output out79;
output out80;
output out81;
output out82;
output out83;
output out84;
output out85;
output out86;
output out87;
output out88;
output out89;
output out90;
output out91;
output out92;
output out93;
output out94;
output out95;
output out96;
output out97;
output out98;
output out99;
output out100;
output out101;
output out102;
output out103;
output out104;
output out105;
output out106;
output out107;
output out108;
output out109;
output out110;
output out111;
output out112;
output out113;
output out114;
output out115;
output out116;
output out117;
output out118;
output out119;
output out120;
output out121;
output out122;
output out123;
output out124;
output out125;
output out126;
output out127;
output out128;
wire var0;
wire var1;
wire var2;
wire var3;
wire var4;
wire var5;
wire var6;
wire var7;
wire var8;
wire var9;
wire var10;
wire var11;
wire var12;
wire var13;
wire var14;
wire var15;
wire var16;
wire var17;
wire var18;
wire var19;
wire var20;
wire var21;
wire var22;
wire var23;
wire var24;
wire var25;
wire var26;
wire var27;
wire var28;
wire var29;
wire var30;
wire var31;
wire var32;
wire var33;
wire var34;
wire var35;
wire var36;
wire var37;
wire var38;
wire var39;
wire var40;
wire var41;
wire var42;
wire var43;
wire var44;
wire var45;
wire var46;
wire var47;
wire var48;
wire var49;
wire var50;
wire var51;
wire var52;
wire var53;
wire var54;
wire var55;
wire var56;
wire var57;
wire var58;
wire var59;
wire var60;
wire var61;
wire var62;
wire var63;
wire var64;
wire var65;
wire var66;
wire var67;
wire var68;
wire var69;
wire var70;
wire var71;
wire var72;
wire var73;
wire var74;
wire var75;
wire var76;
wire var77;
wire var78;
wire var79;
wire var80;
wire var81;
wire var82;
wire var83;
wire var84;
wire var85;
wire var86;
wire var87;
wire var88;
wire var89;
wire var90;
wire var91;
wire var92;
wire var93;
wire var94;
wire var95;
wire var96;
wire var97;
wire var98;
wire var99;
wire var100;
wire var101;
wire var102;
wire var103;
wire var104;
wire var105;
wire var106;
wire var107;
wire var108;
wire var109;
wire var110;
wire var111;
wire var112;
wire var113;
wire var114;
wire var115;
wire var116;
wire var117;
wire var118;
wire var119;
wire var120;
wire var121;
wire var122;
wire var123;
wire var124;
wire var125;
wire var126;
wire var127;
wire var128;
wire var129;
wire var130;
wire var131;
wire var132;
wire var133;
wire var134;
wire var135;
wire var136;
wire var137;
wire var138;
wire var139;
wire var140;
wire var141;
wire var142;
wire var143;
wire var144;
wire var145;
wire var146;
wire var147;
wire var148;
wire var149;
wire var150;
wire var151;
wire var152;
wire var153;
wire var154;
wire var155;
wire var156;
wire var157;
wire var158;
wire var159;
wire var160;
wire var161;
wire var162;
wire var163;
wire var164;
wire var165;
wire var166;
wire var167;
wire var168;
wire var169;
wire var170;
wire var171;
wire var172;
wire var173;
wire var174;
wire var175;
wire var176;
wire var177;
wire var178;
wire var179;
wire var180;
wire var181;
wire var182;
wire var183;
wire var184;
wire var185;
wire var186;
wire var187;
wire var188;
wire var189;
wire var190;
wire var191;
wire var192;
wire var193;
wire var194;
wire var195;
wire var196;
wire var197;
wire var198;
wire var199;
wire var200;
wire var201;
wire var202;
wire var203;
wire var204;
wire var205;
wire var206;
wire var207;
wire var208;
wire var209;
wire var210;
wire var211;
wire var212;
wire var213;
wire var214;
wire var215;
wire var216;
wire var217;
wire var218;
wire var219;
wire var220;
wire var221;
wire var222;
wire var223;
wire var224;
wire var225;
wire var226;
wire var227;
wire var228;
wire var229;
wire var230;
wire var231;
wire var232;
wire var233;
wire var234;
wire var235;
wire var236;
wire var237;
wire var238;
wire var239;
wire var240;
wire var241;
wire var242;
wire var243;
wire var244;
wire var245;
wire var246;
wire var247;
wire var248;
wire var249;
wire var250;
wire var251;
wire var252;
wire var253;
wire var254;
wire var255;
wire var256;
wire var257;
wire var258;
wire var259;
wire var260;
wire var261;
wire var262;
wire var263;
wire var264;
wire var265;
wire var266;
wire var267;
wire var268;
wire var269;
wire var270;
wire var271;
wire var272;
wire var273;
wire var274;
wire var275;
wire var276;
wire var277;
wire var278;
wire var279;
wire var280;
wire var281;
wire var282;
wire var283;
wire var284;
wire var285;
wire var286;
wire var287;
wire var288;
wire var289;
wire var290;
wire var291;
wire var292;
wire var293;
wire var294;
wire var295;
wire var296;
wire var297;
wire var298;
wire var299;
wire var300;
wire var301;
wire var302;
wire var303;
wire var304;
wire var305;
wire var306;
wire var307;
wire var308;
wire var309;
wire var310;
wire var311;
wire var312;
wire var313;
wire var314;
wire var315;
wire var316;
wire var317;
wire var318;
wire var319;
wire var320;
wire var321;
wire var322;
wire var323;
wire var324;
wire var325;
wire var326;
wire var327;
wire var328;
wire var329;
wire var330;
wire var331;
wire var332;
wire var333;
wire var334;
wire var335;
wire var336;
wire var337;
wire var338;
wire var339;
wire var340;
wire var341;
wire var342;
wire var343;
wire var344;
wire var345;
wire var346;
wire var347;
wire var348;
wire var349;
wire var350;
wire var351;
wire var352;
wire var353;
wire var354;
wire var355;
wire var356;
wire var357;
wire var358;
wire var359;
wire var360;
wire var361;
wire var362;
wire var363;
wire var364;
wire var365;
wire var366;
wire var367;
wire var368;
wire var369;
wire var370;
wire var371;
wire var372;
wire var373;
wire var374;
wire var375;
wire var376;
wire var377;
wire var378;
wire var379;
wire var380;
wire var381;
wire var382;
wire var383;
wire var384;
wire var385;
wire var386;
wire var387;
wire var388;
wire var389;
wire var390;
wire var391;
wire var392;
wire var393;
wire var394;
wire var395;
wire var396;
wire var397;
wire var398;
wire var399;
wire var400;
wire var401;
wire var402;
wire var403;
wire var404;
wire var405;
wire var406;
wire var407;
wire var408;
wire var409;
wire var410;
wire var411;
wire var412;
wire var413;
wire var414;
wire var415;
wire var416;
wire var417;
wire var418;
wire var419;
wire var420;
wire var421;
wire var422;
wire var423;
wire var424;
wire var425;
wire var426;
wire var427;
wire var428;
wire var429;
wire var430;
wire var431;
wire var432;
wire var433;
wire var434;
wire var435;
wire var436;
wire var437;
wire var438;
wire var439;
wire var440;
wire var441;
wire var442;
wire var443;
wire var444;
wire var445;
wire var446;
wire var447;
wire var448;
wire var449;
wire var450;
wire var451;
wire var452;
wire var453;
wire var454;
wire var455;
wire var456;
wire var457;
wire var458;
wire var459;
wire var460;
wire var461;
wire var462;
wire var463;
wire var464;
wire var465;
wire var466;
wire var467;
wire var468;
wire var469;
wire var470;
wire var471;
wire var472;
wire var473;
wire var474;
wire var475;
wire var476;
wire var477;
wire var478;
wire var479;
wire var480;
wire var481;
wire var482;
wire var483;
wire var484;
wire var485;
wire var486;
wire var487;
wire var488;
wire var489;
wire var490;
wire var491;
wire var492;
wire var493;
wire var494;
wire var495;
wire var496;
wire var497;
wire var498;
wire var499;
wire var500;
wire var501;
wire var502;
wire var503;
wire var504;
wire var505;
wire var506;
wire var507;
wire var508;
wire var509;
wire var510;
wire var511;
wire var512;
wire var513;
wire var514;
wire var515;
wire var516;
wire var517;
wire var518;
wire var519;
wire var520;
wire var521;
wire var522;
wire var523;
wire var524;
wire var525;
wire var526;
wire var527;
wire var528;
wire var529;
wire var530;
wire var531;
wire var532;
wire var533;
wire var534;
wire var535;
wire var536;
wire var537;
wire var538;
wire var539;
wire var540;
wire var541;
wire var542;
wire var543;
wire var544;
wire var545;
wire var546;
wire var547;
wire var548;
wire var549;
wire var550;
wire var551;
wire var552;
wire var553;
wire var554;
wire var555;
wire var556;
wire var557;
wire var558;
wire var559;
wire var560;
wire var561;
wire var562;
wire var563;
wire var564;
wire var565;
wire var566;
wire var567;
wire var568;
wire var569;
wire var570;
wire var571;
wire var572;
wire var573;
wire var574;
wire var575;
wire var576;
wire var577;
wire var578;
wire var579;
wire var580;
wire var581;
wire var582;
wire var583;
wire var584;
wire var585;
wire var586;
wire var587;
wire var588;
wire var589;
wire var590;
wire var591;
wire var592;
wire var593;
wire var594;
wire var595;
wire var596;
wire var597;
wire var598;
wire var599;
wire var600;
wire var601;
wire var602;
wire var603;
wire var604;
wire var605;
wire var606;
wire var607;
wire var608;
wire var609;
wire var610;
wire var611;
wire var612;
wire var613;
wire var614;
wire var615;
wire var616;
wire var617;
wire var618;
wire var619;
wire var620;
wire var621;
wire var622;
wire var623;
wire var624;
wire var625;
wire var626;
wire var627;
wire var628;
wire var629;
wire var630;
wire var631;
wire var632;
wire var633;
wire var634;
wire var635;
wire var636;
wire var637;
wire var638;
wire var639;
wire var640;
wire var641;
wire var642;
wire var643;
wire var644;
wire var645;
wire var646;
wire var647;
wire var648;
wire var649;
wire var650;
wire var651;
wire var652;
wire var653;
wire var654;
wire var655;
wire var656;
wire var657;
wire var658;
wire var659;
wire var660;
wire var661;
wire var662;
wire var663;
wire var664;
wire var665;
wire var666;
wire var667;
wire var668;
wire var669;
wire var670;
wire var671;
wire var672;
wire var673;
wire var674;
wire var675;
wire var676;
wire var677;
wire var678;
wire var679;
wire var680;
wire var681;
wire var682;
wire var683;
wire var684;
wire var685;
wire var686;
wire var687;
wire var688;
wire var689;
wire var690;
wire var691;
wire var692;
wire var693;
wire var694;
wire var695;
wire var696;
wire var697;
wire var698;
wire var699;
wire var700;
wire var701;
wire var702;
wire var703;
wire var704;
wire var705;
wire var706;
wire var707;
wire var708;
wire var709;
wire var710;
wire var711;
wire var712;
wire var713;
wire var714;
wire var715;
wire var716;
wire var717;
wire var718;
wire var719;
wire var720;
wire var721;
wire var722;
wire var723;
wire var724;
wire var725;
wire var726;
wire var727;
wire var728;
wire var729;
wire var730;
wire var731;
wire var732;
wire var733;
wire var734;
wire var735;
wire var736;
wire var737;
wire var738;
wire var739;
wire var740;
wire var741;
wire var742;
wire var743;
wire var744;
wire var745;
wire var746;
wire var747;
wire var748;
wire var749;
wire var750;
wire var751;
wire var752;
wire var753;
wire var754;
wire var755;
wire var756;
wire var757;
wire var758;
wire var759;
wire var760;
wire var761;
wire var762;
wire var763;
wire var764;
wire var765;
wire var766;
wire var767;
wire var768;
wire var769;
wire var770;
wire var771;
wire var772;
wire var773;
wire var774;
wire var775;
wire var776;
wire var777;
wire var778;
wire var779;
wire var780;
wire var781;
wire var782;
wire var783;
wire var784;
wire var785;
wire var786;
wire var787;
wire var788;
wire var789;
wire var790;
wire var791;
wire var792;
wire var793;
wire var794;
wire var795;
wire var796;
wire var797;
wire var798;
wire var799;
wire var800;
wire var801;
wire var802;
wire var803;
wire var804;
wire var805;
wire var806;
wire var807;
wire var808;
wire var809;
wire var810;
wire var811;
wire var812;
wire var813;
wire var814;
wire var815;
wire var816;
wire var817;
wire var818;
wire var819;
wire var820;
wire var821;
wire var822;
wire var823;
wire var824;
wire var825;
wire var826;
wire var827;
wire var828;
wire var829;
wire var830;
wire var831;
wire var832;
wire var833;
wire var834;
wire var835;
wire var836;
wire var837;
wire var838;
wire var839;
wire var840;
wire var841;
wire var842;
wire var843;
wire var844;
wire var845;
wire var846;
wire var847;
wire var848;
wire var849;
wire var850;
wire var851;
wire var852;
wire var853;
wire var854;
wire var855;
wire var856;
wire var857;
wire var858;
wire var859;
wire var860;
wire var861;
wire var862;
wire var863;
wire var864;
wire var865;
wire var866;
wire var867;
wire var868;
wire var869;
wire var870;
wire var871;
wire var872;
wire var873;
wire var874;
wire var875;
wire var876;
wire var877;
wire var878;
wire var879;
wire var880;
wire var881;
wire var882;
wire var883;
wire var884;
wire var885;
wire var886;
wire var887;
wire var888;
wire var889;
wire var890;
wire var891;
wire var892;
wire var893;
wire var894;
wire var895;
wire var896;
wire var897;
wire var898;
wire var899;
wire var900;
wire var901;
wire var902;
wire var903;
wire var904;
wire var905;
wire var906;
wire var907;
wire var908;
wire var909;
wire var910;
wire var911;
wire var912;
wire var913;
wire var914;
wire var915;
wire var916;
wire var917;
wire var918;
wire var919;
wire var920;
wire var921;
wire var922;
wire var923;
wire var924;
wire var925;
wire var926;
wire var927;
wire var928;
wire var929;
wire var930;
wire var931;
wire var932;
wire var933;
wire var934;
wire var935;
wire var936;
wire var937;
wire var938;
wire var939;
wire var940;
wire var941;
wire var942;
wire var943;
wire var944;
wire var945;
wire var946;
wire var947;
wire var948;
wire var949;
wire var950;
wire var951;
wire var952;
wire var953;
wire var954;
wire var955;
wire var956;
wire var957;
wire var958;
wire var959;
wire var960;
wire var961;
wire var962;
wire var963;
wire var964;
wire var965;
wire var966;
wire var967;
wire var968;
wire var969;
wire var970;
wire var971;
wire var972;
wire var973;
wire var974;
wire var975;
wire var976;
wire var977;
wire var978;
wire var979;
wire var980;
wire var981;
wire var982;
wire var983;
wire var984;
wire var985;
wire var986;
wire var987;
wire var988;
wire var989;
wire var990;
wire var991;
wire var992;
wire var993;
wire var994;
wire var995;
wire var996;
wire var997;
wire var998;
wire var999;
wire var1000;
wire var1001;
wire var1002;
wire var1003;
wire var1004;
wire var1005;
wire var1006;
wire var1007;
wire var1008;
wire var1009;
wire var1010;
wire var1011;
wire var1012;
wire var1013;
wire var1014;
wire var1015;
wire var1016;
wire var1017;
wire var1018;
wire var1019;
wire var1020;
wire var1021;
wire var1022;
wire var1023;
wire var1024;
wire var1025;
wire var1026;
wire var1027;
wire var1028;
wire var1029;
wire var1030;
wire var1031;
wire var1032;
wire var1033;
wire var1034;
wire var1035;
wire var1036;
wire var1037;
wire var1038;
wire var1039;
wire var1040;
wire var1041;
wire var1042;
wire var1043;
wire var1044;
wire var1045;
wire var1046;
wire var1047;
wire var1048;
wire var1049;
wire var1050;
wire var1051;
wire var1052;
wire var1053;
wire var1054;
wire var1055;
wire var1056;
wire var1057;
wire var1058;
wire var1059;
wire var1060;
wire var1061;
wire var1062;
wire var1063;
wire var1064;
wire var1065;
wire var1066;
wire var1067;
wire var1068;
wire var1069;
wire var1070;
wire var1071;
wire var1072;
wire var1073;
wire var1074;
wire var1075;
wire var1076;
wire var1077;
wire var1078;
wire var1079;
wire var1080;
wire var1081;
wire var1082;
wire var1083;
wire var1084;
wire var1085;
wire var1086;
wire var1087;
wire var1088;
wire var1089;
wire var1090;
wire var1091;
wire var1092;
wire var1093;
wire var1094;
wire var1095;
wire var1096;
wire var1097;
wire var1098;
wire var1099;
wire var1100;
wire var1101;
wire var1102;
wire var1103;
wire var1104;
wire var1105;
wire var1106;
wire var1107;
wire var1108;
wire var1109;
wire var1110;
wire var1111;
wire var1112;
wire var1113;
wire var1114;
wire var1115;
wire var1116;
wire var1117;
wire var1118;
wire var1119;
wire var1120;
wire var1121;
wire var1122;
wire var1123;
wire var1124;
wire var1125;
wire var1126;
wire var1127;
wire var1128;
wire var1129;
wire var1130;
wire var1131;
wire var1132;
wire var1133;
wire var1134;
wire var1135;
wire var1136;
wire var1137;
wire var1138;
wire var1139;
wire var1140;
wire var1141;
wire var1142;
wire var1143;
wire var1144;
wire var1145;
wire var1146;
wire var1147;
wire var1148;
wire var1149;
wire var1150;
wire var1151;
wire var1152;
wire var1153;
wire var1154;
wire var1155;
wire var1156;
wire var1157;
wire var1158;
wire var1159;
wire var1160;
wire var1161;
wire var1162;
wire var1163;
wire var1164;
wire var1165;
wire var1166;
wire var1167;
wire var1168;
wire var1169;
wire var1170;
wire var1171;
wire var1172;
wire var1173;
wire var1174;
wire var1175;
wire var1176;
wire var1177;
wire var1178;
wire var1179;
wire var1180;
wire var1181;
wire var1182;
wire var1183;
wire var1184;
wire var1185;
wire var1186;
wire var1187;
wire var1188;
wire var1189;
wire var1190;
wire var1191;
wire var1192;
wire var1193;
wire var1194;
wire var1195;
wire var1196;
wire var1197;
wire var1198;
wire var1199;
wire var1200;
wire var1201;
wire var1202;
wire var1203;
wire var1204;
wire var1205;
wire var1206;
wire var1207;
wire var1208;
wire var1209;
wire var1210;
wire var1211;
wire var1212;
wire var1213;
wire var1214;
wire var1215;
wire var1216;
wire var1217;
wire var1218;
wire var1219;
wire var1220;
wire var1221;
wire var1222;
wire var1223;
wire var1224;
wire var1225;
wire var1226;
wire var1227;
wire var1228;
wire var1229;
wire var1230;
wire var1231;
wire var1232;
wire var1233;
wire var1234;
wire var1235;
wire var1236;
wire var1237;
wire var1238;
wire var1239;
wire var1240;
wire var1241;
wire var1242;
wire var1243;
wire var1244;
wire var1245;
wire var1246;
wire var1247;
wire var1248;
wire var1249;
wire var1250;
wire var1251;
wire var1252;
wire var1253;
wire var1254;
wire var1255;
wire var1256;
wire var1257;
wire var1258;
wire var1259;
wire var1260;
wire var1261;
wire var1262;
wire var1263;
wire var1264;
wire var1265;
wire var1266;
wire var1267;
wire var1268;
wire var1269;
wire var1270;
wire var1271;
wire var1272;
wire var1273;
wire var1274;
wire var1275;
wire var1276;
wire var1277;
wire var1278;
wire var1279;
wire var1280;
wire var1281;
wire var1282;
wire var1283;
wire var1284;
wire var1285;
wire var1286;
wire var1287;
wire var1288;
wire var1289;
wire var1290;
wire var1291;
wire var1292;
wire var1293;
wire var1294;
wire var1295;
wire var1296;
wire var1297;
wire var1298;
wire var1299;
wire var1300;
wire var1301;
wire var1302;
wire var1303;
wire var1304;
wire var1305;
wire var1306;
wire var1307;
wire var1308;
wire var1309;
wire var1310;
wire var1311;
wire var1312;
wire var1313;
wire var1314;
wire var1315;
wire var1316;
wire var1317;
wire var1318;
wire var1319;
wire var1320;
wire var1321;
wire var1322;
wire var1323;
wire var1324;
wire var1325;
wire var1326;
wire var1327;
wire var1328;
wire var1329;
wire var1330;
wire var1331;
wire var1332;
wire var1333;
wire var1334;
wire var1335;
wire var1336;
wire var1337;
wire var1338;
wire var1339;
wire var1340;
wire var1341;
wire var1342;
wire var1343;
wire var1344;
wire var1345;
wire var1346;
wire var1347;
wire var1348;
wire var1349;
wire var1350;
wire var1351;
wire var1352;
wire var1353;
wire var1354;
wire var1355;
wire var1356;
wire var1357;
wire var1358;
wire var1359;
wire var1360;
wire var1361;
wire var1362;
wire var1363;
wire var1364;
wire var1365;
wire var1366;
wire var1367;
wire var1368;
wire var1369;
wire var1370;
wire var1371;
wire var1372;
wire var1373;
wire var1374;
wire var1375;
wire var1376;
wire var1377;
wire var1378;
wire var1379;
wire var1380;
wire var1381;
wire var1382;
wire var1383;
wire var1384;
wire var1385;
wire var1386;
wire var1387;
wire var1388;
wire var1389;
wire var1390;
wire var1391;
wire var1392;
wire var1393;
wire var1394;
wire var1395;
wire var1396;
wire var1397;
wire var1398;
wire var1399;
wire var1400;
wire var1401;
wire var1402;
wire var1403;
wire var1404;
wire var1405;
wire var1406;
wire var1407;
wire var1408;
wire var1409;
wire var1410;
wire var1411;
wire var1412;
wire var1413;
wire var1414;
wire var1415;
wire var1416;
wire var1417;
wire var1418;
wire var1419;
wire var1420;
wire var1421;
wire var1422;
wire var1423;
wire var1424;
wire var1425;
wire var1426;
wire var1427;
wire var1428;
wire var1429;
wire var1430;
wire var1431;
wire var1432;
wire var1433;
wire var1434;
wire var1435;
wire var1436;
wire var1437;
wire var1438;
wire var1439;
wire var1440;
wire var1441;
wire var1442;
wire var1443;
wire var1444;
wire var1445;
wire var1446;
wire var1447;
wire var1448;
wire var1449;
wire var1450;
wire var1451;
wire var1452;
wire var1453;
wire var1454;
wire var1455;
wire var1456;
wire var1457;
wire var1458;
wire var1459;
wire var1460;
wire var1461;
wire var1462;
wire var1463;
wire var1464;
wire var1465;
wire var1466;
wire var1467;
wire var1468;
wire var1469;
wire var1470;
wire var1471;
wire var1472;
wire var1473;
wire var1474;
wire var1475;
wire var1476;
wire var1477;
wire var1478;
wire var1479;
wire var1480;
wire var1481;
wire var1482;
wire var1483;
wire var1484;
wire var1485;
wire var1486;
wire var1487;
wire var1488;
wire var1489;
wire var1490;
wire var1491;
wire var1492;
wire var1493;
wire var1494;
wire var1495;
wire var1496;
wire var1497;
wire var1498;
wire var1499;
wire var1500;
wire var1501;
wire var1502;
wire var1503;
wire var1504;
wire var1505;
wire var1506;
wire var1507;
wire var1508;
wire var1509;
wire var1510;
wire var1511;
wire var1512;
wire var1513;
wire var1514;
wire var1515;
wire var1516;
wire var1517;
wire var1518;
wire var1519;
wire var1520;
wire var1521;
wire var1522;
wire var1523;
wire var1524;
wire var1525;
wire var1526;
wire var1527;
wire var1528;
wire var1529;
wire var1530;
wire var1531;
wire var1532;
wire var1533;
wire var1534;
wire var1535;
wire var1536;
wire var1537;
wire var1538;
wire var1539;
wire var1540;
wire var1541;
wire var1542;
wire var1543;
wire var1544;
wire var1545;
wire var1546;
wire var1547;
wire var1548;
wire var1549;
wire var1550;
wire var1551;
wire var1552;
wire var1553;
wire var1554;
wire var1555;
wire var1556;
wire var1557;
wire var1558;
wire var1559;
wire var1560;
wire var1561;
wire var1562;
wire var1563;
wire var1564;
wire var1565;
wire var1566;
wire var1567;
wire var1568;
wire var1569;
wire var1570;
wire var1571;
wire var1572;
wire var1573;
wire var1574;
wire var1575;
wire var1576;
wire var1577;
wire var1578;
wire var1579;
wire var1580;
wire var1581;
wire var1582;
wire var1583;
wire var1584;
wire var1585;
wire var1586;
wire var1587;
wire var1588;
wire var1589;
wire var1590;
wire var1591;
wire var1592;
wire var1593;
wire var1594;
wire var1595;
wire var1596;
wire var1597;
wire var1598;
wire var1599;
wire var1600;
wire var1601;
wire var1602;
wire var1603;
wire var1604;
wire var1605;
wire var1606;
wire var1607;
wire var1608;
wire var1609;
wire var1610;
wire var1611;
wire var1612;
wire var1613;
wire var1614;
wire var1615;
wire var1616;
wire var1617;
wire var1618;
wire var1619;
wire var1620;
wire var1621;
wire var1622;
wire var1623;
wire var1624;
wire var1625;
wire var1626;
wire var1627;
wire var1628;
wire var1629;
wire var1630;
wire var1631;
wire var1632;
wire var1633;
wire var1634;
wire var1635;
wire var1636;
wire var1637;
wire var1638;
wire var1639;
wire var1640;
wire var1641;
wire var1642;
wire var1643;
wire var1644;
wire var1645;
wire var1646;
wire var1647;
wire var1648;
wire var1649;
wire var1650;
wire var1651;
wire var1652;
wire var1653;
wire var1654;
wire var1655;
wire var1656;
wire var1657;
wire var1658;
wire var1659;
wire var1660;
wire var1661;
wire var1662;
wire var1663;
wire var1664;
wire var1665;
wire var1666;
wire var1667;
wire var1668;
wire var1669;
wire var1670;
wire var1671;
wire var1672;
wire var1673;
wire var1674;
wire var1675;
wire var1676;
wire var1677;
wire var1678;
wire var1679;
wire var1680;
wire var1681;
wire var1682;
wire var1683;
wire var1684;
wire var1685;
wire var1686;
wire var1687;
wire var1688;
wire var1689;
wire var1690;
wire var1691;
wire var1692;
wire var1693;
wire var1694;
wire var1695;
wire var1696;
wire var1697;
wire var1698;
wire var1699;
wire var1700;
wire var1701;
wire var1702;
wire var1703;
wire var1704;
wire var1705;
wire var1706;
wire var1707;
wire var1708;
wire var1709;
wire var1710;
wire var1711;
wire var1712;
wire var1713;
wire var1714;
wire var1715;
wire var1716;
wire var1717;
wire var1718;
wire var1719;
wire var1720;
wire var1721;
wire var1722;
wire var1723;
wire var1724;
wire var1725;
wire var1726;
wire var1727;
wire var1728;
wire var1729;
wire var1730;
wire var1731;
wire var1732;
wire var1733;
wire var1734;
wire var1735;
wire var1736;
wire var1737;
wire var1738;
wire var1739;
wire var1740;
wire var1741;
wire var1742;
wire var1743;
wire var1744;
wire var1745;
wire var1746;
wire var1747;
wire var1748;
wire var1749;
wire var1750;
wire var1751;
wire var1752;
wire var1753;
wire var1754;
wire var1755;
wire var1756;
wire var1757;
wire var1758;
wire var1759;
wire var1760;
wire var1761;
wire var1762;
wire var1763;
wire var1764;
wire var1765;
wire var1766;
wire var1767;
wire var1768;
wire var1769;
wire var1770;
wire var1771;
wire var1772;
wire var1773;
wire var1774;
wire var1775;
wire var1776;
wire var1777;
wire var1778;
wire var1779;
wire var1780;
wire var1781;
wire var1782;
wire var1783;
wire var1784;
wire var1785;
wire var1786;
wire var1787;
wire var1788;
wire var1789;
wire var1790;
wire var1791;
wire var1792;
wire var1793;
wire var1794;
wire var1795;
wire var1796;
wire var1797;
wire var1798;
wire var1799;
wire var1800;
wire var1801;
wire var1802;
wire var1803;
wire var1804;
wire var1805;
wire var1806;
wire var1807;
wire var1808;
wire var1809;
wire var1810;
wire var1811;
wire var1812;
wire var1813;
wire var1814;
wire var1815;
wire var1816;
wire var1817;
wire var1818;
wire var1819;
wire var1820;
wire var1821;
wire var1822;
wire var1823;
wire var1824;
wire var1825;
wire var1826;
wire var1827;
wire var1828;
wire var1829;
wire var1830;
wire var1831;
wire var1832;
wire var1833;
wire var1834;
wire var1835;
wire var1836;
wire var1837;
wire var1838;
wire var1839;
wire var1840;
wire var1841;
wire var1842;
wire var1843;
wire var1844;
wire var1845;
wire var1846;
wire var1847;
wire var1848;
wire var1849;
wire var1850;
wire var1851;
wire var1852;
wire var1853;
wire var1854;
wire var1855;
wire var1856;
wire var1857;
wire var1858;
wire var1859;
wire var1860;
wire var1861;
wire var1862;
wire var1863;
wire var1864;
wire var1865;
wire var1866;
wire var1867;
wire var1868;
wire var1869;
wire var1870;
wire var1871;
wire var1872;
wire var1873;
wire var1874;
wire var1875;
wire var1876;
wire var1877;
wire var1878;
wire var1879;
wire var1880;
wire var1881;
wire var1882;
wire var1883;
wire var1884;
wire var1885;
wire var1886;
wire var1887;
wire var1888;
wire var1889;
wire var1890;
wire var1891;
wire var1892;
wire var1893;
wire var1894;
wire var1895;
wire var1896;
wire var1897;
wire var1898;
wire var1899;
wire var1900;
wire var1901;
wire var1902;
wire var1903;
wire var1904;
wire var1905;
wire var1906;
wire var1907;
wire var1908;
wire var1909;
wire var1910;
wire var1911;
wire var1912;
wire var1913;
wire var1914;
wire var1915;
wire var1916;
wire var1917;
wire var1918;
wire var1919;
wire var1920;
wire var1921;
wire var1922;
wire var1923;
wire var1924;
wire var1925;
wire var1926;
wire var1927;
wire var1928;
wire var1929;
wire var1930;
wire var1931;
wire var1932;
wire var1933;
wire var1934;
wire var1935;
wire var1936;
wire var1937;
wire var1938;
wire var1939;
wire var1940;
wire var1941;
wire var1942;
wire var1943;
wire var1944;
wire var1945;
wire var1946;
wire var1947;
wire var1948;
wire var1949;
wire var1950;
wire var1951;
wire var1952;
wire var1953;
wire var1954;
wire var1955;
wire var1956;
wire var1957;
wire var1958;
wire var1959;
wire var1960;
wire var1961;
wire var1962;
wire var1963;
wire var1964;
wire var1965;
wire var1966;
wire var1967;
wire var1968;
wire var1969;
wire var1970;
wire var1971;
wire var1972;
wire var1973;
wire var1974;
wire var1975;
wire var1976;
wire var1977;
wire var1978;
wire var1979;
wire var1980;
wire var1981;
wire var1982;
wire var1983;
wire var1984;
wire var1985;
wire var1986;
wire var1987;
wire var1988;
wire var1989;
wire var1990;
wire var1991;
wire var1992;
wire var1993;
wire var1994;
wire var1995;
wire var1996;
wire var1997;
wire var1998;
wire var1999;
wire var2000;
wire var2001;
wire var2002;
wire var2003;
wire var2004;
wire var2005;
wire var2006;
wire var2007;
wire var2008;
wire var2009;
wire var2010;
wire var2011;
wire var2012;
wire var2013;
wire var2014;
wire var2015;
wire var2016;
wire var2017;
wire var2018;
wire var2019;
wire var2020;
wire var2021;
wire var2022;
wire var2023;
wire var2024;
wire var2025;
wire var2026;
wire var2027;
wire var2028;
wire var2029;
wire var2030;
wire var2031;
wire var2032;
wire var2033;
wire var2034;
wire var2035;
wire var2036;
wire var2037;
wire var2038;
wire var2039;
wire var2040;
wire var2041;
wire var2042;
wire var2043;
wire var2044;
wire var2045;
wire var2046;
wire var2047;
wire var2048;
wire var2049;
wire var2050;
wire var2051;
wire var2052;
wire var2053;
wire var2054;
wire var2055;
wire var2056;
wire var2057;
wire var2058;
wire var2059;
wire var2060;
wire var2061;
wire var2062;
wire var2063;
wire var2064;
wire var2065;
wire var2066;
wire var2067;
wire var2068;
wire var2069;
wire var2070;
wire var2071;
wire var2072;
wire var2073;
wire var2074;
wire var2075;
wire var2076;
wire var2077;
wire var2078;
wire var2079;
wire var2080;
wire var2081;
wire var2082;
wire var2083;
wire var2084;
wire var2085;
wire var2086;
wire var2087;
wire var2088;
wire var2089;
wire var2090;
wire var2091;
wire var2092;
wire var2093;
wire var2094;
wire var2095;
wire var2096;
wire var2097;
wire var2098;
wire var2099;
wire var2100;
wire var2101;
wire var2102;
wire var2103;
wire var2104;
wire var2105;
wire var2106;
wire var2107;
wire var2108;
wire var2109;
wire var2110;
wire var2111;
wire var2112;
wire var2113;
wire var2114;
wire var2115;
wire var2116;
wire var2117;
wire var2118;
wire var2119;
wire var2120;
wire var2121;
wire var2122;
wire var2123;
wire var2124;
wire var2125;
wire var2126;
wire var2127;
wire var2128;
wire var2129;
wire var2130;
wire var2131;
wire var2132;
wire var2133;
wire var2134;
wire var2135;
wire var2136;
wire var2137;
wire var2138;
wire var2139;
wire var2140;
wire var2141;
wire var2142;
wire var2143;
wire var2144;
wire var2145;
wire var2146;
wire var2147;
wire var2148;
wire var2149;
wire var2150;
wire var2151;
wire var2152;
wire var2153;
wire var2154;
wire var2155;
wire var2156;
wire var2157;
wire var2158;
wire var2159;
wire var2160;
wire var2161;
wire var2162;
wire var2163;
wire var2164;
wire var2165;
wire var2166;
wire var2167;
wire var2168;
wire var2169;
wire var2170;
wire var2171;
wire var2172;
wire var2173;
wire var2174;
wire var2175;
wire var2176;
wire var2177;
wire var2178;
wire var2179;
wire var2180;
wire var2181;
wire var2182;
wire var2183;
wire var2184;
wire var2185;
wire var2186;
wire var2187;
wire var2188;
wire var2189;
wire var2190;
wire var2191;
wire var2192;
wire var2193;
wire var2194;
wire var2195;
wire var2196;
wire var2197;
wire var2198;
wire var2199;
wire var2200;
wire var2201;
wire var2202;
wire var2203;
wire var2204;
wire var2205;
wire var2206;
wire var2207;
wire var2208;
wire var2209;
wire var2210;
wire var2211;
wire var2212;
wire var2213;
wire var2214;
wire var2215;
wire var2216;
wire var2217;
wire var2218;
wire var2219;
wire var2220;
wire var2221;
wire var2222;
wire var2223;
wire var2224;
wire var2225;
wire var2226;
wire var2227;
wire var2228;
wire var2229;
wire var2230;
wire var2231;
wire var2232;
wire var2233;
wire var2234;
wire var2235;
wire var2236;
wire var2237;
wire var2238;
wire var2239;
wire var2240;
wire var2241;
wire var2242;
wire var2243;
wire var2244;
wire var2245;
wire var2246;
wire var2247;
wire var2248;
wire var2249;
wire var2250;
wire var2251;
wire var2252;
wire var2253;
wire var2254;
wire var2255;
wire var2256;
wire var2257;
wire var2258;
wire var2259;
wire var2260;
wire var2261;
wire var2262;
wire var2263;
wire var2264;
wire var2265;
wire var2266;
wire var2267;
wire var2268;
wire var2269;
wire var2270;
wire var2271;
wire var2272;
wire var2273;
wire var2274;
wire var2275;
wire var2276;
wire var2277;
wire var2278;
wire var2279;
wire var2280;
wire var2281;
wire var2282;
wire var2283;
wire var2284;
wire var2285;
wire var2286;
wire var2287;
wire var2288;
wire var2289;
wire var2290;
wire var2291;
wire var2292;
wire var2293;
wire var2294;
wire var2295;
wire var2296;
wire var2297;
wire var2298;
wire var2299;
wire var2300;
wire var2301;
wire var2302;
wire var2303;
wire var2304;
wire var2305;
wire var2306;
wire var2307;
wire var2308;
wire var2309;
wire var2310;
wire var2311;
wire var2312;
wire var2313;
wire var2314;
wire var2315;
wire var2316;
wire var2317;
wire var2318;
wire var2319;
wire var2320;
wire var2321;
wire var2322;
wire var2323;
wire var2324;
wire var2325;
wire var2326;
wire var2327;
wire var2328;
wire var2329;
wire var2330;
wire var2331;
wire var2332;
wire var2333;
wire var2334;
wire var2335;
wire var2336;
wire var2337;
wire var2338;
wire var2339;
wire var2340;
wire var2341;
wire var2342;
wire var2343;
wire var2344;
wire var2345;
wire var2346;
wire var2347;
wire var2348;
wire var2349;
wire var2350;
wire var2351;
wire var2352;
wire var2353;
wire var2354;
wire var2355;
wire var2356;
wire var2357;
wire var2358;
wire var2359;
wire var2360;
wire var2361;
wire var2362;
wire var2363;
wire var2364;
wire var2365;
wire var2366;
wire var2367;
wire var2368;
wire var2369;
wire var2370;
wire var2371;
wire var2372;
wire var2373;
wire var2374;
wire var2375;
wire var2376;
wire var2377;
wire var2378;
wire var2379;
wire var2380;
wire var2381;
wire var2382;
wire var2383;
wire var2384;
wire var2385;
wire var2386;
wire var2387;
wire var2388;
wire var2389;
wire var2390;
wire var2391;
wire var2392;
wire var2393;
wire var2394;
wire var2395;
wire var2396;
wire var2397;
wire var2398;
wire var2399;
wire var2400;
wire var2401;
wire var2402;
wire var2403;
wire var2404;
wire var2405;
wire var2406;
wire var2407;
wire var2408;
wire var2409;
wire var2410;
wire var2411;
wire var2412;
wire var2413;
wire var2414;
wire var2415;
wire var2416;
wire var2417;
wire var2418;
wire var2419;
wire var2420;
wire var2421;
wire var2422;
wire var2423;
wire var2424;
wire var2425;
wire var2426;
wire var2427;
wire var2428;
wire var2429;
wire var2430;
wire var2431;
wire var2432;
wire var2433;
wire var2434;
wire var2435;
wire var2436;
wire var2437;
wire var2438;
wire var2439;
wire var2440;
wire var2441;
wire var2442;
wire var2443;
wire var2444;
wire var2445;
wire var2446;
wire var2447;
wire var2448;
wire var2449;
wire var2450;
wire var2451;
wire var2452;
wire var2453;
wire var2454;
wire var2455;
wire var2456;
wire var2457;
wire var2458;
wire var2459;
wire var2460;
wire var2461;
wire var2462;
wire var2463;
wire var2464;
wire var2465;
wire var2466;
assign var0 = in255 & in127;
assign var1 = in254 & in126;
assign var2 = in253 & in125;
assign var3 = in252 & in124;
assign var4 = in251 & in123;
assign var5 = in250 & in122;
assign var6 = in249 & in121;
assign var7 = in248 & in120;
assign var8 = in247 & in119;
assign var9 = in246 & in118;
assign var10 = in245 & in117;
assign var11 = in244 & in116;
assign var12 = in243 & in115;
assign var13 = in242 & in114;
assign var14 = in241 & in113;
assign var15 = in240 & in112;
assign var16 = in239 & in111;
assign var17 = in238 & in110;
assign var18 = in237 & in109;
assign var19 = in236 & in108;
assign var20 = in235 & in107;
assign var21 = in234 & in106;
assign var22 = in233 & in105;
assign var23 = in232 & in104;
assign var24 = in231 & in103;
assign var25 = in230 & in102;
assign var26 = in229 & in101;
assign var27 = in228 & in100;
assign var28 = in227 & in99;
assign var29 = in226 & in98;
assign var30 = in225 & in97;
assign var31 = in224 & in96;
assign var32 = in223 & in95;
assign var33 = in222 & in94;
assign var34 = in221 & in93;
assign var35 = in220 & in92;
assign var36 = in219 & in91;
assign var37 = in218 & in90;
assign var38 = in217 & in89;
assign var39 = in216 & in88;
assign var40 = in215 & in87;
assign var41 = in214 & in86;
assign var42 = in213 & in85;
assign var43 = in212 & in84;
assign var44 = in211 & in83;
assign var45 = in210 & in82;
assign var46 = in209 & in81;
assign var47 = in208 & in80;
assign var48 = in207 & in79;
assign var49 = in206 & in78;
assign var50 = in205 & in77;
assign var51 = in204 & in76;
assign var52 = in203 & in75;
assign var53 = in202 & in74;
assign var54 = in201 & in73;
assign var55 = in200 & in72;
assign var56 = in199 & in71;
assign var57 = in198 & in70;
assign var58 = in197 & in69;
assign var59 = in196 & in68;
assign var60 = in195 & in67;
assign var61 = in194 & in66;
assign var62 = in193 & in65;
assign var63 = in192 & in64;
assign var64 = in191 & in63;
assign var65 = in190 & in62;
assign var66 = in189 & in61;
assign var67 = in188 & in60;
assign var68 = in187 & in59;
assign var69 = in186 & in58;
assign var70 = in185 & in57;
assign var71 = in184 & in56;
assign var72 = in183 & in55;
assign var73 = in182 & in54;
assign var74 = in181 & in53;
assign var75 = in180 & in52;
assign var76 = in179 & in51;
assign var77 = in178 & in50;
assign var78 = in177 & in49;
assign var79 = in176 & in48;
assign var80 = in175 & in47;
assign var81 = in174 & in46;
assign var82 = in173 & in45;
assign var83 = in172 & in44;
assign var84 = in171 & in43;
assign var85 = in170 & in42;
assign var86 = in169 & in41;
assign var87 = in168 & in40;
assign var88 = in167 & in39;
assign var89 = in166 & in38;
assign var90 = in165 & in37;
assign var91 = in164 & in36;
assign var92 = in163 & in35;
assign var93 = in162 & in34;
assign var94 = in161 & in33;
assign var95 = in160 & in32;
assign var96 = in159 & in31;
assign var97 = in158 & in30;
assign var98 = in157 & in29;
assign var99 = in156 & in28;
assign var100 = in155 & in27;
assign var101 = in154 & in26;
assign var102 = in153 & in25;
assign var103 = in152 & in24;
assign var104 = in151 & in23;
assign var105 = in150 & in22;
assign var106 = in149 & in21;
assign var107 = in148 & in20;
assign var108 = in147 & in19;
assign var109 = in146 & in18;
assign var110 = in145 & in17;
assign var111 = in144 & in16;
assign var112 = in143 & in15;
assign var113 = in142 & in14;
assign var114 = in141 & in13;
assign var115 = in140 & in12;
assign var116 = in139 & in11;
assign var117 = in138 & in10;
assign var118 = in137 & in9;
assign var119 = in136 & in8;
assign var120 = in135 & in7;
assign var121 = in134 & in6;
assign var122 = in133 & in5;
assign var123 = in132 & in4;
assign var124 = in131 & in3;
assign var125 = in130 & in2;
assign var126 = in129 & in1;
assign var127 = in128 & in0;
assign var128 = in255 ^ in127;
assign var129 = in254 ^ in126;
assign var130 = in253 ^ in125;
assign var131 = in252 ^ in124;
assign var132 = in251 ^ in123;
assign var133 = in250 ^ in122;
assign var134 = in249 ^ in121;
assign var135 = in248 ^ in120;
assign var136 = in247 ^ in119;
assign var137 = in246 ^ in118;
assign var138 = in245 ^ in117;
assign var139 = in244 ^ in116;
assign var140 = in243 ^ in115;
assign var141 = in242 ^ in114;
assign var142 = in241 ^ in113;
assign var143 = in240 ^ in112;
assign var144 = in239 ^ in111;
assign var145 = in238 ^ in110;
assign var146 = in237 ^ in109;
assign var147 = in236 ^ in108;
assign var148 = in235 ^ in107;
assign var149 = in234 ^ in106;
assign var150 = in233 ^ in105;
assign var151 = in232 ^ in104;
assign var152 = in231 ^ in103;
assign var153 = in230 ^ in102;
assign var154 = in229 ^ in101;
assign var155 = in228 ^ in100;
assign var156 = in227 ^ in99;
assign var157 = in226 ^ in98;
assign var158 = in225 ^ in97;
assign var159 = in224 ^ in96;
assign var160 = in223 ^ in95;
assign var161 = in222 ^ in94;
assign var162 = in221 ^ in93;
assign var163 = in220 ^ in92;
assign var164 = in219 ^ in91;
assign var165 = in218 ^ in90;
assign var166 = in217 ^ in89;
assign var167 = in216 ^ in88;
assign var168 = in215 ^ in87;
assign var169 = in214 ^ in86;
assign var170 = in213 ^ in85;
assign var171 = in212 ^ in84;
assign var172 = in211 ^ in83;
assign var173 = in210 ^ in82;
assign var174 = in209 ^ in81;
assign var175 = in208 ^ in80;
assign var176 = in207 ^ in79;
assign var177 = in206 ^ in78;
assign var178 = in205 ^ in77;
assign var179 = in204 ^ in76;
assign var180 = in203 ^ in75;
assign var181 = in202 ^ in74;
assign var182 = in201 ^ in73;
assign var183 = in200 ^ in72;
assign var184 = in199 ^ in71;
assign var185 = in198 ^ in70;
assign var186 = in197 ^ in69;
assign var187 = in196 ^ in68;
assign var188 = in195 ^ in67;
assign var189 = in194 ^ in66;
assign var190 = in193 ^ in65;
assign var191 = in192 ^ in64;
assign var192 = in191 ^ in63;
assign var193 = in190 ^ in62;
assign var194 = in189 ^ in61;
assign var195 = in188 ^ in60;
assign var196 = in187 ^ in59;
assign var197 = in186 ^ in58;
assign var198 = in185 ^ in57;
assign var199 = in184 ^ in56;
assign var200 = in183 ^ in55;
assign var201 = in182 ^ in54;
assign var202 = in181 ^ in53;
assign var203 = in180 ^ in52;
assign var204 = in179 ^ in51;
assign var205 = in178 ^ in50;
assign var206 = in177 ^ in49;
assign var207 = in176 ^ in48;
assign var208 = in175 ^ in47;
assign var209 = in174 ^ in46;
assign var210 = in173 ^ in45;
assign var211 = in172 ^ in44;
assign var212 = in171 ^ in43;
assign var213 = in170 ^ in42;
assign var214 = in169 ^ in41;
assign var215 = in168 ^ in40;
assign var216 = in167 ^ in39;
assign var217 = in166 ^ in38;
assign var218 = in165 ^ in37;
assign var219 = in164 ^ in36;
assign var220 = in163 ^ in35;
assign var221 = in162 ^ in34;
assign var222 = in161 ^ in33;
assign var223 = in160 ^ in32;
assign var224 = in159 ^ in31;
assign var225 = in158 ^ in30;
assign var226 = in157 ^ in29;
assign var227 = in156 ^ in28;
assign var228 = in155 ^ in27;
assign var229 = in154 ^ in26;
assign var230 = in153 ^ in25;
assign var231 = in152 ^ in24;
assign var232 = in151 ^ in23;
assign var233 = in150 ^ in22;
assign var234 = in149 ^ in21;
assign var235 = in148 ^ in20;
assign var236 = in147 ^ in19;
assign var237 = in146 ^ in18;
assign var238 = in145 ^ in17;
assign var239 = in144 ^ in16;
assign var240 = in143 ^ in15;
assign var241 = in142 ^ in14;
assign var242 = in141 ^ in13;
assign var243 = in140 ^ in12;
assign var244 = in139 ^ in11;
assign var245 = in138 ^ in10;
assign var246 = in137 ^ in9;
assign var247 = in136 ^ in8;
assign var248 = in135 ^ in7;
assign var249 = in134 ^ in6;
assign var250 = in133 ^ in5;
assign var251 = in132 ^ in4;
assign var252 = in131 ^ in3;
assign var253 = in130 ^ in2;
assign var254 = in129 ^ in1;
assign var255 = in128 ^ in0;
assign var256 = var255 & var126;
assign var257 = var127 | var256;
assign var258 = var255 & var254;
assign var259 = var254 & var125;
assign var260 = var126 | var259;
assign var261 = var254 & var253;
assign var262 = var253 & var124;
assign var263 = var125 | var262;
assign var264 = var253 & var252;
assign var265 = var252 & var123;
assign var266 = var124 | var265;
assign var267 = var252 & var251;
assign var268 = var251 & var122;
assign var269 = var123 | var268;
assign var270 = var251 & var250;
assign var271 = var250 & var121;
assign var272 = var122 | var271;
assign var273 = var250 & var249;
assign var274 = var249 & var120;
assign var275 = var121 | var274;
assign var276 = var249 & var248;
assign var277 = var248 & var119;
assign var278 = var120 | var277;
assign var279 = var248 & var247;
assign var280 = var247 & var118;
assign var281 = var119 | var280;
assign var282 = var247 & var246;
assign var283 = var246 & var117;
assign var284 = var118 | var283;
assign var285 = var246 & var245;
assign var286 = var245 & var116;
assign var287 = var117 | var286;
assign var288 = var245 & var244;
assign var289 = var244 & var115;
assign var290 = var116 | var289;
assign var291 = var244 & var243;
assign var292 = var243 & var114;
assign var293 = var115 | var292;
assign var294 = var243 & var242;
assign var295 = var242 & var113;
assign var296 = var114 | var295;
assign var297 = var242 & var241;
assign var298 = var241 & var112;
assign var299 = var113 | var298;
assign var300 = var241 & var240;
assign var301 = var240 & var111;
assign var302 = var112 | var301;
assign var303 = var240 & var239;
assign var304 = var239 & var110;
assign var305 = var111 | var304;
assign var306 = var239 & var238;
assign var307 = var238 & var109;
assign var308 = var110 | var307;
assign var309 = var238 & var237;
assign var310 = var237 & var108;
assign var311 = var109 | var310;
assign var312 = var237 & var236;
assign var313 = var236 & var107;
assign var314 = var108 | var313;
assign var315 = var236 & var235;
assign var316 = var235 & var106;
assign var317 = var107 | var316;
assign var318 = var235 & var234;
assign var319 = var234 & var105;
assign var320 = var106 | var319;
assign var321 = var234 & var233;
assign var322 = var233 & var104;
assign var323 = var105 | var322;
assign var324 = var233 & var232;
assign var325 = var232 & var103;
assign var326 = var104 | var325;
assign var327 = var232 & var231;
assign var328 = var231 & var102;
assign var329 = var103 | var328;
assign var330 = var231 & var230;
assign var331 = var230 & var101;
assign var332 = var102 | var331;
assign var333 = var230 & var229;
assign var334 = var229 & var100;
assign var335 = var101 | var334;
assign var336 = var229 & var228;
assign var337 = var228 & var99;
assign var338 = var100 | var337;
assign var339 = var228 & var227;
assign var340 = var227 & var98;
assign var341 = var99 | var340;
assign var342 = var227 & var226;
assign var343 = var226 & var97;
assign var344 = var98 | var343;
assign var345 = var226 & var225;
assign var346 = var225 & var96;
assign var347 = var97 | var346;
assign var348 = var225 & var224;
assign var349 = var224 & var95;
assign var350 = var96 | var349;
assign var351 = var224 & var223;
assign var352 = var223 & var94;
assign var353 = var95 | var352;
assign var354 = var223 & var222;
assign var355 = var222 & var93;
assign var356 = var94 | var355;
assign var357 = var222 & var221;
assign var358 = var221 & var92;
assign var359 = var93 | var358;
assign var360 = var221 & var220;
assign var361 = var220 & var91;
assign var362 = var92 | var361;
assign var363 = var220 & var219;
assign var364 = var219 & var90;
assign var365 = var91 | var364;
assign var366 = var219 & var218;
assign var367 = var218 & var89;
assign var368 = var90 | var367;
assign var369 = var218 & var217;
assign var370 = var217 & var88;
assign var371 = var89 | var370;
assign var372 = var217 & var216;
assign var373 = var216 & var87;
assign var374 = var88 | var373;
assign var375 = var216 & var215;
assign var376 = var215 & var86;
assign var377 = var87 | var376;
assign var378 = var215 & var214;
assign var379 = var214 & var85;
assign var380 = var86 | var379;
assign var381 = var214 & var213;
assign var382 = var213 & var84;
assign var383 = var85 | var382;
assign var384 = var213 & var212;
assign var385 = var212 & var83;
assign var386 = var84 | var385;
assign var387 = var212 & var211;
assign var388 = var211 & var82;
assign var389 = var83 | var388;
assign var390 = var211 & var210;
assign var391 = var210 & var81;
assign var392 = var82 | var391;
assign var393 = var210 & var209;
assign var394 = var209 & var80;
assign var395 = var81 | var394;
assign var396 = var209 & var208;
assign var397 = var208 & var79;
assign var398 = var80 | var397;
assign var399 = var208 & var207;
assign var400 = var207 & var78;
assign var401 = var79 | var400;
assign var402 = var207 & var206;
assign var403 = var206 & var77;
assign var404 = var78 | var403;
assign var405 = var206 & var205;
assign var406 = var205 & var76;
assign var407 = var77 | var406;
assign var408 = var205 & var204;
assign var409 = var204 & var75;
assign var410 = var76 | var409;
assign var411 = var204 & var203;
assign var412 = var203 & var74;
assign var413 = var75 | var412;
assign var414 = var203 & var202;
assign var415 = var202 & var73;
assign var416 = var74 | var415;
assign var417 = var202 & var201;
assign var418 = var201 & var72;
assign var419 = var73 | var418;
assign var420 = var201 & var200;
assign var421 = var200 & var71;
assign var422 = var72 | var421;
assign var423 = var200 & var199;
assign var424 = var199 & var70;
assign var425 = var71 | var424;
assign var426 = var199 & var198;
assign var427 = var198 & var69;
assign var428 = var70 | var427;
assign var429 = var198 & var197;
assign var430 = var197 & var68;
assign var431 = var69 | var430;
assign var432 = var197 & var196;
assign var433 = var196 & var67;
assign var434 = var68 | var433;
assign var435 = var196 & var195;
assign var436 = var195 & var66;
assign var437 = var67 | var436;
assign var438 = var195 & var194;
assign var439 = var194 & var65;
assign var440 = var66 | var439;
assign var441 = var194 & var193;
assign var442 = var193 & var64;
assign var443 = var65 | var442;
assign var444 = var193 & var192;
assign var445 = var192 & var63;
assign var446 = var64 | var445;
assign var447 = var192 & var191;
assign var448 = var191 & var62;
assign var449 = var63 | var448;
assign var450 = var191 & var190;
assign var451 = var190 & var61;
assign var452 = var62 | var451;
assign var453 = var190 & var189;
assign var454 = var189 & var60;
assign var455 = var61 | var454;
assign var456 = var189 & var188;
assign var457 = var188 & var59;
assign var458 = var60 | var457;
assign var459 = var188 & var187;
assign var460 = var187 & var58;
assign var461 = var59 | var460;
assign var462 = var187 & var186;
assign var463 = var186 & var57;
assign var464 = var58 | var463;
assign var465 = var186 & var185;
assign var466 = var185 & var56;
assign var467 = var57 | var466;
assign var468 = var185 & var184;
assign var469 = var184 & var55;
assign var470 = var56 | var469;
assign var471 = var184 & var183;
assign var472 = var183 & var54;
assign var473 = var55 | var472;
assign var474 = var183 & var182;
assign var475 = var182 & var53;
assign var476 = var54 | var475;
assign var477 = var182 & var181;
assign var478 = var181 & var52;
assign var479 = var53 | var478;
assign var480 = var181 & var180;
assign var481 = var180 & var51;
assign var482 = var52 | var481;
assign var483 = var180 & var179;
assign var484 = var179 & var50;
assign var485 = var51 | var484;
assign var486 = var179 & var178;
assign var487 = var178 & var49;
assign var488 = var50 | var487;
assign var489 = var178 & var177;
assign var490 = var177 & var48;
assign var491 = var49 | var490;
assign var492 = var177 & var176;
assign var493 = var176 & var47;
assign var494 = var48 | var493;
assign var495 = var176 & var175;
assign var496 = var175 & var46;
assign var497 = var47 | var496;
assign var498 = var175 & var174;
assign var499 = var174 & var45;
assign var500 = var46 | var499;
assign var501 = var174 & var173;
assign var502 = var173 & var44;
assign var503 = var45 | var502;
assign var504 = var173 & var172;
assign var505 = var172 & var43;
assign var506 = var44 | var505;
assign var507 = var172 & var171;
assign var508 = var171 & var42;
assign var509 = var43 | var508;
assign var510 = var171 & var170;
assign var511 = var170 & var41;
assign var512 = var42 | var511;
assign var513 = var170 & var169;
assign var514 = var169 & var40;
assign var515 = var41 | var514;
assign var516 = var169 & var168;
assign var517 = var168 & var39;
assign var518 = var40 | var517;
assign var519 = var168 & var167;
assign var520 = var167 & var38;
assign var521 = var39 | var520;
assign var522 = var167 & var166;
assign var523 = var166 & var37;
assign var524 = var38 | var523;
assign var525 = var166 & var165;
assign var526 = var165 & var36;
assign var527 = var37 | var526;
assign var528 = var165 & var164;
assign var529 = var164 & var35;
assign var530 = var36 | var529;
assign var531 = var164 & var163;
assign var532 = var163 & var34;
assign var533 = var35 | var532;
assign var534 = var163 & var162;
assign var535 = var162 & var33;
assign var536 = var34 | var535;
assign var537 = var162 & var161;
assign var538 = var161 & var32;
assign var539 = var33 | var538;
assign var540 = var161 & var160;
assign var541 = var160 & var31;
assign var542 = var32 | var541;
assign var543 = var160 & var159;
assign var544 = var159 & var30;
assign var545 = var31 | var544;
assign var546 = var159 & var158;
assign var547 = var158 & var29;
assign var548 = var30 | var547;
assign var549 = var158 & var157;
assign var550 = var157 & var28;
assign var551 = var29 | var550;
assign var552 = var157 & var156;
assign var553 = var156 & var27;
assign var554 = var28 | var553;
assign var555 = var156 & var155;
assign var556 = var155 & var26;
assign var557 = var27 | var556;
assign var558 = var155 & var154;
assign var559 = var154 & var25;
assign var560 = var26 | var559;
assign var561 = var154 & var153;
assign var562 = var153 & var24;
assign var563 = var25 | var562;
assign var564 = var153 & var152;
assign var565 = var152 & var23;
assign var566 = var24 | var565;
assign var567 = var152 & var151;
assign var568 = var151 & var22;
assign var569 = var23 | var568;
assign var570 = var151 & var150;
assign var571 = var150 & var21;
assign var572 = var22 | var571;
assign var573 = var150 & var149;
assign var574 = var149 & var20;
assign var575 = var21 | var574;
assign var576 = var149 & var148;
assign var577 = var148 & var19;
assign var578 = var20 | var577;
assign var579 = var148 & var147;
assign var580 = var147 & var18;
assign var581 = var19 | var580;
assign var582 = var147 & var146;
assign var583 = var146 & var17;
assign var584 = var18 | var583;
assign var585 = var146 & var145;
assign var586 = var145 & var16;
assign var587 = var17 | var586;
assign var588 = var145 & var144;
assign var589 = var144 & var15;
assign var590 = var16 | var589;
assign var591 = var144 & var143;
assign var592 = var143 & var14;
assign var593 = var15 | var592;
assign var594 = var143 & var142;
assign var595 = var142 & var13;
assign var596 = var14 | var595;
assign var597 = var142 & var141;
assign var598 = var141 & var12;
assign var599 = var13 | var598;
assign var600 = var141 & var140;
assign var601 = var140 & var11;
assign var602 = var12 | var601;
assign var603 = var140 & var139;
assign var604 = var139 & var10;
assign var605 = var11 | var604;
assign var606 = var139 & var138;
assign var607 = var138 & var9;
assign var608 = var10 | var607;
assign var609 = var138 & var137;
assign var610 = var137 & var8;
assign var611 = var9 | var610;
assign var612 = var137 & var136;
assign var613 = var136 & var7;
assign var614 = var8 | var613;
assign var615 = var136 & var135;
assign var616 = var135 & var6;
assign var617 = var7 | var616;
assign var618 = var135 & var134;
assign var619 = var134 & var5;
assign var620 = var6 | var619;
assign var621 = var134 & var133;
assign var622 = var133 & var4;
assign var623 = var5 | var622;
assign var624 = var133 & var132;
assign var625 = var132 & var3;
assign var626 = var4 | var625;
assign var627 = var132 & var131;
assign var628 = var131 & var2;
assign var629 = var3 | var628;
assign var630 = var131 & var130;
assign var631 = var130 & var1;
assign var632 = var2 | var631;
assign var633 = var130 & var129;
assign var634 = var129 & var0;
assign var635 = var1 | var634;
assign var636 = var258 & var263;
assign var637 = var257 | var636;
assign var638 = var258 & var264;
assign var639 = var261 & var266;
assign var640 = var260 | var639;
assign var641 = var261 & var267;
assign var642 = var264 & var269;
assign var643 = var263 | var642;
assign var644 = var264 & var270;
assign var645 = var267 & var272;
assign var646 = var266 | var645;
assign var647 = var267 & var273;
assign var648 = var270 & var275;
assign var649 = var269 | var648;
assign var650 = var270 & var276;
assign var651 = var273 & var278;
assign var652 = var272 | var651;
assign var653 = var273 & var279;
assign var654 = var276 & var281;
assign var655 = var275 | var654;
assign var656 = var276 & var282;
assign var657 = var279 & var284;
assign var658 = var278 | var657;
assign var659 = var279 & var285;
assign var660 = var282 & var287;
assign var661 = var281 | var660;
assign var662 = var282 & var288;
assign var663 = var285 & var290;
assign var664 = var284 | var663;
assign var665 = var285 & var291;
assign var666 = var288 & var293;
assign var667 = var287 | var666;
assign var668 = var288 & var294;
assign var669 = var291 & var296;
assign var670 = var290 | var669;
assign var671 = var291 & var297;
assign var672 = var294 & var299;
assign var673 = var293 | var672;
assign var674 = var294 & var300;
assign var675 = var297 & var302;
assign var676 = var296 | var675;
assign var677 = var297 & var303;
assign var678 = var300 & var305;
assign var679 = var299 | var678;
assign var680 = var300 & var306;
assign var681 = var303 & var308;
assign var682 = var302 | var681;
assign var683 = var303 & var309;
assign var684 = var306 & var311;
assign var685 = var305 | var684;
assign var686 = var306 & var312;
assign var687 = var309 & var314;
assign var688 = var308 | var687;
assign var689 = var309 & var315;
assign var690 = var312 & var317;
assign var691 = var311 | var690;
assign var692 = var312 & var318;
assign var693 = var315 & var320;
assign var694 = var314 | var693;
assign var695 = var315 & var321;
assign var696 = var318 & var323;
assign var697 = var317 | var696;
assign var698 = var318 & var324;
assign var699 = var321 & var326;
assign var700 = var320 | var699;
assign var701 = var321 & var327;
assign var702 = var324 & var329;
assign var703 = var323 | var702;
assign var704 = var324 & var330;
assign var705 = var327 & var332;
assign var706 = var326 | var705;
assign var707 = var327 & var333;
assign var708 = var330 & var335;
assign var709 = var329 | var708;
assign var710 = var330 & var336;
assign var711 = var333 & var338;
assign var712 = var332 | var711;
assign var713 = var333 & var339;
assign var714 = var336 & var341;
assign var715 = var335 | var714;
assign var716 = var336 & var342;
assign var717 = var339 & var344;
assign var718 = var338 | var717;
assign var719 = var339 & var345;
assign var720 = var342 & var347;
assign var721 = var341 | var720;
assign var722 = var342 & var348;
assign var723 = var345 & var350;
assign var724 = var344 | var723;
assign var725 = var345 & var351;
assign var726 = var348 & var353;
assign var727 = var347 | var726;
assign var728 = var348 & var354;
assign var729 = var351 & var356;
assign var730 = var350 | var729;
assign var731 = var351 & var357;
assign var732 = var354 & var359;
assign var733 = var353 | var732;
assign var734 = var354 & var360;
assign var735 = var357 & var362;
assign var736 = var356 | var735;
assign var737 = var357 & var363;
assign var738 = var360 & var365;
assign var739 = var359 | var738;
assign var740 = var360 & var366;
assign var741 = var363 & var368;
assign var742 = var362 | var741;
assign var743 = var363 & var369;
assign var744 = var366 & var371;
assign var745 = var365 | var744;
assign var746 = var366 & var372;
assign var747 = var369 & var374;
assign var748 = var368 | var747;
assign var749 = var369 & var375;
assign var750 = var372 & var377;
assign var751 = var371 | var750;
assign var752 = var372 & var378;
assign var753 = var375 & var380;
assign var754 = var374 | var753;
assign var755 = var375 & var381;
assign var756 = var378 & var383;
assign var757 = var377 | var756;
assign var758 = var378 & var384;
assign var759 = var381 & var386;
assign var760 = var380 | var759;
assign var761 = var381 & var387;
assign var762 = var384 & var389;
assign var763 = var383 | var762;
assign var764 = var384 & var390;
assign var765 = var387 & var392;
assign var766 = var386 | var765;
assign var767 = var387 & var393;
assign var768 = var390 & var395;
assign var769 = var389 | var768;
assign var770 = var390 & var396;
assign var771 = var393 & var398;
assign var772 = var392 | var771;
assign var773 = var393 & var399;
assign var774 = var396 & var401;
assign var775 = var395 | var774;
assign var776 = var396 & var402;
assign var777 = var399 & var404;
assign var778 = var398 | var777;
assign var779 = var399 & var405;
assign var780 = var402 & var407;
assign var781 = var401 | var780;
assign var782 = var402 & var408;
assign var783 = var405 & var410;
assign var784 = var404 | var783;
assign var785 = var405 & var411;
assign var786 = var408 & var413;
assign var787 = var407 | var786;
assign var788 = var408 & var414;
assign var789 = var411 & var416;
assign var790 = var410 | var789;
assign var791 = var411 & var417;
assign var792 = var414 & var419;
assign var793 = var413 | var792;
assign var794 = var414 & var420;
assign var795 = var417 & var422;
assign var796 = var416 | var795;
assign var797 = var417 & var423;
assign var798 = var420 & var425;
assign var799 = var419 | var798;
assign var800 = var420 & var426;
assign var801 = var423 & var428;
assign var802 = var422 | var801;
assign var803 = var423 & var429;
assign var804 = var426 & var431;
assign var805 = var425 | var804;
assign var806 = var426 & var432;
assign var807 = var429 & var434;
assign var808 = var428 | var807;
assign var809 = var429 & var435;
assign var810 = var432 & var437;
assign var811 = var431 | var810;
assign var812 = var432 & var438;
assign var813 = var435 & var440;
assign var814 = var434 | var813;
assign var815 = var435 & var441;
assign var816 = var438 & var443;
assign var817 = var437 | var816;
assign var818 = var438 & var444;
assign var819 = var441 & var446;
assign var820 = var440 | var819;
assign var821 = var441 & var447;
assign var822 = var444 & var449;
assign var823 = var443 | var822;
assign var824 = var444 & var450;
assign var825 = var447 & var452;
assign var826 = var446 | var825;
assign var827 = var447 & var453;
assign var828 = var450 & var455;
assign var829 = var449 | var828;
assign var830 = var450 & var456;
assign var831 = var453 & var458;
assign var832 = var452 | var831;
assign var833 = var453 & var459;
assign var834 = var456 & var461;
assign var835 = var455 | var834;
assign var836 = var456 & var462;
assign var837 = var459 & var464;
assign var838 = var458 | var837;
assign var839 = var459 & var465;
assign var840 = var462 & var467;
assign var841 = var461 | var840;
assign var842 = var462 & var468;
assign var843 = var465 & var470;
assign var844 = var464 | var843;
assign var845 = var465 & var471;
assign var846 = var468 & var473;
assign var847 = var467 | var846;
assign var848 = var468 & var474;
assign var849 = var471 & var476;
assign var850 = var470 | var849;
assign var851 = var471 & var477;
assign var852 = var474 & var479;
assign var853 = var473 | var852;
assign var854 = var474 & var480;
assign var855 = var477 & var482;
assign var856 = var476 | var855;
assign var857 = var477 & var483;
assign var858 = var480 & var485;
assign var859 = var479 | var858;
assign var860 = var480 & var486;
assign var861 = var483 & var488;
assign var862 = var482 | var861;
assign var863 = var483 & var489;
assign var864 = var486 & var491;
assign var865 = var485 | var864;
assign var866 = var486 & var492;
assign var867 = var489 & var494;
assign var868 = var488 | var867;
assign var869 = var489 & var495;
assign var870 = var492 & var497;
assign var871 = var491 | var870;
assign var872 = var492 & var498;
assign var873 = var495 & var500;
assign var874 = var494 | var873;
assign var875 = var495 & var501;
assign var876 = var498 & var503;
assign var877 = var497 | var876;
assign var878 = var498 & var504;
assign var879 = var501 & var506;
assign var880 = var500 | var879;
assign var881 = var501 & var507;
assign var882 = var504 & var509;
assign var883 = var503 | var882;
assign var884 = var504 & var510;
assign var885 = var507 & var512;
assign var886 = var506 | var885;
assign var887 = var507 & var513;
assign var888 = var510 & var515;
assign var889 = var509 | var888;
assign var890 = var510 & var516;
assign var891 = var513 & var518;
assign var892 = var512 | var891;
assign var893 = var513 & var519;
assign var894 = var516 & var521;
assign var895 = var515 | var894;
assign var896 = var516 & var522;
assign var897 = var519 & var524;
assign var898 = var518 | var897;
assign var899 = var519 & var525;
assign var900 = var522 & var527;
assign var901 = var521 | var900;
assign var902 = var522 & var528;
assign var903 = var525 & var530;
assign var904 = var524 | var903;
assign var905 = var525 & var531;
assign var906 = var528 & var533;
assign var907 = var527 | var906;
assign var908 = var528 & var534;
assign var909 = var531 & var536;
assign var910 = var530 | var909;
assign var911 = var531 & var537;
assign var912 = var534 & var539;
assign var913 = var533 | var912;
assign var914 = var534 & var540;
assign var915 = var537 & var542;
assign var916 = var536 | var915;
assign var917 = var537 & var543;
assign var918 = var540 & var545;
assign var919 = var539 | var918;
assign var920 = var540 & var546;
assign var921 = var543 & var548;
assign var922 = var542 | var921;
assign var923 = var543 & var549;
assign var924 = var546 & var551;
assign var925 = var545 | var924;
assign var926 = var546 & var552;
assign var927 = var549 & var554;
assign var928 = var548 | var927;
assign var929 = var549 & var555;
assign var930 = var552 & var557;
assign var931 = var551 | var930;
assign var932 = var552 & var558;
assign var933 = var555 & var560;
assign var934 = var554 | var933;
assign var935 = var555 & var561;
assign var936 = var558 & var563;
assign var937 = var557 | var936;
assign var938 = var558 & var564;
assign var939 = var561 & var566;
assign var940 = var560 | var939;
assign var941 = var561 & var567;
assign var942 = var564 & var569;
assign var943 = var563 | var942;
assign var944 = var564 & var570;
assign var945 = var567 & var572;
assign var946 = var566 | var945;
assign var947 = var567 & var573;
assign var948 = var570 & var575;
assign var949 = var569 | var948;
assign var950 = var570 & var576;
assign var951 = var573 & var578;
assign var952 = var572 | var951;
assign var953 = var573 & var579;
assign var954 = var576 & var581;
assign var955 = var575 | var954;
assign var956 = var576 & var582;
assign var957 = var579 & var584;
assign var958 = var578 | var957;
assign var959 = var579 & var585;
assign var960 = var582 & var587;
assign var961 = var581 | var960;
assign var962 = var582 & var588;
assign var963 = var585 & var590;
assign var964 = var584 | var963;
assign var965 = var585 & var591;
assign var966 = var588 & var593;
assign var967 = var587 | var966;
assign var968 = var588 & var594;
assign var969 = var591 & var596;
assign var970 = var590 | var969;
assign var971 = var591 & var597;
assign var972 = var594 & var599;
assign var973 = var593 | var972;
assign var974 = var594 & var600;
assign var975 = var597 & var602;
assign var976 = var596 | var975;
assign var977 = var597 & var603;
assign var978 = var600 & var605;
assign var979 = var599 | var978;
assign var980 = var600 & var606;
assign var981 = var603 & var608;
assign var982 = var602 | var981;
assign var983 = var603 & var609;
assign var984 = var606 & var611;
assign var985 = var605 | var984;
assign var986 = var606 & var612;
assign var987 = var609 & var614;
assign var988 = var608 | var987;
assign var989 = var609 & var615;
assign var990 = var612 & var617;
assign var991 = var611 | var990;
assign var992 = var612 & var618;
assign var993 = var615 & var620;
assign var994 = var614 | var993;
assign var995 = var615 & var621;
assign var996 = var618 & var623;
assign var997 = var617 | var996;
assign var998 = var618 & var624;
assign var999 = var621 & var626;
assign var1000 = var620 | var999;
assign var1001 = var621 & var627;
assign var1002 = var624 & var629;
assign var1003 = var623 | var1002;
assign var1004 = var624 & var630;
assign var1005 = var627 & var632;
assign var1006 = var626 | var1005;
assign var1007 = var627 & var633;
assign var1008 = var630 & var635;
assign var1009 = var629 | var1008;
assign var1010 = var633 & var0;
assign var1011 = var632 | var1010;
assign var1012 = var638 & var649;
assign var1013 = var637 | var1012;
assign var1014 = var638 & var650;
assign var1015 = var641 & var652;
assign var1016 = var640 | var1015;
assign var1017 = var641 & var653;
assign var1018 = var644 & var655;
assign var1019 = var643 | var1018;
assign var1020 = var644 & var656;
assign var1021 = var647 & var658;
assign var1022 = var646 | var1021;
assign var1023 = var647 & var659;
assign var1024 = var650 & var661;
assign var1025 = var649 | var1024;
assign var1026 = var650 & var662;
assign var1027 = var653 & var664;
assign var1028 = var652 | var1027;
assign var1029 = var653 & var665;
assign var1030 = var656 & var667;
assign var1031 = var655 | var1030;
assign var1032 = var656 & var668;
assign var1033 = var659 & var670;
assign var1034 = var658 | var1033;
assign var1035 = var659 & var671;
assign var1036 = var662 & var673;
assign var1037 = var661 | var1036;
assign var1038 = var662 & var674;
assign var1039 = var665 & var676;
assign var1040 = var664 | var1039;
assign var1041 = var665 & var677;
assign var1042 = var668 & var679;
assign var1043 = var667 | var1042;
assign var1044 = var668 & var680;
assign var1045 = var671 & var682;
assign var1046 = var670 | var1045;
assign var1047 = var671 & var683;
assign var1048 = var674 & var685;
assign var1049 = var673 | var1048;
assign var1050 = var674 & var686;
assign var1051 = var677 & var688;
assign var1052 = var676 | var1051;
assign var1053 = var677 & var689;
assign var1054 = var680 & var691;
assign var1055 = var679 | var1054;
assign var1056 = var680 & var692;
assign var1057 = var683 & var694;
assign var1058 = var682 | var1057;
assign var1059 = var683 & var695;
assign var1060 = var686 & var697;
assign var1061 = var685 | var1060;
assign var1062 = var686 & var698;
assign var1063 = var689 & var700;
assign var1064 = var688 | var1063;
assign var1065 = var689 & var701;
assign var1066 = var692 & var703;
assign var1067 = var691 | var1066;
assign var1068 = var692 & var704;
assign var1069 = var695 & var706;
assign var1070 = var694 | var1069;
assign var1071 = var695 & var707;
assign var1072 = var698 & var709;
assign var1073 = var697 | var1072;
assign var1074 = var698 & var710;
assign var1075 = var701 & var712;
assign var1076 = var700 | var1075;
assign var1077 = var701 & var713;
assign var1078 = var704 & var715;
assign var1079 = var703 | var1078;
assign var1080 = var704 & var716;
assign var1081 = var707 & var718;
assign var1082 = var706 | var1081;
assign var1083 = var707 & var719;
assign var1084 = var710 & var721;
assign var1085 = var709 | var1084;
assign var1086 = var710 & var722;
assign var1087 = var713 & var724;
assign var1088 = var712 | var1087;
assign var1089 = var713 & var725;
assign var1090 = var716 & var727;
assign var1091 = var715 | var1090;
assign var1092 = var716 & var728;
assign var1093 = var719 & var730;
assign var1094 = var718 | var1093;
assign var1095 = var719 & var731;
assign var1096 = var722 & var733;
assign var1097 = var721 | var1096;
assign var1098 = var722 & var734;
assign var1099 = var725 & var736;
assign var1100 = var724 | var1099;
assign var1101 = var725 & var737;
assign var1102 = var728 & var739;
assign var1103 = var727 | var1102;
assign var1104 = var728 & var740;
assign var1105 = var731 & var742;
assign var1106 = var730 | var1105;
assign var1107 = var731 & var743;
assign var1108 = var734 & var745;
assign var1109 = var733 | var1108;
assign var1110 = var734 & var746;
assign var1111 = var737 & var748;
assign var1112 = var736 | var1111;
assign var1113 = var737 & var749;
assign var1114 = var740 & var751;
assign var1115 = var739 | var1114;
assign var1116 = var740 & var752;
assign var1117 = var743 & var754;
assign var1118 = var742 | var1117;
assign var1119 = var743 & var755;
assign var1120 = var746 & var757;
assign var1121 = var745 | var1120;
assign var1122 = var746 & var758;
assign var1123 = var749 & var760;
assign var1124 = var748 | var1123;
assign var1125 = var749 & var761;
assign var1126 = var752 & var763;
assign var1127 = var751 | var1126;
assign var1128 = var752 & var764;
assign var1129 = var755 & var766;
assign var1130 = var754 | var1129;
assign var1131 = var755 & var767;
assign var1132 = var758 & var769;
assign var1133 = var757 | var1132;
assign var1134 = var758 & var770;
assign var1135 = var761 & var772;
assign var1136 = var760 | var1135;
assign var1137 = var761 & var773;
assign var1138 = var764 & var775;
assign var1139 = var763 | var1138;
assign var1140 = var764 & var776;
assign var1141 = var767 & var778;
assign var1142 = var766 | var1141;
assign var1143 = var767 & var779;
assign var1144 = var770 & var781;
assign var1145 = var769 | var1144;
assign var1146 = var770 & var782;
assign var1147 = var773 & var784;
assign var1148 = var772 | var1147;
assign var1149 = var773 & var785;
assign var1150 = var776 & var787;
assign var1151 = var775 | var1150;
assign var1152 = var776 & var788;
assign var1153 = var779 & var790;
assign var1154 = var778 | var1153;
assign var1155 = var779 & var791;
assign var1156 = var782 & var793;
assign var1157 = var781 | var1156;
assign var1158 = var782 & var794;
assign var1159 = var785 & var796;
assign var1160 = var784 | var1159;
assign var1161 = var785 & var797;
assign var1162 = var788 & var799;
assign var1163 = var787 | var1162;
assign var1164 = var788 & var800;
assign var1165 = var791 & var802;
assign var1166 = var790 | var1165;
assign var1167 = var791 & var803;
assign var1168 = var794 & var805;
assign var1169 = var793 | var1168;
assign var1170 = var794 & var806;
assign var1171 = var797 & var808;
assign var1172 = var796 | var1171;
assign var1173 = var797 & var809;
assign var1174 = var800 & var811;
assign var1175 = var799 | var1174;
assign var1176 = var800 & var812;
assign var1177 = var803 & var814;
assign var1178 = var802 | var1177;
assign var1179 = var803 & var815;
assign var1180 = var806 & var817;
assign var1181 = var805 | var1180;
assign var1182 = var806 & var818;
assign var1183 = var809 & var820;
assign var1184 = var808 | var1183;
assign var1185 = var809 & var821;
assign var1186 = var812 & var823;
assign var1187 = var811 | var1186;
assign var1188 = var812 & var824;
assign var1189 = var815 & var826;
assign var1190 = var814 | var1189;
assign var1191 = var815 & var827;
assign var1192 = var818 & var829;
assign var1193 = var817 | var1192;
assign var1194 = var818 & var830;
assign var1195 = var821 & var832;
assign var1196 = var820 | var1195;
assign var1197 = var821 & var833;
assign var1198 = var824 & var835;
assign var1199 = var823 | var1198;
assign var1200 = var824 & var836;
assign var1201 = var827 & var838;
assign var1202 = var826 | var1201;
assign var1203 = var827 & var839;
assign var1204 = var830 & var841;
assign var1205 = var829 | var1204;
assign var1206 = var830 & var842;
assign var1207 = var833 & var844;
assign var1208 = var832 | var1207;
assign var1209 = var833 & var845;
assign var1210 = var836 & var847;
assign var1211 = var835 | var1210;
assign var1212 = var836 & var848;
assign var1213 = var839 & var850;
assign var1214 = var838 | var1213;
assign var1215 = var839 & var851;
assign var1216 = var842 & var853;
assign var1217 = var841 | var1216;
assign var1218 = var842 & var854;
assign var1219 = var845 & var856;
assign var1220 = var844 | var1219;
assign var1221 = var845 & var857;
assign var1222 = var848 & var859;
assign var1223 = var847 | var1222;
assign var1224 = var848 & var860;
assign var1225 = var851 & var862;
assign var1226 = var850 | var1225;
assign var1227 = var851 & var863;
assign var1228 = var854 & var865;
assign var1229 = var853 | var1228;
assign var1230 = var854 & var866;
assign var1231 = var857 & var868;
assign var1232 = var856 | var1231;
assign var1233 = var857 & var869;
assign var1234 = var860 & var871;
assign var1235 = var859 | var1234;
assign var1236 = var860 & var872;
assign var1237 = var863 & var874;
assign var1238 = var862 | var1237;
assign var1239 = var863 & var875;
assign var1240 = var866 & var877;
assign var1241 = var865 | var1240;
assign var1242 = var866 & var878;
assign var1243 = var869 & var880;
assign var1244 = var868 | var1243;
assign var1245 = var869 & var881;
assign var1246 = var872 & var883;
assign var1247 = var871 | var1246;
assign var1248 = var872 & var884;
assign var1249 = var875 & var886;
assign var1250 = var874 | var1249;
assign var1251 = var875 & var887;
assign var1252 = var878 & var889;
assign var1253 = var877 | var1252;
assign var1254 = var878 & var890;
assign var1255 = var881 & var892;
assign var1256 = var880 | var1255;
assign var1257 = var881 & var893;
assign var1258 = var884 & var895;
assign var1259 = var883 | var1258;
assign var1260 = var884 & var896;
assign var1261 = var887 & var898;
assign var1262 = var886 | var1261;
assign var1263 = var887 & var899;
assign var1264 = var890 & var901;
assign var1265 = var889 | var1264;
assign var1266 = var890 & var902;
assign var1267 = var893 & var904;
assign var1268 = var892 | var1267;
assign var1269 = var893 & var905;
assign var1270 = var896 & var907;
assign var1271 = var895 | var1270;
assign var1272 = var896 & var908;
assign var1273 = var899 & var910;
assign var1274 = var898 | var1273;
assign var1275 = var899 & var911;
assign var1276 = var902 & var913;
assign var1277 = var901 | var1276;
assign var1278 = var902 & var914;
assign var1279 = var905 & var916;
assign var1280 = var904 | var1279;
assign var1281 = var905 & var917;
assign var1282 = var908 & var919;
assign var1283 = var907 | var1282;
assign var1284 = var908 & var920;
assign var1285 = var911 & var922;
assign var1286 = var910 | var1285;
assign var1287 = var911 & var923;
assign var1288 = var914 & var925;
assign var1289 = var913 | var1288;
assign var1290 = var914 & var926;
assign var1291 = var917 & var928;
assign var1292 = var916 | var1291;
assign var1293 = var917 & var929;
assign var1294 = var920 & var931;
assign var1295 = var919 | var1294;
assign var1296 = var920 & var932;
assign var1297 = var923 & var934;
assign var1298 = var922 | var1297;
assign var1299 = var923 & var935;
assign var1300 = var926 & var937;
assign var1301 = var925 | var1300;
assign var1302 = var926 & var938;
assign var1303 = var929 & var940;
assign var1304 = var928 | var1303;
assign var1305 = var929 & var941;
assign var1306 = var932 & var943;
assign var1307 = var931 | var1306;
assign var1308 = var932 & var944;
assign var1309 = var935 & var946;
assign var1310 = var934 | var1309;
assign var1311 = var935 & var947;
assign var1312 = var938 & var949;
assign var1313 = var937 | var1312;
assign var1314 = var938 & var950;
assign var1315 = var941 & var952;
assign var1316 = var940 | var1315;
assign var1317 = var941 & var953;
assign var1318 = var944 & var955;
assign var1319 = var943 | var1318;
assign var1320 = var944 & var956;
assign var1321 = var947 & var958;
assign var1322 = var946 | var1321;
assign var1323 = var947 & var959;
assign var1324 = var950 & var961;
assign var1325 = var949 | var1324;
assign var1326 = var950 & var962;
assign var1327 = var953 & var964;
assign var1328 = var952 | var1327;
assign var1329 = var953 & var965;
assign var1330 = var956 & var967;
assign var1331 = var955 | var1330;
assign var1332 = var956 & var968;
assign var1333 = var959 & var970;
assign var1334 = var958 | var1333;
assign var1335 = var959 & var971;
assign var1336 = var962 & var973;
assign var1337 = var961 | var1336;
assign var1338 = var962 & var974;
assign var1339 = var965 & var976;
assign var1340 = var964 | var1339;
assign var1341 = var965 & var977;
assign var1342 = var968 & var979;
assign var1343 = var967 | var1342;
assign var1344 = var968 & var980;
assign var1345 = var971 & var982;
assign var1346 = var970 | var1345;
assign var1347 = var971 & var983;
assign var1348 = var974 & var985;
assign var1349 = var973 | var1348;
assign var1350 = var974 & var986;
assign var1351 = var977 & var988;
assign var1352 = var976 | var1351;
assign var1353 = var977 & var989;
assign var1354 = var980 & var991;
assign var1355 = var979 | var1354;
assign var1356 = var980 & var992;
assign var1357 = var983 & var994;
assign var1358 = var982 | var1357;
assign var1359 = var983 & var995;
assign var1360 = var986 & var997;
assign var1361 = var985 | var1360;
assign var1362 = var986 & var998;
assign var1363 = var989 & var1000;
assign var1364 = var988 | var1363;
assign var1365 = var989 & var1001;
assign var1366 = var992 & var1003;
assign var1367 = var991 | var1366;
assign var1368 = var992 & var1004;
assign var1369 = var995 & var1006;
assign var1370 = var994 | var1369;
assign var1371 = var995 & var1007;
assign var1372 = var998 & var1009;
assign var1373 = var997 | var1372;
assign var1374 = var1001 & var1011;
assign var1375 = var1000 | var1374;
assign var1376 = var1004 & var635;
assign var1377 = var1003 | var1376;
assign var1378 = var1007 & var0;
assign var1379 = var1006 | var1378;
assign var1380 = var1014 & var1037;
assign var1381 = var1013 | var1380;
assign var1382 = var1014 & var1038;
assign var1383 = var1017 & var1040;
assign var1384 = var1016 | var1383;
assign var1385 = var1017 & var1041;
assign var1386 = var1020 & var1043;
assign var1387 = var1019 | var1386;
assign var1388 = var1020 & var1044;
assign var1389 = var1023 & var1046;
assign var1390 = var1022 | var1389;
assign var1391 = var1023 & var1047;
assign var1392 = var1026 & var1049;
assign var1393 = var1025 | var1392;
assign var1394 = var1026 & var1050;
assign var1395 = var1029 & var1052;
assign var1396 = var1028 | var1395;
assign var1397 = var1029 & var1053;
assign var1398 = var1032 & var1055;
assign var1399 = var1031 | var1398;
assign var1400 = var1032 & var1056;
assign var1401 = var1035 & var1058;
assign var1402 = var1034 | var1401;
assign var1403 = var1035 & var1059;
assign var1404 = var1038 & var1061;
assign var1405 = var1037 | var1404;
assign var1406 = var1038 & var1062;
assign var1407 = var1041 & var1064;
assign var1408 = var1040 | var1407;
assign var1409 = var1041 & var1065;
assign var1410 = var1044 & var1067;
assign var1411 = var1043 | var1410;
assign var1412 = var1044 & var1068;
assign var1413 = var1047 & var1070;
assign var1414 = var1046 | var1413;
assign var1415 = var1047 & var1071;
assign var1416 = var1050 & var1073;
assign var1417 = var1049 | var1416;
assign var1418 = var1050 & var1074;
assign var1419 = var1053 & var1076;
assign var1420 = var1052 | var1419;
assign var1421 = var1053 & var1077;
assign var1422 = var1056 & var1079;
assign var1423 = var1055 | var1422;
assign var1424 = var1056 & var1080;
assign var1425 = var1059 & var1082;
assign var1426 = var1058 | var1425;
assign var1427 = var1059 & var1083;
assign var1428 = var1062 & var1085;
assign var1429 = var1061 | var1428;
assign var1430 = var1062 & var1086;
assign var1431 = var1065 & var1088;
assign var1432 = var1064 | var1431;
assign var1433 = var1065 & var1089;
assign var1434 = var1068 & var1091;
assign var1435 = var1067 | var1434;
assign var1436 = var1068 & var1092;
assign var1437 = var1071 & var1094;
assign var1438 = var1070 | var1437;
assign var1439 = var1071 & var1095;
assign var1440 = var1074 & var1097;
assign var1441 = var1073 | var1440;
assign var1442 = var1074 & var1098;
assign var1443 = var1077 & var1100;
assign var1444 = var1076 | var1443;
assign var1445 = var1077 & var1101;
assign var1446 = var1080 & var1103;
assign var1447 = var1079 | var1446;
assign var1448 = var1080 & var1104;
assign var1449 = var1083 & var1106;
assign var1450 = var1082 | var1449;
assign var1451 = var1083 & var1107;
assign var1452 = var1086 & var1109;
assign var1453 = var1085 | var1452;
assign var1454 = var1086 & var1110;
assign var1455 = var1089 & var1112;
assign var1456 = var1088 | var1455;
assign var1457 = var1089 & var1113;
assign var1458 = var1092 & var1115;
assign var1459 = var1091 | var1458;
assign var1460 = var1092 & var1116;
assign var1461 = var1095 & var1118;
assign var1462 = var1094 | var1461;
assign var1463 = var1095 & var1119;
assign var1464 = var1098 & var1121;
assign var1465 = var1097 | var1464;
assign var1466 = var1098 & var1122;
assign var1467 = var1101 & var1124;
assign var1468 = var1100 | var1467;
assign var1469 = var1101 & var1125;
assign var1470 = var1104 & var1127;
assign var1471 = var1103 | var1470;
assign var1472 = var1104 & var1128;
assign var1473 = var1107 & var1130;
assign var1474 = var1106 | var1473;
assign var1475 = var1107 & var1131;
assign var1476 = var1110 & var1133;
assign var1477 = var1109 | var1476;
assign var1478 = var1110 & var1134;
assign var1479 = var1113 & var1136;
assign var1480 = var1112 | var1479;
assign var1481 = var1113 & var1137;
assign var1482 = var1116 & var1139;
assign var1483 = var1115 | var1482;
assign var1484 = var1116 & var1140;
assign var1485 = var1119 & var1142;
assign var1486 = var1118 | var1485;
assign var1487 = var1119 & var1143;
assign var1488 = var1122 & var1145;
assign var1489 = var1121 | var1488;
assign var1490 = var1122 & var1146;
assign var1491 = var1125 & var1148;
assign var1492 = var1124 | var1491;
assign var1493 = var1125 & var1149;
assign var1494 = var1128 & var1151;
assign var1495 = var1127 | var1494;
assign var1496 = var1128 & var1152;
assign var1497 = var1131 & var1154;
assign var1498 = var1130 | var1497;
assign var1499 = var1131 & var1155;
assign var1500 = var1134 & var1157;
assign var1501 = var1133 | var1500;
assign var1502 = var1134 & var1158;
assign var1503 = var1137 & var1160;
assign var1504 = var1136 | var1503;
assign var1505 = var1137 & var1161;
assign var1506 = var1140 & var1163;
assign var1507 = var1139 | var1506;
assign var1508 = var1140 & var1164;
assign var1509 = var1143 & var1166;
assign var1510 = var1142 | var1509;
assign var1511 = var1143 & var1167;
assign var1512 = var1146 & var1169;
assign var1513 = var1145 | var1512;
assign var1514 = var1146 & var1170;
assign var1515 = var1149 & var1172;
assign var1516 = var1148 | var1515;
assign var1517 = var1149 & var1173;
assign var1518 = var1152 & var1175;
assign var1519 = var1151 | var1518;
assign var1520 = var1152 & var1176;
assign var1521 = var1155 & var1178;
assign var1522 = var1154 | var1521;
assign var1523 = var1155 & var1179;
assign var1524 = var1158 & var1181;
assign var1525 = var1157 | var1524;
assign var1526 = var1158 & var1182;
assign var1527 = var1161 & var1184;
assign var1528 = var1160 | var1527;
assign var1529 = var1161 & var1185;
assign var1530 = var1164 & var1187;
assign var1531 = var1163 | var1530;
assign var1532 = var1164 & var1188;
assign var1533 = var1167 & var1190;
assign var1534 = var1166 | var1533;
assign var1535 = var1167 & var1191;
assign var1536 = var1170 & var1193;
assign var1537 = var1169 | var1536;
assign var1538 = var1170 & var1194;
assign var1539 = var1173 & var1196;
assign var1540 = var1172 | var1539;
assign var1541 = var1173 & var1197;
assign var1542 = var1176 & var1199;
assign var1543 = var1175 | var1542;
assign var1544 = var1176 & var1200;
assign var1545 = var1179 & var1202;
assign var1546 = var1178 | var1545;
assign var1547 = var1179 & var1203;
assign var1548 = var1182 & var1205;
assign var1549 = var1181 | var1548;
assign var1550 = var1182 & var1206;
assign var1551 = var1185 & var1208;
assign var1552 = var1184 | var1551;
assign var1553 = var1185 & var1209;
assign var1554 = var1188 & var1211;
assign var1555 = var1187 | var1554;
assign var1556 = var1188 & var1212;
assign var1557 = var1191 & var1214;
assign var1558 = var1190 | var1557;
assign var1559 = var1191 & var1215;
assign var1560 = var1194 & var1217;
assign var1561 = var1193 | var1560;
assign var1562 = var1194 & var1218;
assign var1563 = var1197 & var1220;
assign var1564 = var1196 | var1563;
assign var1565 = var1197 & var1221;
assign var1566 = var1200 & var1223;
assign var1567 = var1199 | var1566;
assign var1568 = var1200 & var1224;
assign var1569 = var1203 & var1226;
assign var1570 = var1202 | var1569;
assign var1571 = var1203 & var1227;
assign var1572 = var1206 & var1229;
assign var1573 = var1205 | var1572;
assign var1574 = var1206 & var1230;
assign var1575 = var1209 & var1232;
assign var1576 = var1208 | var1575;
assign var1577 = var1209 & var1233;
assign var1578 = var1212 & var1235;
assign var1579 = var1211 | var1578;
assign var1580 = var1212 & var1236;
assign var1581 = var1215 & var1238;
assign var1582 = var1214 | var1581;
assign var1583 = var1215 & var1239;
assign var1584 = var1218 & var1241;
assign var1585 = var1217 | var1584;
assign var1586 = var1218 & var1242;
assign var1587 = var1221 & var1244;
assign var1588 = var1220 | var1587;
assign var1589 = var1221 & var1245;
assign var1590 = var1224 & var1247;
assign var1591 = var1223 | var1590;
assign var1592 = var1224 & var1248;
assign var1593 = var1227 & var1250;
assign var1594 = var1226 | var1593;
assign var1595 = var1227 & var1251;
assign var1596 = var1230 & var1253;
assign var1597 = var1229 | var1596;
assign var1598 = var1230 & var1254;
assign var1599 = var1233 & var1256;
assign var1600 = var1232 | var1599;
assign var1601 = var1233 & var1257;
assign var1602 = var1236 & var1259;
assign var1603 = var1235 | var1602;
assign var1604 = var1236 & var1260;
assign var1605 = var1239 & var1262;
assign var1606 = var1238 | var1605;
assign var1607 = var1239 & var1263;
assign var1608 = var1242 & var1265;
assign var1609 = var1241 | var1608;
assign var1610 = var1242 & var1266;
assign var1611 = var1245 & var1268;
assign var1612 = var1244 | var1611;
assign var1613 = var1245 & var1269;
assign var1614 = var1248 & var1271;
assign var1615 = var1247 | var1614;
assign var1616 = var1248 & var1272;
assign var1617 = var1251 & var1274;
assign var1618 = var1250 | var1617;
assign var1619 = var1251 & var1275;
assign var1620 = var1254 & var1277;
assign var1621 = var1253 | var1620;
assign var1622 = var1254 & var1278;
assign var1623 = var1257 & var1280;
assign var1624 = var1256 | var1623;
assign var1625 = var1257 & var1281;
assign var1626 = var1260 & var1283;
assign var1627 = var1259 | var1626;
assign var1628 = var1260 & var1284;
assign var1629 = var1263 & var1286;
assign var1630 = var1262 | var1629;
assign var1631 = var1263 & var1287;
assign var1632 = var1266 & var1289;
assign var1633 = var1265 | var1632;
assign var1634 = var1266 & var1290;
assign var1635 = var1269 & var1292;
assign var1636 = var1268 | var1635;
assign var1637 = var1269 & var1293;
assign var1638 = var1272 & var1295;
assign var1639 = var1271 | var1638;
assign var1640 = var1272 & var1296;
assign var1641 = var1275 & var1298;
assign var1642 = var1274 | var1641;
assign var1643 = var1275 & var1299;
assign var1644 = var1278 & var1301;
assign var1645 = var1277 | var1644;
assign var1646 = var1278 & var1302;
assign var1647 = var1281 & var1304;
assign var1648 = var1280 | var1647;
assign var1649 = var1281 & var1305;
assign var1650 = var1284 & var1307;
assign var1651 = var1283 | var1650;
assign var1652 = var1284 & var1308;
assign var1653 = var1287 & var1310;
assign var1654 = var1286 | var1653;
assign var1655 = var1287 & var1311;
assign var1656 = var1290 & var1313;
assign var1657 = var1289 | var1656;
assign var1658 = var1290 & var1314;
assign var1659 = var1293 & var1316;
assign var1660 = var1292 | var1659;
assign var1661 = var1293 & var1317;
assign var1662 = var1296 & var1319;
assign var1663 = var1295 | var1662;
assign var1664 = var1296 & var1320;
assign var1665 = var1299 & var1322;
assign var1666 = var1298 | var1665;
assign var1667 = var1299 & var1323;
assign var1668 = var1302 & var1325;
assign var1669 = var1301 | var1668;
assign var1670 = var1302 & var1326;
assign var1671 = var1305 & var1328;
assign var1672 = var1304 | var1671;
assign var1673 = var1305 & var1329;
assign var1674 = var1308 & var1331;
assign var1675 = var1307 | var1674;
assign var1676 = var1308 & var1332;
assign var1677 = var1311 & var1334;
assign var1678 = var1310 | var1677;
assign var1679 = var1311 & var1335;
assign var1680 = var1314 & var1337;
assign var1681 = var1313 | var1680;
assign var1682 = var1314 & var1338;
assign var1683 = var1317 & var1340;
assign var1684 = var1316 | var1683;
assign var1685 = var1317 & var1341;
assign var1686 = var1320 & var1343;
assign var1687 = var1319 | var1686;
assign var1688 = var1320 & var1344;
assign var1689 = var1323 & var1346;
assign var1690 = var1322 | var1689;
assign var1691 = var1323 & var1347;
assign var1692 = var1326 & var1349;
assign var1693 = var1325 | var1692;
assign var1694 = var1326 & var1350;
assign var1695 = var1329 & var1352;
assign var1696 = var1328 | var1695;
assign var1697 = var1329 & var1353;
assign var1698 = var1332 & var1355;
assign var1699 = var1331 | var1698;
assign var1700 = var1332 & var1356;
assign var1701 = var1335 & var1358;
assign var1702 = var1334 | var1701;
assign var1703 = var1335 & var1359;
assign var1704 = var1338 & var1361;
assign var1705 = var1337 | var1704;
assign var1706 = var1338 & var1362;
assign var1707 = var1341 & var1364;
assign var1708 = var1340 | var1707;
assign var1709 = var1341 & var1365;
assign var1710 = var1344 & var1367;
assign var1711 = var1343 | var1710;
assign var1712 = var1344 & var1368;
assign var1713 = var1347 & var1370;
assign var1714 = var1346 | var1713;
assign var1715 = var1347 & var1371;
assign var1716 = var1350 & var1373;
assign var1717 = var1349 | var1716;
assign var1718 = var1353 & var1375;
assign var1719 = var1352 | var1718;
assign var1720 = var1356 & var1377;
assign var1721 = var1355 | var1720;
assign var1722 = var1359 & var1379;
assign var1723 = var1358 | var1722;
assign var1724 = var1362 & var1009;
assign var1725 = var1361 | var1724;
assign var1726 = var1365 & var1011;
assign var1727 = var1364 | var1726;
assign var1728 = var1368 & var635;
assign var1729 = var1367 | var1728;
assign var1730 = var1371 & var0;
assign var1731 = var1370 | var1730;
assign var1732 = var1382 & var1429;
assign var1733 = var1381 | var1732;
assign var1734 = var1382 & var1430;
assign var1735 = var1385 & var1432;
assign var1736 = var1384 | var1735;
assign var1737 = var1385 & var1433;
assign var1738 = var1388 & var1435;
assign var1739 = var1387 | var1738;
assign var1740 = var1388 & var1436;
assign var1741 = var1391 & var1438;
assign var1742 = var1390 | var1741;
assign var1743 = var1391 & var1439;
assign var1744 = var1394 & var1441;
assign var1745 = var1393 | var1744;
assign var1746 = var1394 & var1442;
assign var1747 = var1397 & var1444;
assign var1748 = var1396 | var1747;
assign var1749 = var1397 & var1445;
assign var1750 = var1400 & var1447;
assign var1751 = var1399 | var1750;
assign var1752 = var1400 & var1448;
assign var1753 = var1403 & var1450;
assign var1754 = var1402 | var1753;
assign var1755 = var1403 & var1451;
assign var1756 = var1406 & var1453;
assign var1757 = var1405 | var1756;
assign var1758 = var1406 & var1454;
assign var1759 = var1409 & var1456;
assign var1760 = var1408 | var1759;
assign var1761 = var1409 & var1457;
assign var1762 = var1412 & var1459;
assign var1763 = var1411 | var1762;
assign var1764 = var1412 & var1460;
assign var1765 = var1415 & var1462;
assign var1766 = var1414 | var1765;
assign var1767 = var1415 & var1463;
assign var1768 = var1418 & var1465;
assign var1769 = var1417 | var1768;
assign var1770 = var1418 & var1466;
assign var1771 = var1421 & var1468;
assign var1772 = var1420 | var1771;
assign var1773 = var1421 & var1469;
assign var1774 = var1424 & var1471;
assign var1775 = var1423 | var1774;
assign var1776 = var1424 & var1472;
assign var1777 = var1427 & var1474;
assign var1778 = var1426 | var1777;
assign var1779 = var1427 & var1475;
assign var1780 = var1430 & var1477;
assign var1781 = var1429 | var1780;
assign var1782 = var1430 & var1478;
assign var1783 = var1433 & var1480;
assign var1784 = var1432 | var1783;
assign var1785 = var1433 & var1481;
assign var1786 = var1436 & var1483;
assign var1787 = var1435 | var1786;
assign var1788 = var1436 & var1484;
assign var1789 = var1439 & var1486;
assign var1790 = var1438 | var1789;
assign var1791 = var1439 & var1487;
assign var1792 = var1442 & var1489;
assign var1793 = var1441 | var1792;
assign var1794 = var1442 & var1490;
assign var1795 = var1445 & var1492;
assign var1796 = var1444 | var1795;
assign var1797 = var1445 & var1493;
assign var1798 = var1448 & var1495;
assign var1799 = var1447 | var1798;
assign var1800 = var1448 & var1496;
assign var1801 = var1451 & var1498;
assign var1802 = var1450 | var1801;
assign var1803 = var1451 & var1499;
assign var1804 = var1454 & var1501;
assign var1805 = var1453 | var1804;
assign var1806 = var1454 & var1502;
assign var1807 = var1457 & var1504;
assign var1808 = var1456 | var1807;
assign var1809 = var1457 & var1505;
assign var1810 = var1460 & var1507;
assign var1811 = var1459 | var1810;
assign var1812 = var1460 & var1508;
assign var1813 = var1463 & var1510;
assign var1814 = var1462 | var1813;
assign var1815 = var1463 & var1511;
assign var1816 = var1466 & var1513;
assign var1817 = var1465 | var1816;
assign var1818 = var1466 & var1514;
assign var1819 = var1469 & var1516;
assign var1820 = var1468 | var1819;
assign var1821 = var1469 & var1517;
assign var1822 = var1472 & var1519;
assign var1823 = var1471 | var1822;
assign var1824 = var1472 & var1520;
assign var1825 = var1475 & var1522;
assign var1826 = var1474 | var1825;
assign var1827 = var1475 & var1523;
assign var1828 = var1478 & var1525;
assign var1829 = var1477 | var1828;
assign var1830 = var1478 & var1526;
assign var1831 = var1481 & var1528;
assign var1832 = var1480 | var1831;
assign var1833 = var1481 & var1529;
assign var1834 = var1484 & var1531;
assign var1835 = var1483 | var1834;
assign var1836 = var1484 & var1532;
assign var1837 = var1487 & var1534;
assign var1838 = var1486 | var1837;
assign var1839 = var1487 & var1535;
assign var1840 = var1490 & var1537;
assign var1841 = var1489 | var1840;
assign var1842 = var1490 & var1538;
assign var1843 = var1493 & var1540;
assign var1844 = var1492 | var1843;
assign var1845 = var1493 & var1541;
assign var1846 = var1496 & var1543;
assign var1847 = var1495 | var1846;
assign var1848 = var1496 & var1544;
assign var1849 = var1499 & var1546;
assign var1850 = var1498 | var1849;
assign var1851 = var1499 & var1547;
assign var1852 = var1502 & var1549;
assign var1853 = var1501 | var1852;
assign var1854 = var1502 & var1550;
assign var1855 = var1505 & var1552;
assign var1856 = var1504 | var1855;
assign var1857 = var1505 & var1553;
assign var1858 = var1508 & var1555;
assign var1859 = var1507 | var1858;
assign var1860 = var1508 & var1556;
assign var1861 = var1511 & var1558;
assign var1862 = var1510 | var1861;
assign var1863 = var1511 & var1559;
assign var1864 = var1514 & var1561;
assign var1865 = var1513 | var1864;
assign var1866 = var1514 & var1562;
assign var1867 = var1517 & var1564;
assign var1868 = var1516 | var1867;
assign var1869 = var1517 & var1565;
assign var1870 = var1520 & var1567;
assign var1871 = var1519 | var1870;
assign var1872 = var1520 & var1568;
assign var1873 = var1523 & var1570;
assign var1874 = var1522 | var1873;
assign var1875 = var1523 & var1571;
assign var1876 = var1526 & var1573;
assign var1877 = var1525 | var1876;
assign var1878 = var1526 & var1574;
assign var1879 = var1529 & var1576;
assign var1880 = var1528 | var1879;
assign var1881 = var1529 & var1577;
assign var1882 = var1532 & var1579;
assign var1883 = var1531 | var1882;
assign var1884 = var1532 & var1580;
assign var1885 = var1535 & var1582;
assign var1886 = var1534 | var1885;
assign var1887 = var1535 & var1583;
assign var1888 = var1538 & var1585;
assign var1889 = var1537 | var1888;
assign var1890 = var1538 & var1586;
assign var1891 = var1541 & var1588;
assign var1892 = var1540 | var1891;
assign var1893 = var1541 & var1589;
assign var1894 = var1544 & var1591;
assign var1895 = var1543 | var1894;
assign var1896 = var1544 & var1592;
assign var1897 = var1547 & var1594;
assign var1898 = var1546 | var1897;
assign var1899 = var1547 & var1595;
assign var1900 = var1550 & var1597;
assign var1901 = var1549 | var1900;
assign var1902 = var1550 & var1598;
assign var1903 = var1553 & var1600;
assign var1904 = var1552 | var1903;
assign var1905 = var1553 & var1601;
assign var1906 = var1556 & var1603;
assign var1907 = var1555 | var1906;
assign var1908 = var1556 & var1604;
assign var1909 = var1559 & var1606;
assign var1910 = var1558 | var1909;
assign var1911 = var1559 & var1607;
assign var1912 = var1562 & var1609;
assign var1913 = var1561 | var1912;
assign var1914 = var1562 & var1610;
assign var1915 = var1565 & var1612;
assign var1916 = var1564 | var1915;
assign var1917 = var1565 & var1613;
assign var1918 = var1568 & var1615;
assign var1919 = var1567 | var1918;
assign var1920 = var1568 & var1616;
assign var1921 = var1571 & var1618;
assign var1922 = var1570 | var1921;
assign var1923 = var1571 & var1619;
assign var1924 = var1574 & var1621;
assign var1925 = var1573 | var1924;
assign var1926 = var1574 & var1622;
assign var1927 = var1577 & var1624;
assign var1928 = var1576 | var1927;
assign var1929 = var1577 & var1625;
assign var1930 = var1580 & var1627;
assign var1931 = var1579 | var1930;
assign var1932 = var1580 & var1628;
assign var1933 = var1583 & var1630;
assign var1934 = var1582 | var1933;
assign var1935 = var1583 & var1631;
assign var1936 = var1586 & var1633;
assign var1937 = var1585 | var1936;
assign var1938 = var1586 & var1634;
assign var1939 = var1589 & var1636;
assign var1940 = var1588 | var1939;
assign var1941 = var1589 & var1637;
assign var1942 = var1592 & var1639;
assign var1943 = var1591 | var1942;
assign var1944 = var1592 & var1640;
assign var1945 = var1595 & var1642;
assign var1946 = var1594 | var1945;
assign var1947 = var1595 & var1643;
assign var1948 = var1598 & var1645;
assign var1949 = var1597 | var1948;
assign var1950 = var1598 & var1646;
assign var1951 = var1601 & var1648;
assign var1952 = var1600 | var1951;
assign var1953 = var1601 & var1649;
assign var1954 = var1604 & var1651;
assign var1955 = var1603 | var1954;
assign var1956 = var1604 & var1652;
assign var1957 = var1607 & var1654;
assign var1958 = var1606 | var1957;
assign var1959 = var1607 & var1655;
assign var1960 = var1610 & var1657;
assign var1961 = var1609 | var1960;
assign var1962 = var1610 & var1658;
assign var1963 = var1613 & var1660;
assign var1964 = var1612 | var1963;
assign var1965 = var1613 & var1661;
assign var1966 = var1616 & var1663;
assign var1967 = var1615 | var1966;
assign var1968 = var1616 & var1664;
assign var1969 = var1619 & var1666;
assign var1970 = var1618 | var1969;
assign var1971 = var1619 & var1667;
assign var1972 = var1622 & var1669;
assign var1973 = var1621 | var1972;
assign var1974 = var1622 & var1670;
assign var1975 = var1625 & var1672;
assign var1976 = var1624 | var1975;
assign var1977 = var1625 & var1673;
assign var1978 = var1628 & var1675;
assign var1979 = var1627 | var1978;
assign var1980 = var1628 & var1676;
assign var1981 = var1631 & var1678;
assign var1982 = var1630 | var1981;
assign var1983 = var1631 & var1679;
assign var1984 = var1634 & var1681;
assign var1985 = var1633 | var1984;
assign var1986 = var1634 & var1682;
assign var1987 = var1637 & var1684;
assign var1988 = var1636 | var1987;
assign var1989 = var1637 & var1685;
assign var1990 = var1640 & var1687;
assign var1991 = var1639 | var1990;
assign var1992 = var1640 & var1688;
assign var1993 = var1643 & var1690;
assign var1994 = var1642 | var1993;
assign var1995 = var1643 & var1691;
assign var1996 = var1646 & var1693;
assign var1997 = var1645 | var1996;
assign var1998 = var1646 & var1694;
assign var1999 = var1649 & var1696;
assign var2000 = var1648 | var1999;
assign var2001 = var1649 & var1697;
assign var2002 = var1652 & var1699;
assign var2003 = var1651 | var2002;
assign var2004 = var1652 & var1700;
assign var2005 = var1655 & var1702;
assign var2006 = var1654 | var2005;
assign var2007 = var1655 & var1703;
assign var2008 = var1658 & var1705;
assign var2009 = var1657 | var2008;
assign var2010 = var1658 & var1706;
assign var2011 = var1661 & var1708;
assign var2012 = var1660 | var2011;
assign var2013 = var1661 & var1709;
assign var2014 = var1664 & var1711;
assign var2015 = var1663 | var2014;
assign var2016 = var1664 & var1712;
assign var2017 = var1667 & var1714;
assign var2018 = var1666 | var2017;
assign var2019 = var1667 & var1715;
assign var2020 = var1670 & var1717;
assign var2021 = var1669 | var2020;
assign var2022 = var1673 & var1719;
assign var2023 = var1672 | var2022;
assign var2024 = var1676 & var1721;
assign var2025 = var1675 | var2024;
assign var2026 = var1679 & var1723;
assign var2027 = var1678 | var2026;
assign var2028 = var1682 & var1725;
assign var2029 = var1681 | var2028;
assign var2030 = var1685 & var1727;
assign var2031 = var1684 | var2030;
assign var2032 = var1688 & var1729;
assign var2033 = var1687 | var2032;
assign var2034 = var1691 & var1731;
assign var2035 = var1690 | var2034;
assign var2036 = var1694 & var1373;
assign var2037 = var1693 | var2036;
assign var2038 = var1697 & var1375;
assign var2039 = var1696 | var2038;
assign var2040 = var1700 & var1377;
assign var2041 = var1699 | var2040;
assign var2042 = var1703 & var1379;
assign var2043 = var1702 | var2042;
assign var2044 = var1706 & var1009;
assign var2045 = var1705 | var2044;
assign var2046 = var1709 & var1011;
assign var2047 = var1708 | var2046;
assign var2048 = var1712 & var635;
assign var2049 = var1711 | var2048;
assign var2050 = var1715 & var0;
assign var2051 = var1714 | var2050;
assign var2052 = var1734 & var1829;
assign var2053 = var1733 | var2052;
assign var2054 = var1734 & var1830;
assign var2055 = var1737 & var1832;
assign var2056 = var1736 | var2055;
assign var2057 = var1737 & var1833;
assign var2058 = var1740 & var1835;
assign var2059 = var1739 | var2058;
assign var2060 = var1740 & var1836;
assign var2061 = var1743 & var1838;
assign var2062 = var1742 | var2061;
assign var2063 = var1743 & var1839;
assign var2064 = var1746 & var1841;
assign var2065 = var1745 | var2064;
assign var2066 = var1746 & var1842;
assign var2067 = var1749 & var1844;
assign var2068 = var1748 | var2067;
assign var2069 = var1749 & var1845;
assign var2070 = var1752 & var1847;
assign var2071 = var1751 | var2070;
assign var2072 = var1752 & var1848;
assign var2073 = var1755 & var1850;
assign var2074 = var1754 | var2073;
assign var2075 = var1755 & var1851;
assign var2076 = var1758 & var1853;
assign var2077 = var1757 | var2076;
assign var2078 = var1758 & var1854;
assign var2079 = var1761 & var1856;
assign var2080 = var1760 | var2079;
assign var2081 = var1761 & var1857;
assign var2082 = var1764 & var1859;
assign var2083 = var1763 | var2082;
assign var2084 = var1764 & var1860;
assign var2085 = var1767 & var1862;
assign var2086 = var1766 | var2085;
assign var2087 = var1767 & var1863;
assign var2088 = var1770 & var1865;
assign var2089 = var1769 | var2088;
assign var2090 = var1770 & var1866;
assign var2091 = var1773 & var1868;
assign var2092 = var1772 | var2091;
assign var2093 = var1773 & var1869;
assign var2094 = var1776 & var1871;
assign var2095 = var1775 | var2094;
assign var2096 = var1776 & var1872;
assign var2097 = var1779 & var1874;
assign var2098 = var1778 | var2097;
assign var2099 = var1779 & var1875;
assign var2100 = var1782 & var1877;
assign var2101 = var1781 | var2100;
assign var2102 = var1782 & var1878;
assign var2103 = var1785 & var1880;
assign var2104 = var1784 | var2103;
assign var2105 = var1785 & var1881;
assign var2106 = var1788 & var1883;
assign var2107 = var1787 | var2106;
assign var2108 = var1788 & var1884;
assign var2109 = var1791 & var1886;
assign var2110 = var1790 | var2109;
assign var2111 = var1791 & var1887;
assign var2112 = var1794 & var1889;
assign var2113 = var1793 | var2112;
assign var2114 = var1794 & var1890;
assign var2115 = var1797 & var1892;
assign var2116 = var1796 | var2115;
assign var2117 = var1797 & var1893;
assign var2118 = var1800 & var1895;
assign var2119 = var1799 | var2118;
assign var2120 = var1800 & var1896;
assign var2121 = var1803 & var1898;
assign var2122 = var1802 | var2121;
assign var2123 = var1803 & var1899;
assign var2124 = var1806 & var1901;
assign var2125 = var1805 | var2124;
assign var2126 = var1806 & var1902;
assign var2127 = var1809 & var1904;
assign var2128 = var1808 | var2127;
assign var2129 = var1809 & var1905;
assign var2130 = var1812 & var1907;
assign var2131 = var1811 | var2130;
assign var2132 = var1812 & var1908;
assign var2133 = var1815 & var1910;
assign var2134 = var1814 | var2133;
assign var2135 = var1815 & var1911;
assign var2136 = var1818 & var1913;
assign var2137 = var1817 | var2136;
assign var2138 = var1818 & var1914;
assign var2139 = var1821 & var1916;
assign var2140 = var1820 | var2139;
assign var2141 = var1821 & var1917;
assign var2142 = var1824 & var1919;
assign var2143 = var1823 | var2142;
assign var2144 = var1824 & var1920;
assign var2145 = var1827 & var1922;
assign var2146 = var1826 | var2145;
assign var2147 = var1827 & var1923;
assign var2148 = var1926 & var2021;
assign var2149 = var1925 | var2148;
assign var2150 = var1929 & var2023;
assign var2151 = var1928 | var2150;
assign var2152 = var1932 & var2025;
assign var2153 = var1931 | var2152;
assign var2154 = var1935 & var2027;
assign var2155 = var1934 | var2154;
assign var2156 = var1938 & var2029;
assign var2157 = var1937 | var2156;
assign var2158 = var1941 & var2031;
assign var2159 = var1940 | var2158;
assign var2160 = var1944 & var2033;
assign var2161 = var1943 | var2160;
assign var2162 = var1947 & var2035;
assign var2163 = var1946 | var2162;
assign var2164 = var1950 & var2037;
assign var2165 = var1949 | var2164;
assign var2166 = var1953 & var2039;
assign var2167 = var1952 | var2166;
assign var2168 = var1956 & var2041;
assign var2169 = var1955 | var2168;
assign var2170 = var1959 & var2043;
assign var2171 = var1958 | var2170;
assign var2172 = var1962 & var2045;
assign var2173 = var1961 | var2172;
assign var2174 = var1965 & var2047;
assign var2175 = var1964 | var2174;
assign var2176 = var1968 & var2049;
assign var2177 = var1967 | var2176;
assign var2178 = var1971 & var2051;
assign var2179 = var1970 | var2178;
assign var2180 = var1974 & var1717;
assign var2181 = var1973 | var2180;
assign var2182 = var1977 & var1719;
assign var2183 = var1976 | var2182;
assign var2184 = var1980 & var1721;
assign var2185 = var1979 | var2184;
assign var2186 = var1983 & var1723;
assign var2187 = var1982 | var2186;
assign var2188 = var1986 & var1725;
assign var2189 = var1985 | var2188;
assign var2190 = var1989 & var1727;
assign var2191 = var1988 | var2190;
assign var2192 = var1992 & var1729;
assign var2193 = var1991 | var2192;
assign var2194 = var1995 & var1731;
assign var2195 = var1994 | var2194;
assign var2196 = var1998 & var1373;
assign var2197 = var1997 | var2196;
assign var2198 = var2001 & var1375;
assign var2199 = var2000 | var2198;
assign var2200 = var2004 & var1377;
assign var2201 = var2003 | var2200;
assign var2202 = var2007 & var1379;
assign var2203 = var2006 | var2202;
assign var2204 = var2010 & var1009;
assign var2205 = var2009 | var2204;
assign var2206 = var2013 & var1011;
assign var2207 = var2012 | var2206;
assign var2208 = var2016 & var635;
assign var2209 = var2015 | var2208;
assign var2210 = var2019 & var0;
assign var2211 = var2018 | var2210;
assign var2212 = var2054 & var2149;
assign var2213 = var2053 | var2212;
assign var2214 = var2057 & var2149;
assign var2215 = var2056 | var2214;
assign var2216 = var2060 & var2149;
assign var2217 = var2059 | var2216;
assign var2218 = var2063 & var2149;
assign var2219 = var2062 | var2218;
assign var2220 = var2066 & var2149;
assign var2221 = var2065 | var2220;
assign var2222 = var2069 & var2149;
assign var2223 = var2068 | var2222;
assign var2224 = var2072 & var2149;
assign var2225 = var2071 | var2224;
assign var2226 = var2075 & var2149;
assign var2227 = var2074 | var2226;
assign var2228 = var2078 & var2149;
assign var2229 = var2077 | var2228;
assign var2230 = var2081 & var2149;
assign var2231 = var2080 | var2230;
assign var2232 = var2084 & var2149;
assign var2233 = var2083 | var2232;
assign var2234 = var2087 & var2149;
assign var2235 = var2086 | var2234;
assign var2236 = var2090 & var2149;
assign var2237 = var2089 | var2236;
assign var2238 = var2093 & var2149;
assign var2239 = var2092 | var2238;
assign var2240 = var2096 & var2149;
assign var2241 = var2095 | var2240;
assign var2242 = var2099 & var2149;
assign var2243 = var2098 | var2242;
assign var2244 = var2102 & var2149;
assign var2245 = var2101 | var2244;
assign var2246 = var2105 & var2149;
assign var2247 = var2104 | var2246;
assign var2248 = var2108 & var2149;
assign var2249 = var2107 | var2248;
assign var2250 = var2111 & var2149;
assign var2251 = var2110 | var2250;
assign var2252 = var2114 & var2149;
assign var2253 = var2113 | var2252;
assign var2254 = var2117 & var2149;
assign var2255 = var2116 | var2254;
assign var2256 = var2120 & var2149;
assign var2257 = var2119 | var2256;
assign var2258 = var2123 & var2149;
assign var2259 = var2122 | var2258;
assign var2260 = var2126 & var2149;
assign var2261 = var2125 | var2260;
assign var2262 = var2129 & var2149;
assign var2263 = var2128 | var2262;
assign var2264 = var2132 & var2149;
assign var2265 = var2131 | var2264;
assign var2266 = var2135 & var2149;
assign var2267 = var2134 | var2266;
assign var2268 = var2138 & var2149;
assign var2269 = var2137 | var2268;
assign var2270 = var2141 & var2149;
assign var2271 = var2140 | var2270;
assign var2272 = var2144 & var2149;
assign var2273 = var2143 | var2272;
assign var2274 = var2147 & var2149;
assign var2275 = var2146 | var2274;
assign var2276 = var1830 & var2149;
assign var2277 = var1829 | var2276;
assign var2278 = var1833 & var2149;
assign var2279 = var1832 | var2278;
assign var2280 = var1836 & var2149;
assign var2281 = var1835 | var2280;
assign var2282 = var1839 & var2149;
assign var2283 = var1838 | var2282;
assign var2284 = var1842 & var2149;
assign var2285 = var1841 | var2284;
assign var2286 = var1845 & var2149;
assign var2287 = var1844 | var2286;
assign var2288 = var1848 & var2149;
assign var2289 = var1847 | var2288;
assign var2290 = var1851 & var2149;
assign var2291 = var1850 | var2290;
assign var2292 = var1854 & var2149;
assign var2293 = var1853 | var2292;
assign var2294 = var1857 & var2149;
assign var2295 = var1856 | var2294;
assign var2296 = var1860 & var2149;
assign var2297 = var1859 | var2296;
assign var2298 = var1863 & var2149;
assign var2299 = var1862 | var2298;
assign var2300 = var1866 & var2149;
assign var2301 = var1865 | var2300;
assign var2302 = var1869 & var2149;
assign var2303 = var1868 | var2302;
assign var2304 = var1872 & var2149;
assign var2305 = var1871 | var2304;
assign var2306 = var1875 & var2149;
assign var2307 = var1874 | var2306;
assign var2308 = var1878 & var2149;
assign var2309 = var1877 | var2308;
assign var2310 = var1881 & var2149;
assign var2311 = var1880 | var2310;
assign var2312 = var1884 & var2149;
assign var2313 = var1883 | var2312;
assign var2314 = var1887 & var2149;
assign var2315 = var1886 | var2314;
assign var2316 = var1890 & var2149;
assign var2317 = var1889 | var2316;
assign var2318 = var1893 & var2149;
assign var2319 = var1892 | var2318;
assign var2320 = var1896 & var2149;
assign var2321 = var1895 | var2320;
assign var2322 = var1899 & var2149;
assign var2323 = var1898 | var2322;
assign var2324 = var1902 & var2149;
assign var2325 = var1901 | var2324;
assign var2326 = var1905 & var2149;
assign var2327 = var1904 | var2326;
assign var2328 = var1908 & var2149;
assign var2329 = var1907 | var2328;
assign var2330 = var1911 & var2149;
assign var2331 = var1910 | var2330;
assign var2332 = var1914 & var2149;
assign var2333 = var1913 | var2332;
assign var2334 = var1917 & var2149;
assign var2335 = var1916 | var2334;
assign var2336 = var1920 & var2149;
assign var2337 = var1919 | var2336;
assign var2338 = var1923 & var2149;
assign var2339 = var1922 | var2338;
assign var2340 = var129 ^ var0;
assign var2341 = var130 ^ var635;
assign var2342 = var131 ^ var1011;
assign var2343 = var132 ^ var1009;
assign var2344 = var133 ^ var1379;
assign var2345 = var134 ^ var1377;
assign var2346 = var135 ^ var1375;
assign var2347 = var136 ^ var1373;
assign var2348 = var137 ^ var1731;
assign var2349 = var138 ^ var1729;
assign var2350 = var139 ^ var1727;
assign var2351 = var140 ^ var1725;
assign var2352 = var141 ^ var1723;
assign var2353 = var142 ^ var1721;
assign var2354 = var143 ^ var1719;
assign var2355 = var144 ^ var1717;
assign var2356 = var145 ^ var2051;
assign var2357 = var146 ^ var2049;
assign var2358 = var147 ^ var2047;
assign var2359 = var148 ^ var2045;
assign var2360 = var149 ^ var2043;
assign var2361 = var150 ^ var2041;
assign var2362 = var151 ^ var2039;
assign var2363 = var152 ^ var2037;
assign var2364 = var153 ^ var2035;
assign var2365 = var154 ^ var2033;
assign var2366 = var155 ^ var2031;
assign var2367 = var156 ^ var2029;
assign var2368 = var157 ^ var2027;
assign var2369 = var158 ^ var2025;
assign var2370 = var159 ^ var2023;
assign var2371 = var160 ^ var2021;
assign var2372 = var161 ^ var2211;
assign var2373 = var162 ^ var2209;
assign var2374 = var163 ^ var2207;
assign var2375 = var164 ^ var2205;
assign var2376 = var165 ^ var2203;
assign var2377 = var166 ^ var2201;
assign var2378 = var167 ^ var2199;
assign var2379 = var168 ^ var2197;
assign var2380 = var169 ^ var2195;
assign var2381 = var170 ^ var2193;
assign var2382 = var171 ^ var2191;
assign var2383 = var172 ^ var2189;
assign var2384 = var173 ^ var2187;
assign var2385 = var174 ^ var2185;
assign var2386 = var175 ^ var2183;
assign var2387 = var176 ^ var2181;
assign var2388 = var177 ^ var2179;
assign var2389 = var178 ^ var2177;
assign var2390 = var179 ^ var2175;
assign var2391 = var180 ^ var2173;
assign var2392 = var181 ^ var2171;
assign var2393 = var182 ^ var2169;
assign var2394 = var183 ^ var2167;
assign var2395 = var184 ^ var2165;
assign var2396 = var185 ^ var2163;
assign var2397 = var186 ^ var2161;
assign var2398 = var187 ^ var2159;
assign var2399 = var188 ^ var2157;
assign var2400 = var189 ^ var2155;
assign var2401 = var190 ^ var2153;
assign var2402 = var191 ^ var2151;
assign var2403 = var192 ^ var2149;
assign var2404 = var193 ^ var2339;
assign var2405 = var194 ^ var2337;
assign var2406 = var195 ^ var2335;
assign var2407 = var196 ^ var2333;
assign var2408 = var197 ^ var2331;
assign var2409 = var198 ^ var2329;
assign var2410 = var199 ^ var2327;
assign var2411 = var200 ^ var2325;
assign var2412 = var201 ^ var2323;
assign var2413 = var202 ^ var2321;
assign var2414 = var203 ^ var2319;
assign var2415 = var204 ^ var2317;
assign var2416 = var205 ^ var2315;
assign var2417 = var206 ^ var2313;
assign var2418 = var207 ^ var2311;
assign var2419 = var208 ^ var2309;
assign var2420 = var209 ^ var2307;
assign var2421 = var210 ^ var2305;
assign var2422 = var211 ^ var2303;
assign var2423 = var212 ^ var2301;
assign var2424 = var213 ^ var2299;
assign var2425 = var214 ^ var2297;
assign var2426 = var215 ^ var2295;
assign var2427 = var216 ^ var2293;
assign var2428 = var217 ^ var2291;
assign var2429 = var218 ^ var2289;
assign var2430 = var219 ^ var2287;
assign var2431 = var220 ^ var2285;
assign var2432 = var221 ^ var2283;
assign var2433 = var222 ^ var2281;
assign var2434 = var223 ^ var2279;
assign var2435 = var224 ^ var2277;
assign var2436 = var225 ^ var2275;
assign var2437 = var226 ^ var2273;
assign var2438 = var227 ^ var2271;
assign var2439 = var228 ^ var2269;
assign var2440 = var229 ^ var2267;
assign var2441 = var230 ^ var2265;
assign var2442 = var231 ^ var2263;
assign var2443 = var232 ^ var2261;
assign var2444 = var233 ^ var2259;
assign var2445 = var234 ^ var2257;
assign var2446 = var235 ^ var2255;
assign var2447 = var236 ^ var2253;
assign var2448 = var237 ^ var2251;
assign var2449 = var238 ^ var2249;
assign var2450 = var239 ^ var2247;
assign var2451 = var240 ^ var2245;
assign var2452 = var241 ^ var2243;
assign var2453 = var242 ^ var2241;
assign var2454 = var243 ^ var2239;
assign var2455 = var244 ^ var2237;
assign var2456 = var245 ^ var2235;
assign var2457 = var246 ^ var2233;
assign var2458 = var247 ^ var2231;
assign var2459 = var248 ^ var2229;
assign var2460 = var249 ^ var2227;
assign var2461 = var250 ^ var2225;
assign var2462 = var251 ^ var2223;
assign var2463 = var252 ^ var2221;
assign var2464 = var253 ^ var2219;
assign var2465 = var254 ^ var2217;
assign var2466 = var255 ^ var2215;
assign out0 = var2213;
assign out1 = var2466;
assign out2 = var2465;
assign out3 = var2464;
assign out4 = var2463;
assign out5 = var2462;
assign out6 = var2461;
assign out7 = var2460;
assign out8 = var2459;
assign out9 = var2458;
assign out10 = var2457;
assign out11 = var2456;
assign out12 = var2455;
assign out13 = var2454;
assign out14 = var2453;
assign out15 = var2452;
assign out16 = var2451;
assign out17 = var2450;
assign out18 = var2449;
assign out19 = var2448;
assign out20 = var2447;
assign out21 = var2446;
assign out22 = var2445;
assign out23 = var2444;
assign out24 = var2443;
assign out25 = var2442;
assign out26 = var2441;
assign out27 = var2440;
assign out28 = var2439;
assign out29 = var2438;
assign out30 = var2437;
assign out31 = var2436;
assign out32 = var2435;
assign out33 = var2434;
assign out34 = var2433;
assign out35 = var2432;
assign out36 = var2431;
assign out37 = var2430;
assign out38 = var2429;
assign out39 = var2428;
assign out40 = var2427;
assign out41 = var2426;
assign out42 = var2425;
assign out43 = var2424;
assign out44 = var2423;
assign out45 = var2422;
assign out46 = var2421;
assign out47 = var2420;
assign out48 = var2419;
assign out49 = var2418;
assign out50 = var2417;
assign out51 = var2416;
assign out52 = var2415;
assign out53 = var2414;
assign out54 = var2413;
assign out55 = var2412;
assign out56 = var2411;
assign out57 = var2410;
assign out58 = var2409;
assign out59 = var2408;
assign out60 = var2407;
assign out61 = var2406;
assign out62 = var2405;
assign out63 = var2404;
assign out64 = var2403;
assign out65 = var2402;
assign out66 = var2401;
assign out67 = var2400;
assign out68 = var2399;
assign out69 = var2398;
assign out70 = var2397;
assign out71 = var2396;
assign out72 = var2395;
assign out73 = var2394;
assign out74 = var2393;
assign out75 = var2392;
assign out76 = var2391;
assign out77 = var2390;
assign out78 = var2389;
assign out79 = var2388;
assign out80 = var2387;
assign out81 = var2386;
assign out82 = var2385;
assign out83 = var2384;
assign out84 = var2383;
assign out85 = var2382;
assign out86 = var2381;
assign out87 = var2380;
assign out88 = var2379;
assign out89 = var2378;
assign out90 = var2377;
assign out91 = var2376;
assign out92 = var2375;
assign out93 = var2374;
assign out94 = var2373;
assign out95 = var2372;
assign out96 = var2371;
assign out97 = var2370;
assign out98 = var2369;
assign out99 = var2368;
assign out100 = var2367;
assign out101 = var2366;
assign out102 = var2365;
assign out103 = var2364;
assign out104 = var2363;
assign out105 = var2362;
assign out106 = var2361;
assign out107 = var2360;
assign out108 = var2359;
assign out109 = var2358;
assign out110 = var2357;
assign out111 = var2356;
assign out112 = var2355;
assign out113 = var2354;
assign out114 = var2353;
assign out115 = var2352;
assign out116 = var2351;
assign out117 = var2350;
assign out118 = var2349;
assign out119 = var2348;
assign out120 = var2347;
assign out121 = var2346;
assign out122 = var2345;
assign out123 = var2344;
assign out124 = var2343;
assign out125 = var2342;
assign out126 = var2341;
assign out127 = var2340;
assign out128 = var128;
endmodule 
