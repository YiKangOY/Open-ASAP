module PartialProd(
  input  [63:0] io_multiplicand,
  input  [63:0] io_multiplier,
  output [63:0] io_outs_0,
  output [63:0] io_outs_1,
  output [63:0] io_outs_2,
  output [63:0] io_outs_3,
  output [63:0] io_outs_4,
  output [63:0] io_outs_5,
  output [63:0] io_outs_6,
  output [63:0] io_outs_7,
  output [63:0] io_outs_8,
  output [63:0] io_outs_9,
  output [63:0] io_outs_10,
  output [63:0] io_outs_11,
  output [63:0] io_outs_12,
  output [63:0] io_outs_13,
  output [63:0] io_outs_14,
  output [63:0] io_outs_15,
  output [63:0] io_outs_16,
  output [63:0] io_outs_17,
  output [63:0] io_outs_18,
  output [63:0] io_outs_19,
  output [63:0] io_outs_20,
  output [63:0] io_outs_21,
  output [63:0] io_outs_22,
  output [63:0] io_outs_23,
  output [63:0] io_outs_24,
  output [63:0] io_outs_25,
  output [63:0] io_outs_26,
  output [63:0] io_outs_27,
  output [63:0] io_outs_28,
  output [63:0] io_outs_29,
  output [63:0] io_outs_30,
  output [63:0] io_outs_31,
  output [63:0] io_outs_32,
  output [63:0] io_outs_33,
  output [63:0] io_outs_34,
  output [63:0] io_outs_35,
  output [63:0] io_outs_36,
  output [63:0] io_outs_37,
  output [63:0] io_outs_38,
  output [63:0] io_outs_39,
  output [63:0] io_outs_40,
  output [63:0] io_outs_41,
  output [63:0] io_outs_42,
  output [63:0] io_outs_43,
  output [63:0] io_outs_44,
  output [63:0] io_outs_45,
  output [63:0] io_outs_46,
  output [63:0] io_outs_47,
  output [63:0] io_outs_48,
  output [63:0] io_outs_49,
  output [63:0] io_outs_50,
  output [63:0] io_outs_51,
  output [63:0] io_outs_52,
  output [63:0] io_outs_53,
  output [63:0] io_outs_54,
  output [63:0] io_outs_55,
  output [63:0] io_outs_56,
  output [63:0] io_outs_57,
  output [63:0] io_outs_58,
  output [63:0] io_outs_59,
  output [63:0] io_outs_60,
  output [63:0] io_outs_61,
  output [63:0] io_outs_62,
  output [63:0] io_outs_63
);
  wire  _T_66 = io_multiplicand[0] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_69 = io_multiplicand[1] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_72 = io_multiplicand[2] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_75 = io_multiplicand[3] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_78 = io_multiplicand[4] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_81 = io_multiplicand[5] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_84 = io_multiplicand[6] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_87 = io_multiplicand[7] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_90 = io_multiplicand[8] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_93 = io_multiplicand[9] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_96 = io_multiplicand[10] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_99 = io_multiplicand[11] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_102 = io_multiplicand[12] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_105 = io_multiplicand[13] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_108 = io_multiplicand[14] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_111 = io_multiplicand[15] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_114 = io_multiplicand[16] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_117 = io_multiplicand[17] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_120 = io_multiplicand[18] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_123 = io_multiplicand[19] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_126 = io_multiplicand[20] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_129 = io_multiplicand[21] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_132 = io_multiplicand[22] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_135 = io_multiplicand[23] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_138 = io_multiplicand[24] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_141 = io_multiplicand[25] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_144 = io_multiplicand[26] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_147 = io_multiplicand[27] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_150 = io_multiplicand[28] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_153 = io_multiplicand[29] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_156 = io_multiplicand[30] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_159 = io_multiplicand[31] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_162 = io_multiplicand[32] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_165 = io_multiplicand[33] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_168 = io_multiplicand[34] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_171 = io_multiplicand[35] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_174 = io_multiplicand[36] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_177 = io_multiplicand[37] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_180 = io_multiplicand[38] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_183 = io_multiplicand[39] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_186 = io_multiplicand[40] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_189 = io_multiplicand[41] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_192 = io_multiplicand[42] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_195 = io_multiplicand[43] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_198 = io_multiplicand[44] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_201 = io_multiplicand[45] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_204 = io_multiplicand[46] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_207 = io_multiplicand[47] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_210 = io_multiplicand[48] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_213 = io_multiplicand[49] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_216 = io_multiplicand[50] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_219 = io_multiplicand[51] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_222 = io_multiplicand[52] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_225 = io_multiplicand[53] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_228 = io_multiplicand[54] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_231 = io_multiplicand[55] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_234 = io_multiplicand[56] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_237 = io_multiplicand[57] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_240 = io_multiplicand[58] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_243 = io_multiplicand[59] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_246 = io_multiplicand[60] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_249 = io_multiplicand[61] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_252 = io_multiplicand[62] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_255 = io_multiplicand[63] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire [9:0] _T_264 = {_T_255,_T_252,_T_249,_T_246,_T_243,_T_240,_T_237,_T_234,_T_231,_T_228}; // @[Cat.scala 29:58]
  wire [18:0] _T_273 = {_T_264,_T_225,_T_222,_T_219,_T_216,_T_213,_T_210,_T_207,_T_204,_T_201}; // @[Cat.scala 29:58]
  wire [27:0] _T_282 = {_T_273,_T_198,_T_195,_T_192,_T_189,_T_186,_T_183,_T_180,_T_177,_T_174}; // @[Cat.scala 29:58]
  wire [36:0] _T_291 = {_T_282,_T_171,_T_168,_T_165,_T_162,_T_159,_T_156,_T_153,_T_150,_T_147}; // @[Cat.scala 29:58]
  wire [45:0] _T_300 = {_T_291,_T_144,_T_141,_T_138,_T_135,_T_132,_T_129,_T_126,_T_123,_T_120}; // @[Cat.scala 29:58]
  wire [54:0] _T_309 = {_T_300,_T_117,_T_114,_T_111,_T_108,_T_105,_T_102,_T_99,_T_96,_T_93}; // @[Cat.scala 29:58]
  wire [62:0] _T_317 = {_T_309,_T_90,_T_87,_T_84,_T_81,_T_78,_T_75,_T_72,_T_69}; // @[Cat.scala 29:58]
  wire  _T_385 = io_multiplicand[0] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_388 = io_multiplicand[1] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_391 = io_multiplicand[2] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_394 = io_multiplicand[3] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_397 = io_multiplicand[4] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_400 = io_multiplicand[5] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_403 = io_multiplicand[6] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_406 = io_multiplicand[7] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_409 = io_multiplicand[8] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_412 = io_multiplicand[9] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_415 = io_multiplicand[10] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_418 = io_multiplicand[11] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_421 = io_multiplicand[12] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_424 = io_multiplicand[13] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_427 = io_multiplicand[14] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_430 = io_multiplicand[15] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_433 = io_multiplicand[16] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_436 = io_multiplicand[17] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_439 = io_multiplicand[18] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_442 = io_multiplicand[19] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_445 = io_multiplicand[20] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_448 = io_multiplicand[21] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_451 = io_multiplicand[22] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_454 = io_multiplicand[23] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_457 = io_multiplicand[24] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_460 = io_multiplicand[25] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_463 = io_multiplicand[26] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_466 = io_multiplicand[27] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_469 = io_multiplicand[28] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_472 = io_multiplicand[29] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_475 = io_multiplicand[30] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_478 = io_multiplicand[31] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_481 = io_multiplicand[32] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_484 = io_multiplicand[33] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_487 = io_multiplicand[34] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_490 = io_multiplicand[35] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_493 = io_multiplicand[36] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_496 = io_multiplicand[37] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_499 = io_multiplicand[38] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_502 = io_multiplicand[39] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_505 = io_multiplicand[40] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_508 = io_multiplicand[41] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_511 = io_multiplicand[42] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_514 = io_multiplicand[43] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_517 = io_multiplicand[44] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_520 = io_multiplicand[45] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_523 = io_multiplicand[46] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_526 = io_multiplicand[47] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_529 = io_multiplicand[48] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_532 = io_multiplicand[49] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_535 = io_multiplicand[50] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_538 = io_multiplicand[51] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_541 = io_multiplicand[52] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_544 = io_multiplicand[53] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_547 = io_multiplicand[54] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_550 = io_multiplicand[55] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_553 = io_multiplicand[56] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_556 = io_multiplicand[57] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_559 = io_multiplicand[58] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_562 = io_multiplicand[59] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_565 = io_multiplicand[60] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_568 = io_multiplicand[61] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_571 = io_multiplicand[62] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_574 = io_multiplicand[63] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire [9:0] _T_583 = {_T_574,_T_571,_T_568,_T_565,_T_562,_T_559,_T_556,_T_553,_T_550,_T_547}; // @[Cat.scala 29:58]
  wire [18:0] _T_592 = {_T_583,_T_544,_T_541,_T_538,_T_535,_T_532,_T_529,_T_526,_T_523,_T_520}; // @[Cat.scala 29:58]
  wire [27:0] _T_601 = {_T_592,_T_517,_T_514,_T_511,_T_508,_T_505,_T_502,_T_499,_T_496,_T_493}; // @[Cat.scala 29:58]
  wire [36:0] _T_610 = {_T_601,_T_490,_T_487,_T_484,_T_481,_T_478,_T_475,_T_472,_T_469,_T_466}; // @[Cat.scala 29:58]
  wire [45:0] _T_619 = {_T_610,_T_463,_T_460,_T_457,_T_454,_T_451,_T_448,_T_445,_T_442,_T_439}; // @[Cat.scala 29:58]
  wire [54:0] _T_628 = {_T_619,_T_436,_T_433,_T_430,_T_427,_T_424,_T_421,_T_418,_T_415,_T_412}; // @[Cat.scala 29:58]
  wire [62:0] _T_636 = {_T_628,_T_409,_T_406,_T_403,_T_400,_T_397,_T_394,_T_391,_T_388}; // @[Cat.scala 29:58]
  wire  _T_704 = io_multiplicand[0] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_707 = io_multiplicand[1] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_710 = io_multiplicand[2] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_713 = io_multiplicand[3] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_716 = io_multiplicand[4] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_719 = io_multiplicand[5] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_722 = io_multiplicand[6] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_725 = io_multiplicand[7] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_728 = io_multiplicand[8] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_731 = io_multiplicand[9] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_734 = io_multiplicand[10] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_737 = io_multiplicand[11] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_740 = io_multiplicand[12] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_743 = io_multiplicand[13] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_746 = io_multiplicand[14] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_749 = io_multiplicand[15] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_752 = io_multiplicand[16] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_755 = io_multiplicand[17] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_758 = io_multiplicand[18] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_761 = io_multiplicand[19] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_764 = io_multiplicand[20] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_767 = io_multiplicand[21] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_770 = io_multiplicand[22] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_773 = io_multiplicand[23] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_776 = io_multiplicand[24] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_779 = io_multiplicand[25] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_782 = io_multiplicand[26] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_785 = io_multiplicand[27] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_788 = io_multiplicand[28] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_791 = io_multiplicand[29] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_794 = io_multiplicand[30] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_797 = io_multiplicand[31] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_800 = io_multiplicand[32] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_803 = io_multiplicand[33] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_806 = io_multiplicand[34] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_809 = io_multiplicand[35] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_812 = io_multiplicand[36] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_815 = io_multiplicand[37] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_818 = io_multiplicand[38] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_821 = io_multiplicand[39] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_824 = io_multiplicand[40] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_827 = io_multiplicand[41] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_830 = io_multiplicand[42] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_833 = io_multiplicand[43] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_836 = io_multiplicand[44] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_839 = io_multiplicand[45] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_842 = io_multiplicand[46] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_845 = io_multiplicand[47] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_848 = io_multiplicand[48] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_851 = io_multiplicand[49] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_854 = io_multiplicand[50] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_857 = io_multiplicand[51] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_860 = io_multiplicand[52] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_863 = io_multiplicand[53] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_866 = io_multiplicand[54] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_869 = io_multiplicand[55] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_872 = io_multiplicand[56] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_875 = io_multiplicand[57] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_878 = io_multiplicand[58] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_881 = io_multiplicand[59] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_884 = io_multiplicand[60] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_887 = io_multiplicand[61] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_890 = io_multiplicand[62] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_893 = io_multiplicand[63] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire [9:0] _T_902 = {_T_893,_T_890,_T_887,_T_884,_T_881,_T_878,_T_875,_T_872,_T_869,_T_866}; // @[Cat.scala 29:58]
  wire [18:0] _T_911 = {_T_902,_T_863,_T_860,_T_857,_T_854,_T_851,_T_848,_T_845,_T_842,_T_839}; // @[Cat.scala 29:58]
  wire [27:0] _T_920 = {_T_911,_T_836,_T_833,_T_830,_T_827,_T_824,_T_821,_T_818,_T_815,_T_812}; // @[Cat.scala 29:58]
  wire [36:0] _T_929 = {_T_920,_T_809,_T_806,_T_803,_T_800,_T_797,_T_794,_T_791,_T_788,_T_785}; // @[Cat.scala 29:58]
  wire [45:0] _T_938 = {_T_929,_T_782,_T_779,_T_776,_T_773,_T_770,_T_767,_T_764,_T_761,_T_758}; // @[Cat.scala 29:58]
  wire [54:0] _T_947 = {_T_938,_T_755,_T_752,_T_749,_T_746,_T_743,_T_740,_T_737,_T_734,_T_731}; // @[Cat.scala 29:58]
  wire [62:0] _T_955 = {_T_947,_T_728,_T_725,_T_722,_T_719,_T_716,_T_713,_T_710,_T_707}; // @[Cat.scala 29:58]
  wire  _T_1023 = io_multiplicand[0] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1026 = io_multiplicand[1] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1029 = io_multiplicand[2] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1032 = io_multiplicand[3] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1035 = io_multiplicand[4] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1038 = io_multiplicand[5] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1041 = io_multiplicand[6] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1044 = io_multiplicand[7] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1047 = io_multiplicand[8] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1050 = io_multiplicand[9] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1053 = io_multiplicand[10] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1056 = io_multiplicand[11] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1059 = io_multiplicand[12] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1062 = io_multiplicand[13] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1065 = io_multiplicand[14] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1068 = io_multiplicand[15] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1071 = io_multiplicand[16] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1074 = io_multiplicand[17] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1077 = io_multiplicand[18] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1080 = io_multiplicand[19] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1083 = io_multiplicand[20] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1086 = io_multiplicand[21] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1089 = io_multiplicand[22] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1092 = io_multiplicand[23] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1095 = io_multiplicand[24] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1098 = io_multiplicand[25] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1101 = io_multiplicand[26] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1104 = io_multiplicand[27] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1107 = io_multiplicand[28] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1110 = io_multiplicand[29] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1113 = io_multiplicand[30] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1116 = io_multiplicand[31] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1119 = io_multiplicand[32] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1122 = io_multiplicand[33] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1125 = io_multiplicand[34] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1128 = io_multiplicand[35] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1131 = io_multiplicand[36] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1134 = io_multiplicand[37] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1137 = io_multiplicand[38] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1140 = io_multiplicand[39] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1143 = io_multiplicand[40] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1146 = io_multiplicand[41] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1149 = io_multiplicand[42] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1152 = io_multiplicand[43] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1155 = io_multiplicand[44] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1158 = io_multiplicand[45] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1161 = io_multiplicand[46] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1164 = io_multiplicand[47] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1167 = io_multiplicand[48] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1170 = io_multiplicand[49] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1173 = io_multiplicand[50] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1176 = io_multiplicand[51] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1179 = io_multiplicand[52] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1182 = io_multiplicand[53] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1185 = io_multiplicand[54] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1188 = io_multiplicand[55] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1191 = io_multiplicand[56] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1194 = io_multiplicand[57] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1197 = io_multiplicand[58] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1200 = io_multiplicand[59] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1203 = io_multiplicand[60] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1206 = io_multiplicand[61] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1209 = io_multiplicand[62] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_1212 = io_multiplicand[63] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1221 = {_T_1212,_T_1209,_T_1206,_T_1203,_T_1200,_T_1197,_T_1194,_T_1191,_T_1188,_T_1185}; // @[Cat.scala 29:58]
  wire [18:0] _T_1230 = {_T_1221,_T_1182,_T_1179,_T_1176,_T_1173,_T_1170,_T_1167,_T_1164,_T_1161,_T_1158}; // @[Cat.scala 29:58]
  wire [27:0] _T_1239 = {_T_1230,_T_1155,_T_1152,_T_1149,_T_1146,_T_1143,_T_1140,_T_1137,_T_1134,_T_1131}; // @[Cat.scala 29:58]
  wire [36:0] _T_1248 = {_T_1239,_T_1128,_T_1125,_T_1122,_T_1119,_T_1116,_T_1113,_T_1110,_T_1107,_T_1104}; // @[Cat.scala 29:58]
  wire [45:0] _T_1257 = {_T_1248,_T_1101,_T_1098,_T_1095,_T_1092,_T_1089,_T_1086,_T_1083,_T_1080,_T_1077}; // @[Cat.scala 29:58]
  wire [54:0] _T_1266 = {_T_1257,_T_1074,_T_1071,_T_1068,_T_1065,_T_1062,_T_1059,_T_1056,_T_1053,_T_1050}; // @[Cat.scala 29:58]
  wire [62:0] _T_1274 = {_T_1266,_T_1047,_T_1044,_T_1041,_T_1038,_T_1035,_T_1032,_T_1029,_T_1026}; // @[Cat.scala 29:58]
  wire  _T_1342 = io_multiplicand[0] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1345 = io_multiplicand[1] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1348 = io_multiplicand[2] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1351 = io_multiplicand[3] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1354 = io_multiplicand[4] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1357 = io_multiplicand[5] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1360 = io_multiplicand[6] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1363 = io_multiplicand[7] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1366 = io_multiplicand[8] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1369 = io_multiplicand[9] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1372 = io_multiplicand[10] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1375 = io_multiplicand[11] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1378 = io_multiplicand[12] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1381 = io_multiplicand[13] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1384 = io_multiplicand[14] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1387 = io_multiplicand[15] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1390 = io_multiplicand[16] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1393 = io_multiplicand[17] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1396 = io_multiplicand[18] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1399 = io_multiplicand[19] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1402 = io_multiplicand[20] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1405 = io_multiplicand[21] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1408 = io_multiplicand[22] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1411 = io_multiplicand[23] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1414 = io_multiplicand[24] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1417 = io_multiplicand[25] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1420 = io_multiplicand[26] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1423 = io_multiplicand[27] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1426 = io_multiplicand[28] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1429 = io_multiplicand[29] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1432 = io_multiplicand[30] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1435 = io_multiplicand[31] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1438 = io_multiplicand[32] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1441 = io_multiplicand[33] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1444 = io_multiplicand[34] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1447 = io_multiplicand[35] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1450 = io_multiplicand[36] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1453 = io_multiplicand[37] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1456 = io_multiplicand[38] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1459 = io_multiplicand[39] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1462 = io_multiplicand[40] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1465 = io_multiplicand[41] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1468 = io_multiplicand[42] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1471 = io_multiplicand[43] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1474 = io_multiplicand[44] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1477 = io_multiplicand[45] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1480 = io_multiplicand[46] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1483 = io_multiplicand[47] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1486 = io_multiplicand[48] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1489 = io_multiplicand[49] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1492 = io_multiplicand[50] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1495 = io_multiplicand[51] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1498 = io_multiplicand[52] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1501 = io_multiplicand[53] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1504 = io_multiplicand[54] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1507 = io_multiplicand[55] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1510 = io_multiplicand[56] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1513 = io_multiplicand[57] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1516 = io_multiplicand[58] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1519 = io_multiplicand[59] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1522 = io_multiplicand[60] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1525 = io_multiplicand[61] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1528 = io_multiplicand[62] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_1531 = io_multiplicand[63] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1540 = {_T_1531,_T_1528,_T_1525,_T_1522,_T_1519,_T_1516,_T_1513,_T_1510,_T_1507,_T_1504}; // @[Cat.scala 29:58]
  wire [18:0] _T_1549 = {_T_1540,_T_1501,_T_1498,_T_1495,_T_1492,_T_1489,_T_1486,_T_1483,_T_1480,_T_1477}; // @[Cat.scala 29:58]
  wire [27:0] _T_1558 = {_T_1549,_T_1474,_T_1471,_T_1468,_T_1465,_T_1462,_T_1459,_T_1456,_T_1453,_T_1450}; // @[Cat.scala 29:58]
  wire [36:0] _T_1567 = {_T_1558,_T_1447,_T_1444,_T_1441,_T_1438,_T_1435,_T_1432,_T_1429,_T_1426,_T_1423}; // @[Cat.scala 29:58]
  wire [45:0] _T_1576 = {_T_1567,_T_1420,_T_1417,_T_1414,_T_1411,_T_1408,_T_1405,_T_1402,_T_1399,_T_1396}; // @[Cat.scala 29:58]
  wire [54:0] _T_1585 = {_T_1576,_T_1393,_T_1390,_T_1387,_T_1384,_T_1381,_T_1378,_T_1375,_T_1372,_T_1369}; // @[Cat.scala 29:58]
  wire [62:0] _T_1593 = {_T_1585,_T_1366,_T_1363,_T_1360,_T_1357,_T_1354,_T_1351,_T_1348,_T_1345}; // @[Cat.scala 29:58]
  wire  _T_1661 = io_multiplicand[0] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1664 = io_multiplicand[1] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1667 = io_multiplicand[2] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1670 = io_multiplicand[3] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1673 = io_multiplicand[4] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1676 = io_multiplicand[5] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1679 = io_multiplicand[6] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1682 = io_multiplicand[7] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1685 = io_multiplicand[8] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1688 = io_multiplicand[9] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1691 = io_multiplicand[10] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1694 = io_multiplicand[11] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1697 = io_multiplicand[12] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1700 = io_multiplicand[13] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1703 = io_multiplicand[14] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1706 = io_multiplicand[15] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1709 = io_multiplicand[16] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1712 = io_multiplicand[17] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1715 = io_multiplicand[18] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1718 = io_multiplicand[19] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1721 = io_multiplicand[20] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1724 = io_multiplicand[21] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1727 = io_multiplicand[22] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1730 = io_multiplicand[23] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1733 = io_multiplicand[24] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1736 = io_multiplicand[25] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1739 = io_multiplicand[26] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1742 = io_multiplicand[27] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1745 = io_multiplicand[28] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1748 = io_multiplicand[29] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1751 = io_multiplicand[30] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1754 = io_multiplicand[31] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1757 = io_multiplicand[32] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1760 = io_multiplicand[33] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1763 = io_multiplicand[34] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1766 = io_multiplicand[35] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1769 = io_multiplicand[36] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1772 = io_multiplicand[37] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1775 = io_multiplicand[38] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1778 = io_multiplicand[39] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1781 = io_multiplicand[40] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1784 = io_multiplicand[41] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1787 = io_multiplicand[42] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1790 = io_multiplicand[43] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1793 = io_multiplicand[44] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1796 = io_multiplicand[45] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1799 = io_multiplicand[46] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1802 = io_multiplicand[47] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1805 = io_multiplicand[48] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1808 = io_multiplicand[49] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1811 = io_multiplicand[50] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1814 = io_multiplicand[51] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1817 = io_multiplicand[52] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1820 = io_multiplicand[53] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1823 = io_multiplicand[54] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1826 = io_multiplicand[55] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1829 = io_multiplicand[56] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1832 = io_multiplicand[57] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1835 = io_multiplicand[58] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1838 = io_multiplicand[59] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1841 = io_multiplicand[60] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1844 = io_multiplicand[61] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1847 = io_multiplicand[62] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_1850 = io_multiplicand[63] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1859 = {_T_1850,_T_1847,_T_1844,_T_1841,_T_1838,_T_1835,_T_1832,_T_1829,_T_1826,_T_1823}; // @[Cat.scala 29:58]
  wire [18:0] _T_1868 = {_T_1859,_T_1820,_T_1817,_T_1814,_T_1811,_T_1808,_T_1805,_T_1802,_T_1799,_T_1796}; // @[Cat.scala 29:58]
  wire [27:0] _T_1877 = {_T_1868,_T_1793,_T_1790,_T_1787,_T_1784,_T_1781,_T_1778,_T_1775,_T_1772,_T_1769}; // @[Cat.scala 29:58]
  wire [36:0] _T_1886 = {_T_1877,_T_1766,_T_1763,_T_1760,_T_1757,_T_1754,_T_1751,_T_1748,_T_1745,_T_1742}; // @[Cat.scala 29:58]
  wire [45:0] _T_1895 = {_T_1886,_T_1739,_T_1736,_T_1733,_T_1730,_T_1727,_T_1724,_T_1721,_T_1718,_T_1715}; // @[Cat.scala 29:58]
  wire [54:0] _T_1904 = {_T_1895,_T_1712,_T_1709,_T_1706,_T_1703,_T_1700,_T_1697,_T_1694,_T_1691,_T_1688}; // @[Cat.scala 29:58]
  wire [62:0] _T_1912 = {_T_1904,_T_1685,_T_1682,_T_1679,_T_1676,_T_1673,_T_1670,_T_1667,_T_1664}; // @[Cat.scala 29:58]
  wire  _T_1980 = io_multiplicand[0] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1983 = io_multiplicand[1] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1986 = io_multiplicand[2] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1989 = io_multiplicand[3] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1992 = io_multiplicand[4] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1995 = io_multiplicand[5] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_1998 = io_multiplicand[6] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2001 = io_multiplicand[7] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2004 = io_multiplicand[8] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2007 = io_multiplicand[9] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2010 = io_multiplicand[10] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2013 = io_multiplicand[11] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2016 = io_multiplicand[12] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2019 = io_multiplicand[13] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2022 = io_multiplicand[14] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2025 = io_multiplicand[15] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2028 = io_multiplicand[16] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2031 = io_multiplicand[17] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2034 = io_multiplicand[18] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2037 = io_multiplicand[19] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2040 = io_multiplicand[20] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2043 = io_multiplicand[21] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2046 = io_multiplicand[22] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2049 = io_multiplicand[23] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2052 = io_multiplicand[24] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2055 = io_multiplicand[25] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2058 = io_multiplicand[26] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2061 = io_multiplicand[27] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2064 = io_multiplicand[28] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2067 = io_multiplicand[29] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2070 = io_multiplicand[30] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2073 = io_multiplicand[31] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2076 = io_multiplicand[32] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2079 = io_multiplicand[33] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2082 = io_multiplicand[34] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2085 = io_multiplicand[35] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2088 = io_multiplicand[36] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2091 = io_multiplicand[37] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2094 = io_multiplicand[38] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2097 = io_multiplicand[39] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2100 = io_multiplicand[40] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2103 = io_multiplicand[41] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2106 = io_multiplicand[42] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2109 = io_multiplicand[43] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2112 = io_multiplicand[44] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2115 = io_multiplicand[45] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2118 = io_multiplicand[46] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2121 = io_multiplicand[47] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2124 = io_multiplicand[48] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2127 = io_multiplicand[49] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2130 = io_multiplicand[50] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2133 = io_multiplicand[51] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2136 = io_multiplicand[52] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2139 = io_multiplicand[53] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2142 = io_multiplicand[54] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2145 = io_multiplicand[55] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2148 = io_multiplicand[56] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2151 = io_multiplicand[57] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2154 = io_multiplicand[58] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2157 = io_multiplicand[59] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2160 = io_multiplicand[60] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2163 = io_multiplicand[61] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2166 = io_multiplicand[62] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_2169 = io_multiplicand[63] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire [9:0] _T_2178 = {_T_2169,_T_2166,_T_2163,_T_2160,_T_2157,_T_2154,_T_2151,_T_2148,_T_2145,_T_2142}; // @[Cat.scala 29:58]
  wire [18:0] _T_2187 = {_T_2178,_T_2139,_T_2136,_T_2133,_T_2130,_T_2127,_T_2124,_T_2121,_T_2118,_T_2115}; // @[Cat.scala 29:58]
  wire [27:0] _T_2196 = {_T_2187,_T_2112,_T_2109,_T_2106,_T_2103,_T_2100,_T_2097,_T_2094,_T_2091,_T_2088}; // @[Cat.scala 29:58]
  wire [36:0] _T_2205 = {_T_2196,_T_2085,_T_2082,_T_2079,_T_2076,_T_2073,_T_2070,_T_2067,_T_2064,_T_2061}; // @[Cat.scala 29:58]
  wire [45:0] _T_2214 = {_T_2205,_T_2058,_T_2055,_T_2052,_T_2049,_T_2046,_T_2043,_T_2040,_T_2037,_T_2034}; // @[Cat.scala 29:58]
  wire [54:0] _T_2223 = {_T_2214,_T_2031,_T_2028,_T_2025,_T_2022,_T_2019,_T_2016,_T_2013,_T_2010,_T_2007}; // @[Cat.scala 29:58]
  wire [62:0] _T_2231 = {_T_2223,_T_2004,_T_2001,_T_1998,_T_1995,_T_1992,_T_1989,_T_1986,_T_1983}; // @[Cat.scala 29:58]
  wire  _T_2299 = io_multiplicand[0] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2302 = io_multiplicand[1] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2305 = io_multiplicand[2] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2308 = io_multiplicand[3] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2311 = io_multiplicand[4] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2314 = io_multiplicand[5] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2317 = io_multiplicand[6] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2320 = io_multiplicand[7] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2323 = io_multiplicand[8] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2326 = io_multiplicand[9] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2329 = io_multiplicand[10] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2332 = io_multiplicand[11] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2335 = io_multiplicand[12] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2338 = io_multiplicand[13] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2341 = io_multiplicand[14] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2344 = io_multiplicand[15] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2347 = io_multiplicand[16] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2350 = io_multiplicand[17] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2353 = io_multiplicand[18] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2356 = io_multiplicand[19] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2359 = io_multiplicand[20] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2362 = io_multiplicand[21] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2365 = io_multiplicand[22] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2368 = io_multiplicand[23] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2371 = io_multiplicand[24] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2374 = io_multiplicand[25] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2377 = io_multiplicand[26] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2380 = io_multiplicand[27] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2383 = io_multiplicand[28] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2386 = io_multiplicand[29] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2389 = io_multiplicand[30] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2392 = io_multiplicand[31] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2395 = io_multiplicand[32] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2398 = io_multiplicand[33] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2401 = io_multiplicand[34] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2404 = io_multiplicand[35] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2407 = io_multiplicand[36] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2410 = io_multiplicand[37] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2413 = io_multiplicand[38] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2416 = io_multiplicand[39] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2419 = io_multiplicand[40] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2422 = io_multiplicand[41] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2425 = io_multiplicand[42] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2428 = io_multiplicand[43] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2431 = io_multiplicand[44] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2434 = io_multiplicand[45] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2437 = io_multiplicand[46] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2440 = io_multiplicand[47] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2443 = io_multiplicand[48] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2446 = io_multiplicand[49] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2449 = io_multiplicand[50] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2452 = io_multiplicand[51] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2455 = io_multiplicand[52] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2458 = io_multiplicand[53] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2461 = io_multiplicand[54] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2464 = io_multiplicand[55] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2467 = io_multiplicand[56] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2470 = io_multiplicand[57] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2473 = io_multiplicand[58] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2476 = io_multiplicand[59] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2479 = io_multiplicand[60] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2482 = io_multiplicand[61] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2485 = io_multiplicand[62] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_2488 = io_multiplicand[63] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire [9:0] _T_2497 = {_T_2488,_T_2485,_T_2482,_T_2479,_T_2476,_T_2473,_T_2470,_T_2467,_T_2464,_T_2461}; // @[Cat.scala 29:58]
  wire [18:0] _T_2506 = {_T_2497,_T_2458,_T_2455,_T_2452,_T_2449,_T_2446,_T_2443,_T_2440,_T_2437,_T_2434}; // @[Cat.scala 29:58]
  wire [27:0] _T_2515 = {_T_2506,_T_2431,_T_2428,_T_2425,_T_2422,_T_2419,_T_2416,_T_2413,_T_2410,_T_2407}; // @[Cat.scala 29:58]
  wire [36:0] _T_2524 = {_T_2515,_T_2404,_T_2401,_T_2398,_T_2395,_T_2392,_T_2389,_T_2386,_T_2383,_T_2380}; // @[Cat.scala 29:58]
  wire [45:0] _T_2533 = {_T_2524,_T_2377,_T_2374,_T_2371,_T_2368,_T_2365,_T_2362,_T_2359,_T_2356,_T_2353}; // @[Cat.scala 29:58]
  wire [54:0] _T_2542 = {_T_2533,_T_2350,_T_2347,_T_2344,_T_2341,_T_2338,_T_2335,_T_2332,_T_2329,_T_2326}; // @[Cat.scala 29:58]
  wire [62:0] _T_2550 = {_T_2542,_T_2323,_T_2320,_T_2317,_T_2314,_T_2311,_T_2308,_T_2305,_T_2302}; // @[Cat.scala 29:58]
  wire  _T_2618 = io_multiplicand[0] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2621 = io_multiplicand[1] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2624 = io_multiplicand[2] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2627 = io_multiplicand[3] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2630 = io_multiplicand[4] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2633 = io_multiplicand[5] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2636 = io_multiplicand[6] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2639 = io_multiplicand[7] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2642 = io_multiplicand[8] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2645 = io_multiplicand[9] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2648 = io_multiplicand[10] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2651 = io_multiplicand[11] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2654 = io_multiplicand[12] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2657 = io_multiplicand[13] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2660 = io_multiplicand[14] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2663 = io_multiplicand[15] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2666 = io_multiplicand[16] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2669 = io_multiplicand[17] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2672 = io_multiplicand[18] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2675 = io_multiplicand[19] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2678 = io_multiplicand[20] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2681 = io_multiplicand[21] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2684 = io_multiplicand[22] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2687 = io_multiplicand[23] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2690 = io_multiplicand[24] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2693 = io_multiplicand[25] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2696 = io_multiplicand[26] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2699 = io_multiplicand[27] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2702 = io_multiplicand[28] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2705 = io_multiplicand[29] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2708 = io_multiplicand[30] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2711 = io_multiplicand[31] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2714 = io_multiplicand[32] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2717 = io_multiplicand[33] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2720 = io_multiplicand[34] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2723 = io_multiplicand[35] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2726 = io_multiplicand[36] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2729 = io_multiplicand[37] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2732 = io_multiplicand[38] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2735 = io_multiplicand[39] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2738 = io_multiplicand[40] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2741 = io_multiplicand[41] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2744 = io_multiplicand[42] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2747 = io_multiplicand[43] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2750 = io_multiplicand[44] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2753 = io_multiplicand[45] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2756 = io_multiplicand[46] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2759 = io_multiplicand[47] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2762 = io_multiplicand[48] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2765 = io_multiplicand[49] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2768 = io_multiplicand[50] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2771 = io_multiplicand[51] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2774 = io_multiplicand[52] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2777 = io_multiplicand[53] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2780 = io_multiplicand[54] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2783 = io_multiplicand[55] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2786 = io_multiplicand[56] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2789 = io_multiplicand[57] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2792 = io_multiplicand[58] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2795 = io_multiplicand[59] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2798 = io_multiplicand[60] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2801 = io_multiplicand[61] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2804 = io_multiplicand[62] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_2807 = io_multiplicand[63] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire [9:0] _T_2816 = {_T_2807,_T_2804,_T_2801,_T_2798,_T_2795,_T_2792,_T_2789,_T_2786,_T_2783,_T_2780}; // @[Cat.scala 29:58]
  wire [18:0] _T_2825 = {_T_2816,_T_2777,_T_2774,_T_2771,_T_2768,_T_2765,_T_2762,_T_2759,_T_2756,_T_2753}; // @[Cat.scala 29:58]
  wire [27:0] _T_2834 = {_T_2825,_T_2750,_T_2747,_T_2744,_T_2741,_T_2738,_T_2735,_T_2732,_T_2729,_T_2726}; // @[Cat.scala 29:58]
  wire [36:0] _T_2843 = {_T_2834,_T_2723,_T_2720,_T_2717,_T_2714,_T_2711,_T_2708,_T_2705,_T_2702,_T_2699}; // @[Cat.scala 29:58]
  wire [45:0] _T_2852 = {_T_2843,_T_2696,_T_2693,_T_2690,_T_2687,_T_2684,_T_2681,_T_2678,_T_2675,_T_2672}; // @[Cat.scala 29:58]
  wire [54:0] _T_2861 = {_T_2852,_T_2669,_T_2666,_T_2663,_T_2660,_T_2657,_T_2654,_T_2651,_T_2648,_T_2645}; // @[Cat.scala 29:58]
  wire [62:0] _T_2869 = {_T_2861,_T_2642,_T_2639,_T_2636,_T_2633,_T_2630,_T_2627,_T_2624,_T_2621}; // @[Cat.scala 29:58]
  wire  _T_2937 = io_multiplicand[0] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2940 = io_multiplicand[1] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2943 = io_multiplicand[2] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2946 = io_multiplicand[3] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2949 = io_multiplicand[4] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2952 = io_multiplicand[5] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2955 = io_multiplicand[6] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2958 = io_multiplicand[7] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2961 = io_multiplicand[8] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2964 = io_multiplicand[9] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2967 = io_multiplicand[10] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2970 = io_multiplicand[11] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2973 = io_multiplicand[12] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2976 = io_multiplicand[13] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2979 = io_multiplicand[14] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2982 = io_multiplicand[15] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2985 = io_multiplicand[16] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2988 = io_multiplicand[17] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2991 = io_multiplicand[18] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2994 = io_multiplicand[19] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_2997 = io_multiplicand[20] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3000 = io_multiplicand[21] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3003 = io_multiplicand[22] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3006 = io_multiplicand[23] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3009 = io_multiplicand[24] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3012 = io_multiplicand[25] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3015 = io_multiplicand[26] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3018 = io_multiplicand[27] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3021 = io_multiplicand[28] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3024 = io_multiplicand[29] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3027 = io_multiplicand[30] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3030 = io_multiplicand[31] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3033 = io_multiplicand[32] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3036 = io_multiplicand[33] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3039 = io_multiplicand[34] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3042 = io_multiplicand[35] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3045 = io_multiplicand[36] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3048 = io_multiplicand[37] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3051 = io_multiplicand[38] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3054 = io_multiplicand[39] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3057 = io_multiplicand[40] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3060 = io_multiplicand[41] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3063 = io_multiplicand[42] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3066 = io_multiplicand[43] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3069 = io_multiplicand[44] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3072 = io_multiplicand[45] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3075 = io_multiplicand[46] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3078 = io_multiplicand[47] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3081 = io_multiplicand[48] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3084 = io_multiplicand[49] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3087 = io_multiplicand[50] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3090 = io_multiplicand[51] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3093 = io_multiplicand[52] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3096 = io_multiplicand[53] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3099 = io_multiplicand[54] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3102 = io_multiplicand[55] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3105 = io_multiplicand[56] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3108 = io_multiplicand[57] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3111 = io_multiplicand[58] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3114 = io_multiplicand[59] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3117 = io_multiplicand[60] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3120 = io_multiplicand[61] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3123 = io_multiplicand[62] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_3126 = io_multiplicand[63] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire [9:0] _T_3135 = {_T_3126,_T_3123,_T_3120,_T_3117,_T_3114,_T_3111,_T_3108,_T_3105,_T_3102,_T_3099}; // @[Cat.scala 29:58]
  wire [18:0] _T_3144 = {_T_3135,_T_3096,_T_3093,_T_3090,_T_3087,_T_3084,_T_3081,_T_3078,_T_3075,_T_3072}; // @[Cat.scala 29:58]
  wire [27:0] _T_3153 = {_T_3144,_T_3069,_T_3066,_T_3063,_T_3060,_T_3057,_T_3054,_T_3051,_T_3048,_T_3045}; // @[Cat.scala 29:58]
  wire [36:0] _T_3162 = {_T_3153,_T_3042,_T_3039,_T_3036,_T_3033,_T_3030,_T_3027,_T_3024,_T_3021,_T_3018}; // @[Cat.scala 29:58]
  wire [45:0] _T_3171 = {_T_3162,_T_3015,_T_3012,_T_3009,_T_3006,_T_3003,_T_3000,_T_2997,_T_2994,_T_2991}; // @[Cat.scala 29:58]
  wire [54:0] _T_3180 = {_T_3171,_T_2988,_T_2985,_T_2982,_T_2979,_T_2976,_T_2973,_T_2970,_T_2967,_T_2964}; // @[Cat.scala 29:58]
  wire [62:0] _T_3188 = {_T_3180,_T_2961,_T_2958,_T_2955,_T_2952,_T_2949,_T_2946,_T_2943,_T_2940}; // @[Cat.scala 29:58]
  wire  _T_3256 = io_multiplicand[0] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3259 = io_multiplicand[1] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3262 = io_multiplicand[2] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3265 = io_multiplicand[3] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3268 = io_multiplicand[4] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3271 = io_multiplicand[5] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3274 = io_multiplicand[6] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3277 = io_multiplicand[7] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3280 = io_multiplicand[8] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3283 = io_multiplicand[9] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3286 = io_multiplicand[10] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3289 = io_multiplicand[11] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3292 = io_multiplicand[12] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3295 = io_multiplicand[13] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3298 = io_multiplicand[14] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3301 = io_multiplicand[15] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3304 = io_multiplicand[16] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3307 = io_multiplicand[17] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3310 = io_multiplicand[18] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3313 = io_multiplicand[19] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3316 = io_multiplicand[20] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3319 = io_multiplicand[21] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3322 = io_multiplicand[22] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3325 = io_multiplicand[23] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3328 = io_multiplicand[24] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3331 = io_multiplicand[25] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3334 = io_multiplicand[26] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3337 = io_multiplicand[27] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3340 = io_multiplicand[28] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3343 = io_multiplicand[29] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3346 = io_multiplicand[30] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3349 = io_multiplicand[31] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3352 = io_multiplicand[32] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3355 = io_multiplicand[33] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3358 = io_multiplicand[34] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3361 = io_multiplicand[35] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3364 = io_multiplicand[36] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3367 = io_multiplicand[37] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3370 = io_multiplicand[38] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3373 = io_multiplicand[39] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3376 = io_multiplicand[40] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3379 = io_multiplicand[41] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3382 = io_multiplicand[42] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3385 = io_multiplicand[43] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3388 = io_multiplicand[44] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3391 = io_multiplicand[45] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3394 = io_multiplicand[46] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3397 = io_multiplicand[47] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3400 = io_multiplicand[48] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3403 = io_multiplicand[49] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3406 = io_multiplicand[50] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3409 = io_multiplicand[51] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3412 = io_multiplicand[52] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3415 = io_multiplicand[53] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3418 = io_multiplicand[54] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3421 = io_multiplicand[55] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3424 = io_multiplicand[56] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3427 = io_multiplicand[57] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3430 = io_multiplicand[58] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3433 = io_multiplicand[59] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3436 = io_multiplicand[60] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3439 = io_multiplicand[61] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3442 = io_multiplicand[62] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_3445 = io_multiplicand[63] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire [9:0] _T_3454 = {_T_3445,_T_3442,_T_3439,_T_3436,_T_3433,_T_3430,_T_3427,_T_3424,_T_3421,_T_3418}; // @[Cat.scala 29:58]
  wire [18:0] _T_3463 = {_T_3454,_T_3415,_T_3412,_T_3409,_T_3406,_T_3403,_T_3400,_T_3397,_T_3394,_T_3391}; // @[Cat.scala 29:58]
  wire [27:0] _T_3472 = {_T_3463,_T_3388,_T_3385,_T_3382,_T_3379,_T_3376,_T_3373,_T_3370,_T_3367,_T_3364}; // @[Cat.scala 29:58]
  wire [36:0] _T_3481 = {_T_3472,_T_3361,_T_3358,_T_3355,_T_3352,_T_3349,_T_3346,_T_3343,_T_3340,_T_3337}; // @[Cat.scala 29:58]
  wire [45:0] _T_3490 = {_T_3481,_T_3334,_T_3331,_T_3328,_T_3325,_T_3322,_T_3319,_T_3316,_T_3313,_T_3310}; // @[Cat.scala 29:58]
  wire [54:0] _T_3499 = {_T_3490,_T_3307,_T_3304,_T_3301,_T_3298,_T_3295,_T_3292,_T_3289,_T_3286,_T_3283}; // @[Cat.scala 29:58]
  wire [62:0] _T_3507 = {_T_3499,_T_3280,_T_3277,_T_3274,_T_3271,_T_3268,_T_3265,_T_3262,_T_3259}; // @[Cat.scala 29:58]
  wire  _T_3575 = io_multiplicand[0] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3578 = io_multiplicand[1] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3581 = io_multiplicand[2] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3584 = io_multiplicand[3] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3587 = io_multiplicand[4] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3590 = io_multiplicand[5] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3593 = io_multiplicand[6] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3596 = io_multiplicand[7] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3599 = io_multiplicand[8] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3602 = io_multiplicand[9] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3605 = io_multiplicand[10] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3608 = io_multiplicand[11] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3611 = io_multiplicand[12] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3614 = io_multiplicand[13] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3617 = io_multiplicand[14] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3620 = io_multiplicand[15] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3623 = io_multiplicand[16] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3626 = io_multiplicand[17] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3629 = io_multiplicand[18] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3632 = io_multiplicand[19] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3635 = io_multiplicand[20] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3638 = io_multiplicand[21] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3641 = io_multiplicand[22] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3644 = io_multiplicand[23] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3647 = io_multiplicand[24] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3650 = io_multiplicand[25] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3653 = io_multiplicand[26] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3656 = io_multiplicand[27] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3659 = io_multiplicand[28] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3662 = io_multiplicand[29] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3665 = io_multiplicand[30] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3668 = io_multiplicand[31] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3671 = io_multiplicand[32] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3674 = io_multiplicand[33] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3677 = io_multiplicand[34] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3680 = io_multiplicand[35] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3683 = io_multiplicand[36] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3686 = io_multiplicand[37] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3689 = io_multiplicand[38] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3692 = io_multiplicand[39] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3695 = io_multiplicand[40] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3698 = io_multiplicand[41] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3701 = io_multiplicand[42] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3704 = io_multiplicand[43] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3707 = io_multiplicand[44] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3710 = io_multiplicand[45] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3713 = io_multiplicand[46] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3716 = io_multiplicand[47] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3719 = io_multiplicand[48] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3722 = io_multiplicand[49] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3725 = io_multiplicand[50] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3728 = io_multiplicand[51] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3731 = io_multiplicand[52] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3734 = io_multiplicand[53] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3737 = io_multiplicand[54] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3740 = io_multiplicand[55] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3743 = io_multiplicand[56] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3746 = io_multiplicand[57] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3749 = io_multiplicand[58] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3752 = io_multiplicand[59] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3755 = io_multiplicand[60] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3758 = io_multiplicand[61] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3761 = io_multiplicand[62] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_3764 = io_multiplicand[63] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire [9:0] _T_3773 = {_T_3764,_T_3761,_T_3758,_T_3755,_T_3752,_T_3749,_T_3746,_T_3743,_T_3740,_T_3737}; // @[Cat.scala 29:58]
  wire [18:0] _T_3782 = {_T_3773,_T_3734,_T_3731,_T_3728,_T_3725,_T_3722,_T_3719,_T_3716,_T_3713,_T_3710}; // @[Cat.scala 29:58]
  wire [27:0] _T_3791 = {_T_3782,_T_3707,_T_3704,_T_3701,_T_3698,_T_3695,_T_3692,_T_3689,_T_3686,_T_3683}; // @[Cat.scala 29:58]
  wire [36:0] _T_3800 = {_T_3791,_T_3680,_T_3677,_T_3674,_T_3671,_T_3668,_T_3665,_T_3662,_T_3659,_T_3656}; // @[Cat.scala 29:58]
  wire [45:0] _T_3809 = {_T_3800,_T_3653,_T_3650,_T_3647,_T_3644,_T_3641,_T_3638,_T_3635,_T_3632,_T_3629}; // @[Cat.scala 29:58]
  wire [54:0] _T_3818 = {_T_3809,_T_3626,_T_3623,_T_3620,_T_3617,_T_3614,_T_3611,_T_3608,_T_3605,_T_3602}; // @[Cat.scala 29:58]
  wire [62:0] _T_3826 = {_T_3818,_T_3599,_T_3596,_T_3593,_T_3590,_T_3587,_T_3584,_T_3581,_T_3578}; // @[Cat.scala 29:58]
  wire  _T_3894 = io_multiplicand[0] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3897 = io_multiplicand[1] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3900 = io_multiplicand[2] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3903 = io_multiplicand[3] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3906 = io_multiplicand[4] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3909 = io_multiplicand[5] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3912 = io_multiplicand[6] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3915 = io_multiplicand[7] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3918 = io_multiplicand[8] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3921 = io_multiplicand[9] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3924 = io_multiplicand[10] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3927 = io_multiplicand[11] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3930 = io_multiplicand[12] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3933 = io_multiplicand[13] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3936 = io_multiplicand[14] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3939 = io_multiplicand[15] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3942 = io_multiplicand[16] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3945 = io_multiplicand[17] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3948 = io_multiplicand[18] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3951 = io_multiplicand[19] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3954 = io_multiplicand[20] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3957 = io_multiplicand[21] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3960 = io_multiplicand[22] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3963 = io_multiplicand[23] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3966 = io_multiplicand[24] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3969 = io_multiplicand[25] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3972 = io_multiplicand[26] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3975 = io_multiplicand[27] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3978 = io_multiplicand[28] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3981 = io_multiplicand[29] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3984 = io_multiplicand[30] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3987 = io_multiplicand[31] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3990 = io_multiplicand[32] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3993 = io_multiplicand[33] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3996 = io_multiplicand[34] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_3999 = io_multiplicand[35] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4002 = io_multiplicand[36] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4005 = io_multiplicand[37] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4008 = io_multiplicand[38] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4011 = io_multiplicand[39] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4014 = io_multiplicand[40] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4017 = io_multiplicand[41] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4020 = io_multiplicand[42] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4023 = io_multiplicand[43] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4026 = io_multiplicand[44] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4029 = io_multiplicand[45] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4032 = io_multiplicand[46] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4035 = io_multiplicand[47] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4038 = io_multiplicand[48] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4041 = io_multiplicand[49] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4044 = io_multiplicand[50] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4047 = io_multiplicand[51] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4050 = io_multiplicand[52] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4053 = io_multiplicand[53] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4056 = io_multiplicand[54] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4059 = io_multiplicand[55] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4062 = io_multiplicand[56] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4065 = io_multiplicand[57] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4068 = io_multiplicand[58] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4071 = io_multiplicand[59] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4074 = io_multiplicand[60] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4077 = io_multiplicand[61] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4080 = io_multiplicand[62] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_4083 = io_multiplicand[63] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire [9:0] _T_4092 = {_T_4083,_T_4080,_T_4077,_T_4074,_T_4071,_T_4068,_T_4065,_T_4062,_T_4059,_T_4056}; // @[Cat.scala 29:58]
  wire [18:0] _T_4101 = {_T_4092,_T_4053,_T_4050,_T_4047,_T_4044,_T_4041,_T_4038,_T_4035,_T_4032,_T_4029}; // @[Cat.scala 29:58]
  wire [27:0] _T_4110 = {_T_4101,_T_4026,_T_4023,_T_4020,_T_4017,_T_4014,_T_4011,_T_4008,_T_4005,_T_4002}; // @[Cat.scala 29:58]
  wire [36:0] _T_4119 = {_T_4110,_T_3999,_T_3996,_T_3993,_T_3990,_T_3987,_T_3984,_T_3981,_T_3978,_T_3975}; // @[Cat.scala 29:58]
  wire [45:0] _T_4128 = {_T_4119,_T_3972,_T_3969,_T_3966,_T_3963,_T_3960,_T_3957,_T_3954,_T_3951,_T_3948}; // @[Cat.scala 29:58]
  wire [54:0] _T_4137 = {_T_4128,_T_3945,_T_3942,_T_3939,_T_3936,_T_3933,_T_3930,_T_3927,_T_3924,_T_3921}; // @[Cat.scala 29:58]
  wire [62:0] _T_4145 = {_T_4137,_T_3918,_T_3915,_T_3912,_T_3909,_T_3906,_T_3903,_T_3900,_T_3897}; // @[Cat.scala 29:58]
  wire  _T_4213 = io_multiplicand[0] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4216 = io_multiplicand[1] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4219 = io_multiplicand[2] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4222 = io_multiplicand[3] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4225 = io_multiplicand[4] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4228 = io_multiplicand[5] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4231 = io_multiplicand[6] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4234 = io_multiplicand[7] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4237 = io_multiplicand[8] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4240 = io_multiplicand[9] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4243 = io_multiplicand[10] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4246 = io_multiplicand[11] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4249 = io_multiplicand[12] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4252 = io_multiplicand[13] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4255 = io_multiplicand[14] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4258 = io_multiplicand[15] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4261 = io_multiplicand[16] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4264 = io_multiplicand[17] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4267 = io_multiplicand[18] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4270 = io_multiplicand[19] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4273 = io_multiplicand[20] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4276 = io_multiplicand[21] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4279 = io_multiplicand[22] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4282 = io_multiplicand[23] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4285 = io_multiplicand[24] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4288 = io_multiplicand[25] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4291 = io_multiplicand[26] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4294 = io_multiplicand[27] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4297 = io_multiplicand[28] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4300 = io_multiplicand[29] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4303 = io_multiplicand[30] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4306 = io_multiplicand[31] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4309 = io_multiplicand[32] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4312 = io_multiplicand[33] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4315 = io_multiplicand[34] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4318 = io_multiplicand[35] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4321 = io_multiplicand[36] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4324 = io_multiplicand[37] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4327 = io_multiplicand[38] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4330 = io_multiplicand[39] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4333 = io_multiplicand[40] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4336 = io_multiplicand[41] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4339 = io_multiplicand[42] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4342 = io_multiplicand[43] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4345 = io_multiplicand[44] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4348 = io_multiplicand[45] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4351 = io_multiplicand[46] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4354 = io_multiplicand[47] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4357 = io_multiplicand[48] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4360 = io_multiplicand[49] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4363 = io_multiplicand[50] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4366 = io_multiplicand[51] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4369 = io_multiplicand[52] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4372 = io_multiplicand[53] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4375 = io_multiplicand[54] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4378 = io_multiplicand[55] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4381 = io_multiplicand[56] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4384 = io_multiplicand[57] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4387 = io_multiplicand[58] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4390 = io_multiplicand[59] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4393 = io_multiplicand[60] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4396 = io_multiplicand[61] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4399 = io_multiplicand[62] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_4402 = io_multiplicand[63] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire [9:0] _T_4411 = {_T_4402,_T_4399,_T_4396,_T_4393,_T_4390,_T_4387,_T_4384,_T_4381,_T_4378,_T_4375}; // @[Cat.scala 29:58]
  wire [18:0] _T_4420 = {_T_4411,_T_4372,_T_4369,_T_4366,_T_4363,_T_4360,_T_4357,_T_4354,_T_4351,_T_4348}; // @[Cat.scala 29:58]
  wire [27:0] _T_4429 = {_T_4420,_T_4345,_T_4342,_T_4339,_T_4336,_T_4333,_T_4330,_T_4327,_T_4324,_T_4321}; // @[Cat.scala 29:58]
  wire [36:0] _T_4438 = {_T_4429,_T_4318,_T_4315,_T_4312,_T_4309,_T_4306,_T_4303,_T_4300,_T_4297,_T_4294}; // @[Cat.scala 29:58]
  wire [45:0] _T_4447 = {_T_4438,_T_4291,_T_4288,_T_4285,_T_4282,_T_4279,_T_4276,_T_4273,_T_4270,_T_4267}; // @[Cat.scala 29:58]
  wire [54:0] _T_4456 = {_T_4447,_T_4264,_T_4261,_T_4258,_T_4255,_T_4252,_T_4249,_T_4246,_T_4243,_T_4240}; // @[Cat.scala 29:58]
  wire [62:0] _T_4464 = {_T_4456,_T_4237,_T_4234,_T_4231,_T_4228,_T_4225,_T_4222,_T_4219,_T_4216}; // @[Cat.scala 29:58]
  wire  _T_4532 = io_multiplicand[0] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4535 = io_multiplicand[1] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4538 = io_multiplicand[2] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4541 = io_multiplicand[3] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4544 = io_multiplicand[4] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4547 = io_multiplicand[5] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4550 = io_multiplicand[6] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4553 = io_multiplicand[7] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4556 = io_multiplicand[8] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4559 = io_multiplicand[9] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4562 = io_multiplicand[10] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4565 = io_multiplicand[11] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4568 = io_multiplicand[12] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4571 = io_multiplicand[13] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4574 = io_multiplicand[14] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4577 = io_multiplicand[15] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4580 = io_multiplicand[16] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4583 = io_multiplicand[17] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4586 = io_multiplicand[18] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4589 = io_multiplicand[19] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4592 = io_multiplicand[20] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4595 = io_multiplicand[21] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4598 = io_multiplicand[22] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4601 = io_multiplicand[23] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4604 = io_multiplicand[24] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4607 = io_multiplicand[25] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4610 = io_multiplicand[26] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4613 = io_multiplicand[27] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4616 = io_multiplicand[28] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4619 = io_multiplicand[29] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4622 = io_multiplicand[30] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4625 = io_multiplicand[31] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4628 = io_multiplicand[32] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4631 = io_multiplicand[33] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4634 = io_multiplicand[34] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4637 = io_multiplicand[35] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4640 = io_multiplicand[36] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4643 = io_multiplicand[37] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4646 = io_multiplicand[38] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4649 = io_multiplicand[39] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4652 = io_multiplicand[40] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4655 = io_multiplicand[41] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4658 = io_multiplicand[42] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4661 = io_multiplicand[43] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4664 = io_multiplicand[44] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4667 = io_multiplicand[45] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4670 = io_multiplicand[46] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4673 = io_multiplicand[47] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4676 = io_multiplicand[48] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4679 = io_multiplicand[49] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4682 = io_multiplicand[50] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4685 = io_multiplicand[51] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4688 = io_multiplicand[52] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4691 = io_multiplicand[53] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4694 = io_multiplicand[54] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4697 = io_multiplicand[55] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4700 = io_multiplicand[56] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4703 = io_multiplicand[57] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4706 = io_multiplicand[58] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4709 = io_multiplicand[59] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4712 = io_multiplicand[60] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4715 = io_multiplicand[61] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4718 = io_multiplicand[62] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_4721 = io_multiplicand[63] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire [9:0] _T_4730 = {_T_4721,_T_4718,_T_4715,_T_4712,_T_4709,_T_4706,_T_4703,_T_4700,_T_4697,_T_4694}; // @[Cat.scala 29:58]
  wire [18:0] _T_4739 = {_T_4730,_T_4691,_T_4688,_T_4685,_T_4682,_T_4679,_T_4676,_T_4673,_T_4670,_T_4667}; // @[Cat.scala 29:58]
  wire [27:0] _T_4748 = {_T_4739,_T_4664,_T_4661,_T_4658,_T_4655,_T_4652,_T_4649,_T_4646,_T_4643,_T_4640}; // @[Cat.scala 29:58]
  wire [36:0] _T_4757 = {_T_4748,_T_4637,_T_4634,_T_4631,_T_4628,_T_4625,_T_4622,_T_4619,_T_4616,_T_4613}; // @[Cat.scala 29:58]
  wire [45:0] _T_4766 = {_T_4757,_T_4610,_T_4607,_T_4604,_T_4601,_T_4598,_T_4595,_T_4592,_T_4589,_T_4586}; // @[Cat.scala 29:58]
  wire [54:0] _T_4775 = {_T_4766,_T_4583,_T_4580,_T_4577,_T_4574,_T_4571,_T_4568,_T_4565,_T_4562,_T_4559}; // @[Cat.scala 29:58]
  wire [62:0] _T_4783 = {_T_4775,_T_4556,_T_4553,_T_4550,_T_4547,_T_4544,_T_4541,_T_4538,_T_4535}; // @[Cat.scala 29:58]
  wire  _T_4851 = io_multiplicand[0] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4854 = io_multiplicand[1] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4857 = io_multiplicand[2] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4860 = io_multiplicand[3] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4863 = io_multiplicand[4] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4866 = io_multiplicand[5] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4869 = io_multiplicand[6] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4872 = io_multiplicand[7] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4875 = io_multiplicand[8] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4878 = io_multiplicand[9] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4881 = io_multiplicand[10] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4884 = io_multiplicand[11] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4887 = io_multiplicand[12] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4890 = io_multiplicand[13] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4893 = io_multiplicand[14] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4896 = io_multiplicand[15] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4899 = io_multiplicand[16] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4902 = io_multiplicand[17] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4905 = io_multiplicand[18] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4908 = io_multiplicand[19] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4911 = io_multiplicand[20] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4914 = io_multiplicand[21] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4917 = io_multiplicand[22] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4920 = io_multiplicand[23] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4923 = io_multiplicand[24] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4926 = io_multiplicand[25] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4929 = io_multiplicand[26] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4932 = io_multiplicand[27] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4935 = io_multiplicand[28] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4938 = io_multiplicand[29] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4941 = io_multiplicand[30] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4944 = io_multiplicand[31] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4947 = io_multiplicand[32] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4950 = io_multiplicand[33] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4953 = io_multiplicand[34] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4956 = io_multiplicand[35] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4959 = io_multiplicand[36] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4962 = io_multiplicand[37] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4965 = io_multiplicand[38] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4968 = io_multiplicand[39] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4971 = io_multiplicand[40] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4974 = io_multiplicand[41] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4977 = io_multiplicand[42] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4980 = io_multiplicand[43] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4983 = io_multiplicand[44] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4986 = io_multiplicand[45] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4989 = io_multiplicand[46] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4992 = io_multiplicand[47] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4995 = io_multiplicand[48] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_4998 = io_multiplicand[49] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_5001 = io_multiplicand[50] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_5004 = io_multiplicand[51] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_5007 = io_multiplicand[52] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_5010 = io_multiplicand[53] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_5013 = io_multiplicand[54] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_5016 = io_multiplicand[55] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_5019 = io_multiplicand[56] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_5022 = io_multiplicand[57] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_5025 = io_multiplicand[58] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_5028 = io_multiplicand[59] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_5031 = io_multiplicand[60] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_5034 = io_multiplicand[61] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_5037 = io_multiplicand[62] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_5040 = io_multiplicand[63] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire [9:0] _T_5049 = {_T_5040,_T_5037,_T_5034,_T_5031,_T_5028,_T_5025,_T_5022,_T_5019,_T_5016,_T_5013}; // @[Cat.scala 29:58]
  wire [18:0] _T_5058 = {_T_5049,_T_5010,_T_5007,_T_5004,_T_5001,_T_4998,_T_4995,_T_4992,_T_4989,_T_4986}; // @[Cat.scala 29:58]
  wire [27:0] _T_5067 = {_T_5058,_T_4983,_T_4980,_T_4977,_T_4974,_T_4971,_T_4968,_T_4965,_T_4962,_T_4959}; // @[Cat.scala 29:58]
  wire [36:0] _T_5076 = {_T_5067,_T_4956,_T_4953,_T_4950,_T_4947,_T_4944,_T_4941,_T_4938,_T_4935,_T_4932}; // @[Cat.scala 29:58]
  wire [45:0] _T_5085 = {_T_5076,_T_4929,_T_4926,_T_4923,_T_4920,_T_4917,_T_4914,_T_4911,_T_4908,_T_4905}; // @[Cat.scala 29:58]
  wire [54:0] _T_5094 = {_T_5085,_T_4902,_T_4899,_T_4896,_T_4893,_T_4890,_T_4887,_T_4884,_T_4881,_T_4878}; // @[Cat.scala 29:58]
  wire [62:0] _T_5102 = {_T_5094,_T_4875,_T_4872,_T_4869,_T_4866,_T_4863,_T_4860,_T_4857,_T_4854}; // @[Cat.scala 29:58]
  wire  _T_5170 = io_multiplicand[0] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5173 = io_multiplicand[1] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5176 = io_multiplicand[2] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5179 = io_multiplicand[3] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5182 = io_multiplicand[4] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5185 = io_multiplicand[5] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5188 = io_multiplicand[6] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5191 = io_multiplicand[7] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5194 = io_multiplicand[8] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5197 = io_multiplicand[9] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5200 = io_multiplicand[10] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5203 = io_multiplicand[11] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5206 = io_multiplicand[12] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5209 = io_multiplicand[13] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5212 = io_multiplicand[14] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5215 = io_multiplicand[15] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5218 = io_multiplicand[16] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5221 = io_multiplicand[17] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5224 = io_multiplicand[18] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5227 = io_multiplicand[19] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5230 = io_multiplicand[20] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5233 = io_multiplicand[21] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5236 = io_multiplicand[22] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5239 = io_multiplicand[23] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5242 = io_multiplicand[24] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5245 = io_multiplicand[25] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5248 = io_multiplicand[26] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5251 = io_multiplicand[27] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5254 = io_multiplicand[28] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5257 = io_multiplicand[29] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5260 = io_multiplicand[30] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5263 = io_multiplicand[31] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5266 = io_multiplicand[32] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5269 = io_multiplicand[33] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5272 = io_multiplicand[34] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5275 = io_multiplicand[35] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5278 = io_multiplicand[36] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5281 = io_multiplicand[37] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5284 = io_multiplicand[38] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5287 = io_multiplicand[39] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5290 = io_multiplicand[40] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5293 = io_multiplicand[41] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5296 = io_multiplicand[42] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5299 = io_multiplicand[43] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5302 = io_multiplicand[44] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5305 = io_multiplicand[45] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5308 = io_multiplicand[46] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5311 = io_multiplicand[47] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5314 = io_multiplicand[48] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5317 = io_multiplicand[49] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5320 = io_multiplicand[50] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5323 = io_multiplicand[51] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5326 = io_multiplicand[52] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5329 = io_multiplicand[53] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5332 = io_multiplicand[54] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5335 = io_multiplicand[55] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5338 = io_multiplicand[56] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5341 = io_multiplicand[57] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5344 = io_multiplicand[58] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5347 = io_multiplicand[59] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5350 = io_multiplicand[60] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5353 = io_multiplicand[61] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5356 = io_multiplicand[62] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire  _T_5359 = io_multiplicand[63] & io_multiplier[16]; // @[partialprod.scala 16:36]
  wire [9:0] _T_5368 = {_T_5359,_T_5356,_T_5353,_T_5350,_T_5347,_T_5344,_T_5341,_T_5338,_T_5335,_T_5332}; // @[Cat.scala 29:58]
  wire [18:0] _T_5377 = {_T_5368,_T_5329,_T_5326,_T_5323,_T_5320,_T_5317,_T_5314,_T_5311,_T_5308,_T_5305}; // @[Cat.scala 29:58]
  wire [27:0] _T_5386 = {_T_5377,_T_5302,_T_5299,_T_5296,_T_5293,_T_5290,_T_5287,_T_5284,_T_5281,_T_5278}; // @[Cat.scala 29:58]
  wire [36:0] _T_5395 = {_T_5386,_T_5275,_T_5272,_T_5269,_T_5266,_T_5263,_T_5260,_T_5257,_T_5254,_T_5251}; // @[Cat.scala 29:58]
  wire [45:0] _T_5404 = {_T_5395,_T_5248,_T_5245,_T_5242,_T_5239,_T_5236,_T_5233,_T_5230,_T_5227,_T_5224}; // @[Cat.scala 29:58]
  wire [54:0] _T_5413 = {_T_5404,_T_5221,_T_5218,_T_5215,_T_5212,_T_5209,_T_5206,_T_5203,_T_5200,_T_5197}; // @[Cat.scala 29:58]
  wire [62:0] _T_5421 = {_T_5413,_T_5194,_T_5191,_T_5188,_T_5185,_T_5182,_T_5179,_T_5176,_T_5173}; // @[Cat.scala 29:58]
  wire  _T_5489 = io_multiplicand[0] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5492 = io_multiplicand[1] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5495 = io_multiplicand[2] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5498 = io_multiplicand[3] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5501 = io_multiplicand[4] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5504 = io_multiplicand[5] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5507 = io_multiplicand[6] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5510 = io_multiplicand[7] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5513 = io_multiplicand[8] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5516 = io_multiplicand[9] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5519 = io_multiplicand[10] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5522 = io_multiplicand[11] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5525 = io_multiplicand[12] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5528 = io_multiplicand[13] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5531 = io_multiplicand[14] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5534 = io_multiplicand[15] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5537 = io_multiplicand[16] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5540 = io_multiplicand[17] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5543 = io_multiplicand[18] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5546 = io_multiplicand[19] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5549 = io_multiplicand[20] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5552 = io_multiplicand[21] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5555 = io_multiplicand[22] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5558 = io_multiplicand[23] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5561 = io_multiplicand[24] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5564 = io_multiplicand[25] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5567 = io_multiplicand[26] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5570 = io_multiplicand[27] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5573 = io_multiplicand[28] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5576 = io_multiplicand[29] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5579 = io_multiplicand[30] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5582 = io_multiplicand[31] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5585 = io_multiplicand[32] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5588 = io_multiplicand[33] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5591 = io_multiplicand[34] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5594 = io_multiplicand[35] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5597 = io_multiplicand[36] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5600 = io_multiplicand[37] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5603 = io_multiplicand[38] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5606 = io_multiplicand[39] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5609 = io_multiplicand[40] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5612 = io_multiplicand[41] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5615 = io_multiplicand[42] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5618 = io_multiplicand[43] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5621 = io_multiplicand[44] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5624 = io_multiplicand[45] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5627 = io_multiplicand[46] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5630 = io_multiplicand[47] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5633 = io_multiplicand[48] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5636 = io_multiplicand[49] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5639 = io_multiplicand[50] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5642 = io_multiplicand[51] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5645 = io_multiplicand[52] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5648 = io_multiplicand[53] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5651 = io_multiplicand[54] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5654 = io_multiplicand[55] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5657 = io_multiplicand[56] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5660 = io_multiplicand[57] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5663 = io_multiplicand[58] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5666 = io_multiplicand[59] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5669 = io_multiplicand[60] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5672 = io_multiplicand[61] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5675 = io_multiplicand[62] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire  _T_5678 = io_multiplicand[63] & io_multiplier[17]; // @[partialprod.scala 16:36]
  wire [9:0] _T_5687 = {_T_5678,_T_5675,_T_5672,_T_5669,_T_5666,_T_5663,_T_5660,_T_5657,_T_5654,_T_5651}; // @[Cat.scala 29:58]
  wire [18:0] _T_5696 = {_T_5687,_T_5648,_T_5645,_T_5642,_T_5639,_T_5636,_T_5633,_T_5630,_T_5627,_T_5624}; // @[Cat.scala 29:58]
  wire [27:0] _T_5705 = {_T_5696,_T_5621,_T_5618,_T_5615,_T_5612,_T_5609,_T_5606,_T_5603,_T_5600,_T_5597}; // @[Cat.scala 29:58]
  wire [36:0] _T_5714 = {_T_5705,_T_5594,_T_5591,_T_5588,_T_5585,_T_5582,_T_5579,_T_5576,_T_5573,_T_5570}; // @[Cat.scala 29:58]
  wire [45:0] _T_5723 = {_T_5714,_T_5567,_T_5564,_T_5561,_T_5558,_T_5555,_T_5552,_T_5549,_T_5546,_T_5543}; // @[Cat.scala 29:58]
  wire [54:0] _T_5732 = {_T_5723,_T_5540,_T_5537,_T_5534,_T_5531,_T_5528,_T_5525,_T_5522,_T_5519,_T_5516}; // @[Cat.scala 29:58]
  wire [62:0] _T_5740 = {_T_5732,_T_5513,_T_5510,_T_5507,_T_5504,_T_5501,_T_5498,_T_5495,_T_5492}; // @[Cat.scala 29:58]
  wire  _T_5808 = io_multiplicand[0] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5811 = io_multiplicand[1] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5814 = io_multiplicand[2] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5817 = io_multiplicand[3] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5820 = io_multiplicand[4] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5823 = io_multiplicand[5] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5826 = io_multiplicand[6] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5829 = io_multiplicand[7] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5832 = io_multiplicand[8] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5835 = io_multiplicand[9] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5838 = io_multiplicand[10] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5841 = io_multiplicand[11] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5844 = io_multiplicand[12] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5847 = io_multiplicand[13] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5850 = io_multiplicand[14] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5853 = io_multiplicand[15] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5856 = io_multiplicand[16] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5859 = io_multiplicand[17] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5862 = io_multiplicand[18] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5865 = io_multiplicand[19] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5868 = io_multiplicand[20] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5871 = io_multiplicand[21] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5874 = io_multiplicand[22] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5877 = io_multiplicand[23] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5880 = io_multiplicand[24] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5883 = io_multiplicand[25] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5886 = io_multiplicand[26] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5889 = io_multiplicand[27] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5892 = io_multiplicand[28] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5895 = io_multiplicand[29] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5898 = io_multiplicand[30] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5901 = io_multiplicand[31] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5904 = io_multiplicand[32] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5907 = io_multiplicand[33] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5910 = io_multiplicand[34] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5913 = io_multiplicand[35] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5916 = io_multiplicand[36] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5919 = io_multiplicand[37] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5922 = io_multiplicand[38] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5925 = io_multiplicand[39] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5928 = io_multiplicand[40] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5931 = io_multiplicand[41] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5934 = io_multiplicand[42] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5937 = io_multiplicand[43] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5940 = io_multiplicand[44] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5943 = io_multiplicand[45] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5946 = io_multiplicand[46] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5949 = io_multiplicand[47] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5952 = io_multiplicand[48] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5955 = io_multiplicand[49] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5958 = io_multiplicand[50] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5961 = io_multiplicand[51] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5964 = io_multiplicand[52] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5967 = io_multiplicand[53] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5970 = io_multiplicand[54] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5973 = io_multiplicand[55] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5976 = io_multiplicand[56] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5979 = io_multiplicand[57] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5982 = io_multiplicand[58] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5985 = io_multiplicand[59] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5988 = io_multiplicand[60] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5991 = io_multiplicand[61] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5994 = io_multiplicand[62] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire  _T_5997 = io_multiplicand[63] & io_multiplier[18]; // @[partialprod.scala 16:36]
  wire [9:0] _T_6006 = {_T_5997,_T_5994,_T_5991,_T_5988,_T_5985,_T_5982,_T_5979,_T_5976,_T_5973,_T_5970}; // @[Cat.scala 29:58]
  wire [18:0] _T_6015 = {_T_6006,_T_5967,_T_5964,_T_5961,_T_5958,_T_5955,_T_5952,_T_5949,_T_5946,_T_5943}; // @[Cat.scala 29:58]
  wire [27:0] _T_6024 = {_T_6015,_T_5940,_T_5937,_T_5934,_T_5931,_T_5928,_T_5925,_T_5922,_T_5919,_T_5916}; // @[Cat.scala 29:58]
  wire [36:0] _T_6033 = {_T_6024,_T_5913,_T_5910,_T_5907,_T_5904,_T_5901,_T_5898,_T_5895,_T_5892,_T_5889}; // @[Cat.scala 29:58]
  wire [45:0] _T_6042 = {_T_6033,_T_5886,_T_5883,_T_5880,_T_5877,_T_5874,_T_5871,_T_5868,_T_5865,_T_5862}; // @[Cat.scala 29:58]
  wire [54:0] _T_6051 = {_T_6042,_T_5859,_T_5856,_T_5853,_T_5850,_T_5847,_T_5844,_T_5841,_T_5838,_T_5835}; // @[Cat.scala 29:58]
  wire [62:0] _T_6059 = {_T_6051,_T_5832,_T_5829,_T_5826,_T_5823,_T_5820,_T_5817,_T_5814,_T_5811}; // @[Cat.scala 29:58]
  wire  _T_6127 = io_multiplicand[0] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6130 = io_multiplicand[1] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6133 = io_multiplicand[2] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6136 = io_multiplicand[3] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6139 = io_multiplicand[4] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6142 = io_multiplicand[5] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6145 = io_multiplicand[6] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6148 = io_multiplicand[7] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6151 = io_multiplicand[8] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6154 = io_multiplicand[9] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6157 = io_multiplicand[10] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6160 = io_multiplicand[11] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6163 = io_multiplicand[12] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6166 = io_multiplicand[13] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6169 = io_multiplicand[14] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6172 = io_multiplicand[15] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6175 = io_multiplicand[16] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6178 = io_multiplicand[17] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6181 = io_multiplicand[18] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6184 = io_multiplicand[19] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6187 = io_multiplicand[20] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6190 = io_multiplicand[21] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6193 = io_multiplicand[22] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6196 = io_multiplicand[23] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6199 = io_multiplicand[24] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6202 = io_multiplicand[25] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6205 = io_multiplicand[26] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6208 = io_multiplicand[27] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6211 = io_multiplicand[28] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6214 = io_multiplicand[29] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6217 = io_multiplicand[30] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6220 = io_multiplicand[31] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6223 = io_multiplicand[32] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6226 = io_multiplicand[33] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6229 = io_multiplicand[34] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6232 = io_multiplicand[35] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6235 = io_multiplicand[36] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6238 = io_multiplicand[37] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6241 = io_multiplicand[38] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6244 = io_multiplicand[39] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6247 = io_multiplicand[40] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6250 = io_multiplicand[41] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6253 = io_multiplicand[42] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6256 = io_multiplicand[43] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6259 = io_multiplicand[44] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6262 = io_multiplicand[45] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6265 = io_multiplicand[46] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6268 = io_multiplicand[47] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6271 = io_multiplicand[48] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6274 = io_multiplicand[49] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6277 = io_multiplicand[50] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6280 = io_multiplicand[51] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6283 = io_multiplicand[52] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6286 = io_multiplicand[53] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6289 = io_multiplicand[54] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6292 = io_multiplicand[55] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6295 = io_multiplicand[56] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6298 = io_multiplicand[57] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6301 = io_multiplicand[58] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6304 = io_multiplicand[59] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6307 = io_multiplicand[60] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6310 = io_multiplicand[61] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6313 = io_multiplicand[62] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire  _T_6316 = io_multiplicand[63] & io_multiplier[19]; // @[partialprod.scala 16:36]
  wire [9:0] _T_6325 = {_T_6316,_T_6313,_T_6310,_T_6307,_T_6304,_T_6301,_T_6298,_T_6295,_T_6292,_T_6289}; // @[Cat.scala 29:58]
  wire [18:0] _T_6334 = {_T_6325,_T_6286,_T_6283,_T_6280,_T_6277,_T_6274,_T_6271,_T_6268,_T_6265,_T_6262}; // @[Cat.scala 29:58]
  wire [27:0] _T_6343 = {_T_6334,_T_6259,_T_6256,_T_6253,_T_6250,_T_6247,_T_6244,_T_6241,_T_6238,_T_6235}; // @[Cat.scala 29:58]
  wire [36:0] _T_6352 = {_T_6343,_T_6232,_T_6229,_T_6226,_T_6223,_T_6220,_T_6217,_T_6214,_T_6211,_T_6208}; // @[Cat.scala 29:58]
  wire [45:0] _T_6361 = {_T_6352,_T_6205,_T_6202,_T_6199,_T_6196,_T_6193,_T_6190,_T_6187,_T_6184,_T_6181}; // @[Cat.scala 29:58]
  wire [54:0] _T_6370 = {_T_6361,_T_6178,_T_6175,_T_6172,_T_6169,_T_6166,_T_6163,_T_6160,_T_6157,_T_6154}; // @[Cat.scala 29:58]
  wire [62:0] _T_6378 = {_T_6370,_T_6151,_T_6148,_T_6145,_T_6142,_T_6139,_T_6136,_T_6133,_T_6130}; // @[Cat.scala 29:58]
  wire  _T_6446 = io_multiplicand[0] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6449 = io_multiplicand[1] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6452 = io_multiplicand[2] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6455 = io_multiplicand[3] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6458 = io_multiplicand[4] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6461 = io_multiplicand[5] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6464 = io_multiplicand[6] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6467 = io_multiplicand[7] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6470 = io_multiplicand[8] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6473 = io_multiplicand[9] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6476 = io_multiplicand[10] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6479 = io_multiplicand[11] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6482 = io_multiplicand[12] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6485 = io_multiplicand[13] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6488 = io_multiplicand[14] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6491 = io_multiplicand[15] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6494 = io_multiplicand[16] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6497 = io_multiplicand[17] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6500 = io_multiplicand[18] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6503 = io_multiplicand[19] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6506 = io_multiplicand[20] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6509 = io_multiplicand[21] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6512 = io_multiplicand[22] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6515 = io_multiplicand[23] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6518 = io_multiplicand[24] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6521 = io_multiplicand[25] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6524 = io_multiplicand[26] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6527 = io_multiplicand[27] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6530 = io_multiplicand[28] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6533 = io_multiplicand[29] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6536 = io_multiplicand[30] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6539 = io_multiplicand[31] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6542 = io_multiplicand[32] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6545 = io_multiplicand[33] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6548 = io_multiplicand[34] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6551 = io_multiplicand[35] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6554 = io_multiplicand[36] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6557 = io_multiplicand[37] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6560 = io_multiplicand[38] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6563 = io_multiplicand[39] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6566 = io_multiplicand[40] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6569 = io_multiplicand[41] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6572 = io_multiplicand[42] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6575 = io_multiplicand[43] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6578 = io_multiplicand[44] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6581 = io_multiplicand[45] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6584 = io_multiplicand[46] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6587 = io_multiplicand[47] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6590 = io_multiplicand[48] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6593 = io_multiplicand[49] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6596 = io_multiplicand[50] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6599 = io_multiplicand[51] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6602 = io_multiplicand[52] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6605 = io_multiplicand[53] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6608 = io_multiplicand[54] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6611 = io_multiplicand[55] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6614 = io_multiplicand[56] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6617 = io_multiplicand[57] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6620 = io_multiplicand[58] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6623 = io_multiplicand[59] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6626 = io_multiplicand[60] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6629 = io_multiplicand[61] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6632 = io_multiplicand[62] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire  _T_6635 = io_multiplicand[63] & io_multiplier[20]; // @[partialprod.scala 16:36]
  wire [9:0] _T_6644 = {_T_6635,_T_6632,_T_6629,_T_6626,_T_6623,_T_6620,_T_6617,_T_6614,_T_6611,_T_6608}; // @[Cat.scala 29:58]
  wire [18:0] _T_6653 = {_T_6644,_T_6605,_T_6602,_T_6599,_T_6596,_T_6593,_T_6590,_T_6587,_T_6584,_T_6581}; // @[Cat.scala 29:58]
  wire [27:0] _T_6662 = {_T_6653,_T_6578,_T_6575,_T_6572,_T_6569,_T_6566,_T_6563,_T_6560,_T_6557,_T_6554}; // @[Cat.scala 29:58]
  wire [36:0] _T_6671 = {_T_6662,_T_6551,_T_6548,_T_6545,_T_6542,_T_6539,_T_6536,_T_6533,_T_6530,_T_6527}; // @[Cat.scala 29:58]
  wire [45:0] _T_6680 = {_T_6671,_T_6524,_T_6521,_T_6518,_T_6515,_T_6512,_T_6509,_T_6506,_T_6503,_T_6500}; // @[Cat.scala 29:58]
  wire [54:0] _T_6689 = {_T_6680,_T_6497,_T_6494,_T_6491,_T_6488,_T_6485,_T_6482,_T_6479,_T_6476,_T_6473}; // @[Cat.scala 29:58]
  wire [62:0] _T_6697 = {_T_6689,_T_6470,_T_6467,_T_6464,_T_6461,_T_6458,_T_6455,_T_6452,_T_6449}; // @[Cat.scala 29:58]
  wire  _T_6765 = io_multiplicand[0] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6768 = io_multiplicand[1] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6771 = io_multiplicand[2] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6774 = io_multiplicand[3] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6777 = io_multiplicand[4] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6780 = io_multiplicand[5] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6783 = io_multiplicand[6] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6786 = io_multiplicand[7] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6789 = io_multiplicand[8] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6792 = io_multiplicand[9] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6795 = io_multiplicand[10] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6798 = io_multiplicand[11] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6801 = io_multiplicand[12] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6804 = io_multiplicand[13] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6807 = io_multiplicand[14] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6810 = io_multiplicand[15] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6813 = io_multiplicand[16] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6816 = io_multiplicand[17] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6819 = io_multiplicand[18] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6822 = io_multiplicand[19] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6825 = io_multiplicand[20] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6828 = io_multiplicand[21] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6831 = io_multiplicand[22] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6834 = io_multiplicand[23] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6837 = io_multiplicand[24] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6840 = io_multiplicand[25] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6843 = io_multiplicand[26] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6846 = io_multiplicand[27] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6849 = io_multiplicand[28] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6852 = io_multiplicand[29] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6855 = io_multiplicand[30] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6858 = io_multiplicand[31] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6861 = io_multiplicand[32] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6864 = io_multiplicand[33] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6867 = io_multiplicand[34] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6870 = io_multiplicand[35] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6873 = io_multiplicand[36] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6876 = io_multiplicand[37] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6879 = io_multiplicand[38] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6882 = io_multiplicand[39] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6885 = io_multiplicand[40] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6888 = io_multiplicand[41] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6891 = io_multiplicand[42] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6894 = io_multiplicand[43] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6897 = io_multiplicand[44] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6900 = io_multiplicand[45] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6903 = io_multiplicand[46] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6906 = io_multiplicand[47] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6909 = io_multiplicand[48] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6912 = io_multiplicand[49] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6915 = io_multiplicand[50] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6918 = io_multiplicand[51] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6921 = io_multiplicand[52] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6924 = io_multiplicand[53] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6927 = io_multiplicand[54] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6930 = io_multiplicand[55] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6933 = io_multiplicand[56] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6936 = io_multiplicand[57] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6939 = io_multiplicand[58] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6942 = io_multiplicand[59] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6945 = io_multiplicand[60] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6948 = io_multiplicand[61] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6951 = io_multiplicand[62] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire  _T_6954 = io_multiplicand[63] & io_multiplier[21]; // @[partialprod.scala 16:36]
  wire [9:0] _T_6963 = {_T_6954,_T_6951,_T_6948,_T_6945,_T_6942,_T_6939,_T_6936,_T_6933,_T_6930,_T_6927}; // @[Cat.scala 29:58]
  wire [18:0] _T_6972 = {_T_6963,_T_6924,_T_6921,_T_6918,_T_6915,_T_6912,_T_6909,_T_6906,_T_6903,_T_6900}; // @[Cat.scala 29:58]
  wire [27:0] _T_6981 = {_T_6972,_T_6897,_T_6894,_T_6891,_T_6888,_T_6885,_T_6882,_T_6879,_T_6876,_T_6873}; // @[Cat.scala 29:58]
  wire [36:0] _T_6990 = {_T_6981,_T_6870,_T_6867,_T_6864,_T_6861,_T_6858,_T_6855,_T_6852,_T_6849,_T_6846}; // @[Cat.scala 29:58]
  wire [45:0] _T_6999 = {_T_6990,_T_6843,_T_6840,_T_6837,_T_6834,_T_6831,_T_6828,_T_6825,_T_6822,_T_6819}; // @[Cat.scala 29:58]
  wire [54:0] _T_7008 = {_T_6999,_T_6816,_T_6813,_T_6810,_T_6807,_T_6804,_T_6801,_T_6798,_T_6795,_T_6792}; // @[Cat.scala 29:58]
  wire [62:0] _T_7016 = {_T_7008,_T_6789,_T_6786,_T_6783,_T_6780,_T_6777,_T_6774,_T_6771,_T_6768}; // @[Cat.scala 29:58]
  wire  _T_7084 = io_multiplicand[0] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7087 = io_multiplicand[1] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7090 = io_multiplicand[2] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7093 = io_multiplicand[3] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7096 = io_multiplicand[4] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7099 = io_multiplicand[5] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7102 = io_multiplicand[6] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7105 = io_multiplicand[7] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7108 = io_multiplicand[8] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7111 = io_multiplicand[9] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7114 = io_multiplicand[10] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7117 = io_multiplicand[11] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7120 = io_multiplicand[12] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7123 = io_multiplicand[13] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7126 = io_multiplicand[14] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7129 = io_multiplicand[15] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7132 = io_multiplicand[16] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7135 = io_multiplicand[17] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7138 = io_multiplicand[18] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7141 = io_multiplicand[19] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7144 = io_multiplicand[20] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7147 = io_multiplicand[21] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7150 = io_multiplicand[22] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7153 = io_multiplicand[23] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7156 = io_multiplicand[24] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7159 = io_multiplicand[25] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7162 = io_multiplicand[26] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7165 = io_multiplicand[27] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7168 = io_multiplicand[28] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7171 = io_multiplicand[29] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7174 = io_multiplicand[30] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7177 = io_multiplicand[31] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7180 = io_multiplicand[32] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7183 = io_multiplicand[33] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7186 = io_multiplicand[34] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7189 = io_multiplicand[35] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7192 = io_multiplicand[36] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7195 = io_multiplicand[37] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7198 = io_multiplicand[38] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7201 = io_multiplicand[39] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7204 = io_multiplicand[40] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7207 = io_multiplicand[41] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7210 = io_multiplicand[42] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7213 = io_multiplicand[43] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7216 = io_multiplicand[44] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7219 = io_multiplicand[45] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7222 = io_multiplicand[46] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7225 = io_multiplicand[47] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7228 = io_multiplicand[48] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7231 = io_multiplicand[49] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7234 = io_multiplicand[50] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7237 = io_multiplicand[51] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7240 = io_multiplicand[52] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7243 = io_multiplicand[53] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7246 = io_multiplicand[54] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7249 = io_multiplicand[55] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7252 = io_multiplicand[56] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7255 = io_multiplicand[57] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7258 = io_multiplicand[58] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7261 = io_multiplicand[59] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7264 = io_multiplicand[60] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7267 = io_multiplicand[61] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7270 = io_multiplicand[62] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire  _T_7273 = io_multiplicand[63] & io_multiplier[22]; // @[partialprod.scala 16:36]
  wire [9:0] _T_7282 = {_T_7273,_T_7270,_T_7267,_T_7264,_T_7261,_T_7258,_T_7255,_T_7252,_T_7249,_T_7246}; // @[Cat.scala 29:58]
  wire [18:0] _T_7291 = {_T_7282,_T_7243,_T_7240,_T_7237,_T_7234,_T_7231,_T_7228,_T_7225,_T_7222,_T_7219}; // @[Cat.scala 29:58]
  wire [27:0] _T_7300 = {_T_7291,_T_7216,_T_7213,_T_7210,_T_7207,_T_7204,_T_7201,_T_7198,_T_7195,_T_7192}; // @[Cat.scala 29:58]
  wire [36:0] _T_7309 = {_T_7300,_T_7189,_T_7186,_T_7183,_T_7180,_T_7177,_T_7174,_T_7171,_T_7168,_T_7165}; // @[Cat.scala 29:58]
  wire [45:0] _T_7318 = {_T_7309,_T_7162,_T_7159,_T_7156,_T_7153,_T_7150,_T_7147,_T_7144,_T_7141,_T_7138}; // @[Cat.scala 29:58]
  wire [54:0] _T_7327 = {_T_7318,_T_7135,_T_7132,_T_7129,_T_7126,_T_7123,_T_7120,_T_7117,_T_7114,_T_7111}; // @[Cat.scala 29:58]
  wire [62:0] _T_7335 = {_T_7327,_T_7108,_T_7105,_T_7102,_T_7099,_T_7096,_T_7093,_T_7090,_T_7087}; // @[Cat.scala 29:58]
  wire  _T_7403 = io_multiplicand[0] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7406 = io_multiplicand[1] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7409 = io_multiplicand[2] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7412 = io_multiplicand[3] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7415 = io_multiplicand[4] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7418 = io_multiplicand[5] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7421 = io_multiplicand[6] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7424 = io_multiplicand[7] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7427 = io_multiplicand[8] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7430 = io_multiplicand[9] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7433 = io_multiplicand[10] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7436 = io_multiplicand[11] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7439 = io_multiplicand[12] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7442 = io_multiplicand[13] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7445 = io_multiplicand[14] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7448 = io_multiplicand[15] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7451 = io_multiplicand[16] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7454 = io_multiplicand[17] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7457 = io_multiplicand[18] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7460 = io_multiplicand[19] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7463 = io_multiplicand[20] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7466 = io_multiplicand[21] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7469 = io_multiplicand[22] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7472 = io_multiplicand[23] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7475 = io_multiplicand[24] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7478 = io_multiplicand[25] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7481 = io_multiplicand[26] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7484 = io_multiplicand[27] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7487 = io_multiplicand[28] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7490 = io_multiplicand[29] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7493 = io_multiplicand[30] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7496 = io_multiplicand[31] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7499 = io_multiplicand[32] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7502 = io_multiplicand[33] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7505 = io_multiplicand[34] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7508 = io_multiplicand[35] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7511 = io_multiplicand[36] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7514 = io_multiplicand[37] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7517 = io_multiplicand[38] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7520 = io_multiplicand[39] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7523 = io_multiplicand[40] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7526 = io_multiplicand[41] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7529 = io_multiplicand[42] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7532 = io_multiplicand[43] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7535 = io_multiplicand[44] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7538 = io_multiplicand[45] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7541 = io_multiplicand[46] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7544 = io_multiplicand[47] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7547 = io_multiplicand[48] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7550 = io_multiplicand[49] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7553 = io_multiplicand[50] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7556 = io_multiplicand[51] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7559 = io_multiplicand[52] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7562 = io_multiplicand[53] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7565 = io_multiplicand[54] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7568 = io_multiplicand[55] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7571 = io_multiplicand[56] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7574 = io_multiplicand[57] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7577 = io_multiplicand[58] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7580 = io_multiplicand[59] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7583 = io_multiplicand[60] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7586 = io_multiplicand[61] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7589 = io_multiplicand[62] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire  _T_7592 = io_multiplicand[63] & io_multiplier[23]; // @[partialprod.scala 16:36]
  wire [9:0] _T_7601 = {_T_7592,_T_7589,_T_7586,_T_7583,_T_7580,_T_7577,_T_7574,_T_7571,_T_7568,_T_7565}; // @[Cat.scala 29:58]
  wire [18:0] _T_7610 = {_T_7601,_T_7562,_T_7559,_T_7556,_T_7553,_T_7550,_T_7547,_T_7544,_T_7541,_T_7538}; // @[Cat.scala 29:58]
  wire [27:0] _T_7619 = {_T_7610,_T_7535,_T_7532,_T_7529,_T_7526,_T_7523,_T_7520,_T_7517,_T_7514,_T_7511}; // @[Cat.scala 29:58]
  wire [36:0] _T_7628 = {_T_7619,_T_7508,_T_7505,_T_7502,_T_7499,_T_7496,_T_7493,_T_7490,_T_7487,_T_7484}; // @[Cat.scala 29:58]
  wire [45:0] _T_7637 = {_T_7628,_T_7481,_T_7478,_T_7475,_T_7472,_T_7469,_T_7466,_T_7463,_T_7460,_T_7457}; // @[Cat.scala 29:58]
  wire [54:0] _T_7646 = {_T_7637,_T_7454,_T_7451,_T_7448,_T_7445,_T_7442,_T_7439,_T_7436,_T_7433,_T_7430}; // @[Cat.scala 29:58]
  wire [62:0] _T_7654 = {_T_7646,_T_7427,_T_7424,_T_7421,_T_7418,_T_7415,_T_7412,_T_7409,_T_7406}; // @[Cat.scala 29:58]
  wire  _T_7722 = io_multiplicand[0] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7725 = io_multiplicand[1] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7728 = io_multiplicand[2] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7731 = io_multiplicand[3] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7734 = io_multiplicand[4] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7737 = io_multiplicand[5] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7740 = io_multiplicand[6] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7743 = io_multiplicand[7] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7746 = io_multiplicand[8] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7749 = io_multiplicand[9] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7752 = io_multiplicand[10] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7755 = io_multiplicand[11] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7758 = io_multiplicand[12] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7761 = io_multiplicand[13] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7764 = io_multiplicand[14] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7767 = io_multiplicand[15] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7770 = io_multiplicand[16] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7773 = io_multiplicand[17] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7776 = io_multiplicand[18] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7779 = io_multiplicand[19] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7782 = io_multiplicand[20] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7785 = io_multiplicand[21] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7788 = io_multiplicand[22] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7791 = io_multiplicand[23] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7794 = io_multiplicand[24] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7797 = io_multiplicand[25] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7800 = io_multiplicand[26] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7803 = io_multiplicand[27] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7806 = io_multiplicand[28] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7809 = io_multiplicand[29] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7812 = io_multiplicand[30] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7815 = io_multiplicand[31] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7818 = io_multiplicand[32] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7821 = io_multiplicand[33] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7824 = io_multiplicand[34] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7827 = io_multiplicand[35] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7830 = io_multiplicand[36] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7833 = io_multiplicand[37] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7836 = io_multiplicand[38] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7839 = io_multiplicand[39] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7842 = io_multiplicand[40] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7845 = io_multiplicand[41] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7848 = io_multiplicand[42] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7851 = io_multiplicand[43] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7854 = io_multiplicand[44] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7857 = io_multiplicand[45] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7860 = io_multiplicand[46] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7863 = io_multiplicand[47] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7866 = io_multiplicand[48] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7869 = io_multiplicand[49] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7872 = io_multiplicand[50] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7875 = io_multiplicand[51] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7878 = io_multiplicand[52] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7881 = io_multiplicand[53] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7884 = io_multiplicand[54] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7887 = io_multiplicand[55] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7890 = io_multiplicand[56] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7893 = io_multiplicand[57] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7896 = io_multiplicand[58] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7899 = io_multiplicand[59] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7902 = io_multiplicand[60] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7905 = io_multiplicand[61] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7908 = io_multiplicand[62] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire  _T_7911 = io_multiplicand[63] & io_multiplier[24]; // @[partialprod.scala 16:36]
  wire [9:0] _T_7920 = {_T_7911,_T_7908,_T_7905,_T_7902,_T_7899,_T_7896,_T_7893,_T_7890,_T_7887,_T_7884}; // @[Cat.scala 29:58]
  wire [18:0] _T_7929 = {_T_7920,_T_7881,_T_7878,_T_7875,_T_7872,_T_7869,_T_7866,_T_7863,_T_7860,_T_7857}; // @[Cat.scala 29:58]
  wire [27:0] _T_7938 = {_T_7929,_T_7854,_T_7851,_T_7848,_T_7845,_T_7842,_T_7839,_T_7836,_T_7833,_T_7830}; // @[Cat.scala 29:58]
  wire [36:0] _T_7947 = {_T_7938,_T_7827,_T_7824,_T_7821,_T_7818,_T_7815,_T_7812,_T_7809,_T_7806,_T_7803}; // @[Cat.scala 29:58]
  wire [45:0] _T_7956 = {_T_7947,_T_7800,_T_7797,_T_7794,_T_7791,_T_7788,_T_7785,_T_7782,_T_7779,_T_7776}; // @[Cat.scala 29:58]
  wire [54:0] _T_7965 = {_T_7956,_T_7773,_T_7770,_T_7767,_T_7764,_T_7761,_T_7758,_T_7755,_T_7752,_T_7749}; // @[Cat.scala 29:58]
  wire [62:0] _T_7973 = {_T_7965,_T_7746,_T_7743,_T_7740,_T_7737,_T_7734,_T_7731,_T_7728,_T_7725}; // @[Cat.scala 29:58]
  wire  _T_8041 = io_multiplicand[0] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8044 = io_multiplicand[1] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8047 = io_multiplicand[2] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8050 = io_multiplicand[3] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8053 = io_multiplicand[4] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8056 = io_multiplicand[5] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8059 = io_multiplicand[6] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8062 = io_multiplicand[7] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8065 = io_multiplicand[8] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8068 = io_multiplicand[9] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8071 = io_multiplicand[10] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8074 = io_multiplicand[11] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8077 = io_multiplicand[12] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8080 = io_multiplicand[13] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8083 = io_multiplicand[14] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8086 = io_multiplicand[15] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8089 = io_multiplicand[16] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8092 = io_multiplicand[17] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8095 = io_multiplicand[18] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8098 = io_multiplicand[19] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8101 = io_multiplicand[20] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8104 = io_multiplicand[21] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8107 = io_multiplicand[22] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8110 = io_multiplicand[23] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8113 = io_multiplicand[24] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8116 = io_multiplicand[25] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8119 = io_multiplicand[26] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8122 = io_multiplicand[27] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8125 = io_multiplicand[28] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8128 = io_multiplicand[29] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8131 = io_multiplicand[30] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8134 = io_multiplicand[31] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8137 = io_multiplicand[32] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8140 = io_multiplicand[33] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8143 = io_multiplicand[34] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8146 = io_multiplicand[35] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8149 = io_multiplicand[36] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8152 = io_multiplicand[37] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8155 = io_multiplicand[38] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8158 = io_multiplicand[39] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8161 = io_multiplicand[40] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8164 = io_multiplicand[41] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8167 = io_multiplicand[42] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8170 = io_multiplicand[43] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8173 = io_multiplicand[44] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8176 = io_multiplicand[45] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8179 = io_multiplicand[46] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8182 = io_multiplicand[47] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8185 = io_multiplicand[48] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8188 = io_multiplicand[49] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8191 = io_multiplicand[50] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8194 = io_multiplicand[51] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8197 = io_multiplicand[52] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8200 = io_multiplicand[53] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8203 = io_multiplicand[54] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8206 = io_multiplicand[55] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8209 = io_multiplicand[56] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8212 = io_multiplicand[57] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8215 = io_multiplicand[58] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8218 = io_multiplicand[59] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8221 = io_multiplicand[60] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8224 = io_multiplicand[61] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8227 = io_multiplicand[62] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire  _T_8230 = io_multiplicand[63] & io_multiplier[25]; // @[partialprod.scala 16:36]
  wire [9:0] _T_8239 = {_T_8230,_T_8227,_T_8224,_T_8221,_T_8218,_T_8215,_T_8212,_T_8209,_T_8206,_T_8203}; // @[Cat.scala 29:58]
  wire [18:0] _T_8248 = {_T_8239,_T_8200,_T_8197,_T_8194,_T_8191,_T_8188,_T_8185,_T_8182,_T_8179,_T_8176}; // @[Cat.scala 29:58]
  wire [27:0] _T_8257 = {_T_8248,_T_8173,_T_8170,_T_8167,_T_8164,_T_8161,_T_8158,_T_8155,_T_8152,_T_8149}; // @[Cat.scala 29:58]
  wire [36:0] _T_8266 = {_T_8257,_T_8146,_T_8143,_T_8140,_T_8137,_T_8134,_T_8131,_T_8128,_T_8125,_T_8122}; // @[Cat.scala 29:58]
  wire [45:0] _T_8275 = {_T_8266,_T_8119,_T_8116,_T_8113,_T_8110,_T_8107,_T_8104,_T_8101,_T_8098,_T_8095}; // @[Cat.scala 29:58]
  wire [54:0] _T_8284 = {_T_8275,_T_8092,_T_8089,_T_8086,_T_8083,_T_8080,_T_8077,_T_8074,_T_8071,_T_8068}; // @[Cat.scala 29:58]
  wire [62:0] _T_8292 = {_T_8284,_T_8065,_T_8062,_T_8059,_T_8056,_T_8053,_T_8050,_T_8047,_T_8044}; // @[Cat.scala 29:58]
  wire  _T_8360 = io_multiplicand[0] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8363 = io_multiplicand[1] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8366 = io_multiplicand[2] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8369 = io_multiplicand[3] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8372 = io_multiplicand[4] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8375 = io_multiplicand[5] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8378 = io_multiplicand[6] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8381 = io_multiplicand[7] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8384 = io_multiplicand[8] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8387 = io_multiplicand[9] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8390 = io_multiplicand[10] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8393 = io_multiplicand[11] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8396 = io_multiplicand[12] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8399 = io_multiplicand[13] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8402 = io_multiplicand[14] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8405 = io_multiplicand[15] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8408 = io_multiplicand[16] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8411 = io_multiplicand[17] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8414 = io_multiplicand[18] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8417 = io_multiplicand[19] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8420 = io_multiplicand[20] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8423 = io_multiplicand[21] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8426 = io_multiplicand[22] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8429 = io_multiplicand[23] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8432 = io_multiplicand[24] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8435 = io_multiplicand[25] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8438 = io_multiplicand[26] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8441 = io_multiplicand[27] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8444 = io_multiplicand[28] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8447 = io_multiplicand[29] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8450 = io_multiplicand[30] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8453 = io_multiplicand[31] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8456 = io_multiplicand[32] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8459 = io_multiplicand[33] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8462 = io_multiplicand[34] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8465 = io_multiplicand[35] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8468 = io_multiplicand[36] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8471 = io_multiplicand[37] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8474 = io_multiplicand[38] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8477 = io_multiplicand[39] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8480 = io_multiplicand[40] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8483 = io_multiplicand[41] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8486 = io_multiplicand[42] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8489 = io_multiplicand[43] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8492 = io_multiplicand[44] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8495 = io_multiplicand[45] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8498 = io_multiplicand[46] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8501 = io_multiplicand[47] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8504 = io_multiplicand[48] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8507 = io_multiplicand[49] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8510 = io_multiplicand[50] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8513 = io_multiplicand[51] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8516 = io_multiplicand[52] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8519 = io_multiplicand[53] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8522 = io_multiplicand[54] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8525 = io_multiplicand[55] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8528 = io_multiplicand[56] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8531 = io_multiplicand[57] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8534 = io_multiplicand[58] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8537 = io_multiplicand[59] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8540 = io_multiplicand[60] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8543 = io_multiplicand[61] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8546 = io_multiplicand[62] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire  _T_8549 = io_multiplicand[63] & io_multiplier[26]; // @[partialprod.scala 16:36]
  wire [9:0] _T_8558 = {_T_8549,_T_8546,_T_8543,_T_8540,_T_8537,_T_8534,_T_8531,_T_8528,_T_8525,_T_8522}; // @[Cat.scala 29:58]
  wire [18:0] _T_8567 = {_T_8558,_T_8519,_T_8516,_T_8513,_T_8510,_T_8507,_T_8504,_T_8501,_T_8498,_T_8495}; // @[Cat.scala 29:58]
  wire [27:0] _T_8576 = {_T_8567,_T_8492,_T_8489,_T_8486,_T_8483,_T_8480,_T_8477,_T_8474,_T_8471,_T_8468}; // @[Cat.scala 29:58]
  wire [36:0] _T_8585 = {_T_8576,_T_8465,_T_8462,_T_8459,_T_8456,_T_8453,_T_8450,_T_8447,_T_8444,_T_8441}; // @[Cat.scala 29:58]
  wire [45:0] _T_8594 = {_T_8585,_T_8438,_T_8435,_T_8432,_T_8429,_T_8426,_T_8423,_T_8420,_T_8417,_T_8414}; // @[Cat.scala 29:58]
  wire [54:0] _T_8603 = {_T_8594,_T_8411,_T_8408,_T_8405,_T_8402,_T_8399,_T_8396,_T_8393,_T_8390,_T_8387}; // @[Cat.scala 29:58]
  wire [62:0] _T_8611 = {_T_8603,_T_8384,_T_8381,_T_8378,_T_8375,_T_8372,_T_8369,_T_8366,_T_8363}; // @[Cat.scala 29:58]
  wire  _T_8679 = io_multiplicand[0] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8682 = io_multiplicand[1] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8685 = io_multiplicand[2] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8688 = io_multiplicand[3] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8691 = io_multiplicand[4] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8694 = io_multiplicand[5] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8697 = io_multiplicand[6] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8700 = io_multiplicand[7] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8703 = io_multiplicand[8] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8706 = io_multiplicand[9] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8709 = io_multiplicand[10] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8712 = io_multiplicand[11] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8715 = io_multiplicand[12] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8718 = io_multiplicand[13] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8721 = io_multiplicand[14] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8724 = io_multiplicand[15] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8727 = io_multiplicand[16] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8730 = io_multiplicand[17] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8733 = io_multiplicand[18] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8736 = io_multiplicand[19] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8739 = io_multiplicand[20] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8742 = io_multiplicand[21] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8745 = io_multiplicand[22] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8748 = io_multiplicand[23] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8751 = io_multiplicand[24] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8754 = io_multiplicand[25] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8757 = io_multiplicand[26] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8760 = io_multiplicand[27] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8763 = io_multiplicand[28] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8766 = io_multiplicand[29] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8769 = io_multiplicand[30] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8772 = io_multiplicand[31] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8775 = io_multiplicand[32] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8778 = io_multiplicand[33] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8781 = io_multiplicand[34] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8784 = io_multiplicand[35] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8787 = io_multiplicand[36] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8790 = io_multiplicand[37] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8793 = io_multiplicand[38] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8796 = io_multiplicand[39] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8799 = io_multiplicand[40] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8802 = io_multiplicand[41] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8805 = io_multiplicand[42] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8808 = io_multiplicand[43] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8811 = io_multiplicand[44] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8814 = io_multiplicand[45] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8817 = io_multiplicand[46] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8820 = io_multiplicand[47] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8823 = io_multiplicand[48] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8826 = io_multiplicand[49] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8829 = io_multiplicand[50] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8832 = io_multiplicand[51] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8835 = io_multiplicand[52] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8838 = io_multiplicand[53] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8841 = io_multiplicand[54] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8844 = io_multiplicand[55] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8847 = io_multiplicand[56] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8850 = io_multiplicand[57] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8853 = io_multiplicand[58] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8856 = io_multiplicand[59] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8859 = io_multiplicand[60] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8862 = io_multiplicand[61] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8865 = io_multiplicand[62] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire  _T_8868 = io_multiplicand[63] & io_multiplier[27]; // @[partialprod.scala 16:36]
  wire [9:0] _T_8877 = {_T_8868,_T_8865,_T_8862,_T_8859,_T_8856,_T_8853,_T_8850,_T_8847,_T_8844,_T_8841}; // @[Cat.scala 29:58]
  wire [18:0] _T_8886 = {_T_8877,_T_8838,_T_8835,_T_8832,_T_8829,_T_8826,_T_8823,_T_8820,_T_8817,_T_8814}; // @[Cat.scala 29:58]
  wire [27:0] _T_8895 = {_T_8886,_T_8811,_T_8808,_T_8805,_T_8802,_T_8799,_T_8796,_T_8793,_T_8790,_T_8787}; // @[Cat.scala 29:58]
  wire [36:0] _T_8904 = {_T_8895,_T_8784,_T_8781,_T_8778,_T_8775,_T_8772,_T_8769,_T_8766,_T_8763,_T_8760}; // @[Cat.scala 29:58]
  wire [45:0] _T_8913 = {_T_8904,_T_8757,_T_8754,_T_8751,_T_8748,_T_8745,_T_8742,_T_8739,_T_8736,_T_8733}; // @[Cat.scala 29:58]
  wire [54:0] _T_8922 = {_T_8913,_T_8730,_T_8727,_T_8724,_T_8721,_T_8718,_T_8715,_T_8712,_T_8709,_T_8706}; // @[Cat.scala 29:58]
  wire [62:0] _T_8930 = {_T_8922,_T_8703,_T_8700,_T_8697,_T_8694,_T_8691,_T_8688,_T_8685,_T_8682}; // @[Cat.scala 29:58]
  wire  _T_8998 = io_multiplicand[0] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9001 = io_multiplicand[1] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9004 = io_multiplicand[2] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9007 = io_multiplicand[3] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9010 = io_multiplicand[4] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9013 = io_multiplicand[5] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9016 = io_multiplicand[6] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9019 = io_multiplicand[7] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9022 = io_multiplicand[8] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9025 = io_multiplicand[9] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9028 = io_multiplicand[10] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9031 = io_multiplicand[11] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9034 = io_multiplicand[12] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9037 = io_multiplicand[13] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9040 = io_multiplicand[14] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9043 = io_multiplicand[15] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9046 = io_multiplicand[16] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9049 = io_multiplicand[17] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9052 = io_multiplicand[18] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9055 = io_multiplicand[19] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9058 = io_multiplicand[20] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9061 = io_multiplicand[21] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9064 = io_multiplicand[22] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9067 = io_multiplicand[23] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9070 = io_multiplicand[24] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9073 = io_multiplicand[25] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9076 = io_multiplicand[26] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9079 = io_multiplicand[27] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9082 = io_multiplicand[28] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9085 = io_multiplicand[29] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9088 = io_multiplicand[30] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9091 = io_multiplicand[31] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9094 = io_multiplicand[32] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9097 = io_multiplicand[33] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9100 = io_multiplicand[34] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9103 = io_multiplicand[35] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9106 = io_multiplicand[36] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9109 = io_multiplicand[37] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9112 = io_multiplicand[38] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9115 = io_multiplicand[39] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9118 = io_multiplicand[40] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9121 = io_multiplicand[41] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9124 = io_multiplicand[42] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9127 = io_multiplicand[43] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9130 = io_multiplicand[44] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9133 = io_multiplicand[45] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9136 = io_multiplicand[46] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9139 = io_multiplicand[47] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9142 = io_multiplicand[48] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9145 = io_multiplicand[49] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9148 = io_multiplicand[50] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9151 = io_multiplicand[51] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9154 = io_multiplicand[52] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9157 = io_multiplicand[53] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9160 = io_multiplicand[54] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9163 = io_multiplicand[55] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9166 = io_multiplicand[56] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9169 = io_multiplicand[57] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9172 = io_multiplicand[58] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9175 = io_multiplicand[59] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9178 = io_multiplicand[60] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9181 = io_multiplicand[61] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9184 = io_multiplicand[62] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire  _T_9187 = io_multiplicand[63] & io_multiplier[28]; // @[partialprod.scala 16:36]
  wire [9:0] _T_9196 = {_T_9187,_T_9184,_T_9181,_T_9178,_T_9175,_T_9172,_T_9169,_T_9166,_T_9163,_T_9160}; // @[Cat.scala 29:58]
  wire [18:0] _T_9205 = {_T_9196,_T_9157,_T_9154,_T_9151,_T_9148,_T_9145,_T_9142,_T_9139,_T_9136,_T_9133}; // @[Cat.scala 29:58]
  wire [27:0] _T_9214 = {_T_9205,_T_9130,_T_9127,_T_9124,_T_9121,_T_9118,_T_9115,_T_9112,_T_9109,_T_9106}; // @[Cat.scala 29:58]
  wire [36:0] _T_9223 = {_T_9214,_T_9103,_T_9100,_T_9097,_T_9094,_T_9091,_T_9088,_T_9085,_T_9082,_T_9079}; // @[Cat.scala 29:58]
  wire [45:0] _T_9232 = {_T_9223,_T_9076,_T_9073,_T_9070,_T_9067,_T_9064,_T_9061,_T_9058,_T_9055,_T_9052}; // @[Cat.scala 29:58]
  wire [54:0] _T_9241 = {_T_9232,_T_9049,_T_9046,_T_9043,_T_9040,_T_9037,_T_9034,_T_9031,_T_9028,_T_9025}; // @[Cat.scala 29:58]
  wire [62:0] _T_9249 = {_T_9241,_T_9022,_T_9019,_T_9016,_T_9013,_T_9010,_T_9007,_T_9004,_T_9001}; // @[Cat.scala 29:58]
  wire  _T_9317 = io_multiplicand[0] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9320 = io_multiplicand[1] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9323 = io_multiplicand[2] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9326 = io_multiplicand[3] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9329 = io_multiplicand[4] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9332 = io_multiplicand[5] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9335 = io_multiplicand[6] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9338 = io_multiplicand[7] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9341 = io_multiplicand[8] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9344 = io_multiplicand[9] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9347 = io_multiplicand[10] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9350 = io_multiplicand[11] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9353 = io_multiplicand[12] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9356 = io_multiplicand[13] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9359 = io_multiplicand[14] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9362 = io_multiplicand[15] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9365 = io_multiplicand[16] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9368 = io_multiplicand[17] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9371 = io_multiplicand[18] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9374 = io_multiplicand[19] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9377 = io_multiplicand[20] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9380 = io_multiplicand[21] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9383 = io_multiplicand[22] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9386 = io_multiplicand[23] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9389 = io_multiplicand[24] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9392 = io_multiplicand[25] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9395 = io_multiplicand[26] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9398 = io_multiplicand[27] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9401 = io_multiplicand[28] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9404 = io_multiplicand[29] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9407 = io_multiplicand[30] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9410 = io_multiplicand[31] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9413 = io_multiplicand[32] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9416 = io_multiplicand[33] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9419 = io_multiplicand[34] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9422 = io_multiplicand[35] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9425 = io_multiplicand[36] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9428 = io_multiplicand[37] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9431 = io_multiplicand[38] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9434 = io_multiplicand[39] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9437 = io_multiplicand[40] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9440 = io_multiplicand[41] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9443 = io_multiplicand[42] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9446 = io_multiplicand[43] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9449 = io_multiplicand[44] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9452 = io_multiplicand[45] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9455 = io_multiplicand[46] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9458 = io_multiplicand[47] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9461 = io_multiplicand[48] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9464 = io_multiplicand[49] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9467 = io_multiplicand[50] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9470 = io_multiplicand[51] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9473 = io_multiplicand[52] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9476 = io_multiplicand[53] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9479 = io_multiplicand[54] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9482 = io_multiplicand[55] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9485 = io_multiplicand[56] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9488 = io_multiplicand[57] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9491 = io_multiplicand[58] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9494 = io_multiplicand[59] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9497 = io_multiplicand[60] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9500 = io_multiplicand[61] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9503 = io_multiplicand[62] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire  _T_9506 = io_multiplicand[63] & io_multiplier[29]; // @[partialprod.scala 16:36]
  wire [9:0] _T_9515 = {_T_9506,_T_9503,_T_9500,_T_9497,_T_9494,_T_9491,_T_9488,_T_9485,_T_9482,_T_9479}; // @[Cat.scala 29:58]
  wire [18:0] _T_9524 = {_T_9515,_T_9476,_T_9473,_T_9470,_T_9467,_T_9464,_T_9461,_T_9458,_T_9455,_T_9452}; // @[Cat.scala 29:58]
  wire [27:0] _T_9533 = {_T_9524,_T_9449,_T_9446,_T_9443,_T_9440,_T_9437,_T_9434,_T_9431,_T_9428,_T_9425}; // @[Cat.scala 29:58]
  wire [36:0] _T_9542 = {_T_9533,_T_9422,_T_9419,_T_9416,_T_9413,_T_9410,_T_9407,_T_9404,_T_9401,_T_9398}; // @[Cat.scala 29:58]
  wire [45:0] _T_9551 = {_T_9542,_T_9395,_T_9392,_T_9389,_T_9386,_T_9383,_T_9380,_T_9377,_T_9374,_T_9371}; // @[Cat.scala 29:58]
  wire [54:0] _T_9560 = {_T_9551,_T_9368,_T_9365,_T_9362,_T_9359,_T_9356,_T_9353,_T_9350,_T_9347,_T_9344}; // @[Cat.scala 29:58]
  wire [62:0] _T_9568 = {_T_9560,_T_9341,_T_9338,_T_9335,_T_9332,_T_9329,_T_9326,_T_9323,_T_9320}; // @[Cat.scala 29:58]
  wire  _T_9636 = io_multiplicand[0] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9639 = io_multiplicand[1] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9642 = io_multiplicand[2] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9645 = io_multiplicand[3] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9648 = io_multiplicand[4] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9651 = io_multiplicand[5] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9654 = io_multiplicand[6] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9657 = io_multiplicand[7] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9660 = io_multiplicand[8] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9663 = io_multiplicand[9] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9666 = io_multiplicand[10] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9669 = io_multiplicand[11] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9672 = io_multiplicand[12] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9675 = io_multiplicand[13] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9678 = io_multiplicand[14] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9681 = io_multiplicand[15] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9684 = io_multiplicand[16] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9687 = io_multiplicand[17] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9690 = io_multiplicand[18] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9693 = io_multiplicand[19] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9696 = io_multiplicand[20] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9699 = io_multiplicand[21] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9702 = io_multiplicand[22] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9705 = io_multiplicand[23] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9708 = io_multiplicand[24] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9711 = io_multiplicand[25] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9714 = io_multiplicand[26] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9717 = io_multiplicand[27] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9720 = io_multiplicand[28] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9723 = io_multiplicand[29] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9726 = io_multiplicand[30] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9729 = io_multiplicand[31] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9732 = io_multiplicand[32] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9735 = io_multiplicand[33] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9738 = io_multiplicand[34] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9741 = io_multiplicand[35] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9744 = io_multiplicand[36] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9747 = io_multiplicand[37] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9750 = io_multiplicand[38] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9753 = io_multiplicand[39] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9756 = io_multiplicand[40] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9759 = io_multiplicand[41] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9762 = io_multiplicand[42] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9765 = io_multiplicand[43] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9768 = io_multiplicand[44] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9771 = io_multiplicand[45] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9774 = io_multiplicand[46] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9777 = io_multiplicand[47] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9780 = io_multiplicand[48] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9783 = io_multiplicand[49] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9786 = io_multiplicand[50] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9789 = io_multiplicand[51] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9792 = io_multiplicand[52] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9795 = io_multiplicand[53] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9798 = io_multiplicand[54] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9801 = io_multiplicand[55] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9804 = io_multiplicand[56] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9807 = io_multiplicand[57] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9810 = io_multiplicand[58] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9813 = io_multiplicand[59] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9816 = io_multiplicand[60] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9819 = io_multiplicand[61] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9822 = io_multiplicand[62] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire  _T_9825 = io_multiplicand[63] & io_multiplier[30]; // @[partialprod.scala 16:36]
  wire [9:0] _T_9834 = {_T_9825,_T_9822,_T_9819,_T_9816,_T_9813,_T_9810,_T_9807,_T_9804,_T_9801,_T_9798}; // @[Cat.scala 29:58]
  wire [18:0] _T_9843 = {_T_9834,_T_9795,_T_9792,_T_9789,_T_9786,_T_9783,_T_9780,_T_9777,_T_9774,_T_9771}; // @[Cat.scala 29:58]
  wire [27:0] _T_9852 = {_T_9843,_T_9768,_T_9765,_T_9762,_T_9759,_T_9756,_T_9753,_T_9750,_T_9747,_T_9744}; // @[Cat.scala 29:58]
  wire [36:0] _T_9861 = {_T_9852,_T_9741,_T_9738,_T_9735,_T_9732,_T_9729,_T_9726,_T_9723,_T_9720,_T_9717}; // @[Cat.scala 29:58]
  wire [45:0] _T_9870 = {_T_9861,_T_9714,_T_9711,_T_9708,_T_9705,_T_9702,_T_9699,_T_9696,_T_9693,_T_9690}; // @[Cat.scala 29:58]
  wire [54:0] _T_9879 = {_T_9870,_T_9687,_T_9684,_T_9681,_T_9678,_T_9675,_T_9672,_T_9669,_T_9666,_T_9663}; // @[Cat.scala 29:58]
  wire [62:0] _T_9887 = {_T_9879,_T_9660,_T_9657,_T_9654,_T_9651,_T_9648,_T_9645,_T_9642,_T_9639}; // @[Cat.scala 29:58]
  wire  _T_9955 = io_multiplicand[0] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_9958 = io_multiplicand[1] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_9961 = io_multiplicand[2] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_9964 = io_multiplicand[3] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_9967 = io_multiplicand[4] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_9970 = io_multiplicand[5] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_9973 = io_multiplicand[6] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_9976 = io_multiplicand[7] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_9979 = io_multiplicand[8] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_9982 = io_multiplicand[9] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_9985 = io_multiplicand[10] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_9988 = io_multiplicand[11] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_9991 = io_multiplicand[12] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_9994 = io_multiplicand[13] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_9997 = io_multiplicand[14] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10000 = io_multiplicand[15] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10003 = io_multiplicand[16] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10006 = io_multiplicand[17] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10009 = io_multiplicand[18] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10012 = io_multiplicand[19] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10015 = io_multiplicand[20] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10018 = io_multiplicand[21] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10021 = io_multiplicand[22] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10024 = io_multiplicand[23] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10027 = io_multiplicand[24] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10030 = io_multiplicand[25] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10033 = io_multiplicand[26] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10036 = io_multiplicand[27] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10039 = io_multiplicand[28] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10042 = io_multiplicand[29] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10045 = io_multiplicand[30] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10048 = io_multiplicand[31] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10051 = io_multiplicand[32] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10054 = io_multiplicand[33] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10057 = io_multiplicand[34] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10060 = io_multiplicand[35] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10063 = io_multiplicand[36] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10066 = io_multiplicand[37] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10069 = io_multiplicand[38] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10072 = io_multiplicand[39] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10075 = io_multiplicand[40] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10078 = io_multiplicand[41] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10081 = io_multiplicand[42] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10084 = io_multiplicand[43] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10087 = io_multiplicand[44] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10090 = io_multiplicand[45] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10093 = io_multiplicand[46] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10096 = io_multiplicand[47] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10099 = io_multiplicand[48] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10102 = io_multiplicand[49] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10105 = io_multiplicand[50] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10108 = io_multiplicand[51] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10111 = io_multiplicand[52] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10114 = io_multiplicand[53] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10117 = io_multiplicand[54] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10120 = io_multiplicand[55] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10123 = io_multiplicand[56] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10126 = io_multiplicand[57] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10129 = io_multiplicand[58] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10132 = io_multiplicand[59] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10135 = io_multiplicand[60] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10138 = io_multiplicand[61] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10141 = io_multiplicand[62] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire  _T_10144 = io_multiplicand[63] & io_multiplier[31]; // @[partialprod.scala 16:36]
  wire [9:0] _T_10153 = {_T_10144,_T_10141,_T_10138,_T_10135,_T_10132,_T_10129,_T_10126,_T_10123,_T_10120,_T_10117}; // @[Cat.scala 29:58]
  wire [18:0] _T_10162 = {_T_10153,_T_10114,_T_10111,_T_10108,_T_10105,_T_10102,_T_10099,_T_10096,_T_10093,_T_10090}; // @[Cat.scala 29:58]
  wire [27:0] _T_10171 = {_T_10162,_T_10087,_T_10084,_T_10081,_T_10078,_T_10075,_T_10072,_T_10069,_T_10066,_T_10063}; // @[Cat.scala 29:58]
  wire [36:0] _T_10180 = {_T_10171,_T_10060,_T_10057,_T_10054,_T_10051,_T_10048,_T_10045,_T_10042,_T_10039,_T_10036}; // @[Cat.scala 29:58]
  wire [45:0] _T_10189 = {_T_10180,_T_10033,_T_10030,_T_10027,_T_10024,_T_10021,_T_10018,_T_10015,_T_10012,_T_10009}; // @[Cat.scala 29:58]
  wire [54:0] _T_10198 = {_T_10189,_T_10006,_T_10003,_T_10000,_T_9997,_T_9994,_T_9991,_T_9988,_T_9985,_T_9982}; // @[Cat.scala 29:58]
  wire [62:0] _T_10206 = {_T_10198,_T_9979,_T_9976,_T_9973,_T_9970,_T_9967,_T_9964,_T_9961,_T_9958}; // @[Cat.scala 29:58]
  wire  _T_10274 = io_multiplicand[0] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10277 = io_multiplicand[1] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10280 = io_multiplicand[2] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10283 = io_multiplicand[3] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10286 = io_multiplicand[4] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10289 = io_multiplicand[5] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10292 = io_multiplicand[6] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10295 = io_multiplicand[7] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10298 = io_multiplicand[8] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10301 = io_multiplicand[9] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10304 = io_multiplicand[10] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10307 = io_multiplicand[11] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10310 = io_multiplicand[12] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10313 = io_multiplicand[13] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10316 = io_multiplicand[14] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10319 = io_multiplicand[15] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10322 = io_multiplicand[16] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10325 = io_multiplicand[17] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10328 = io_multiplicand[18] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10331 = io_multiplicand[19] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10334 = io_multiplicand[20] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10337 = io_multiplicand[21] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10340 = io_multiplicand[22] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10343 = io_multiplicand[23] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10346 = io_multiplicand[24] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10349 = io_multiplicand[25] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10352 = io_multiplicand[26] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10355 = io_multiplicand[27] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10358 = io_multiplicand[28] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10361 = io_multiplicand[29] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10364 = io_multiplicand[30] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10367 = io_multiplicand[31] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10370 = io_multiplicand[32] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10373 = io_multiplicand[33] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10376 = io_multiplicand[34] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10379 = io_multiplicand[35] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10382 = io_multiplicand[36] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10385 = io_multiplicand[37] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10388 = io_multiplicand[38] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10391 = io_multiplicand[39] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10394 = io_multiplicand[40] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10397 = io_multiplicand[41] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10400 = io_multiplicand[42] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10403 = io_multiplicand[43] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10406 = io_multiplicand[44] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10409 = io_multiplicand[45] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10412 = io_multiplicand[46] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10415 = io_multiplicand[47] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10418 = io_multiplicand[48] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10421 = io_multiplicand[49] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10424 = io_multiplicand[50] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10427 = io_multiplicand[51] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10430 = io_multiplicand[52] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10433 = io_multiplicand[53] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10436 = io_multiplicand[54] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10439 = io_multiplicand[55] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10442 = io_multiplicand[56] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10445 = io_multiplicand[57] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10448 = io_multiplicand[58] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10451 = io_multiplicand[59] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10454 = io_multiplicand[60] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10457 = io_multiplicand[61] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10460 = io_multiplicand[62] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire  _T_10463 = io_multiplicand[63] & io_multiplier[32]; // @[partialprod.scala 16:36]
  wire [9:0] _T_10472 = {_T_10463,_T_10460,_T_10457,_T_10454,_T_10451,_T_10448,_T_10445,_T_10442,_T_10439,_T_10436}; // @[Cat.scala 29:58]
  wire [18:0] _T_10481 = {_T_10472,_T_10433,_T_10430,_T_10427,_T_10424,_T_10421,_T_10418,_T_10415,_T_10412,_T_10409}; // @[Cat.scala 29:58]
  wire [27:0] _T_10490 = {_T_10481,_T_10406,_T_10403,_T_10400,_T_10397,_T_10394,_T_10391,_T_10388,_T_10385,_T_10382}; // @[Cat.scala 29:58]
  wire [36:0] _T_10499 = {_T_10490,_T_10379,_T_10376,_T_10373,_T_10370,_T_10367,_T_10364,_T_10361,_T_10358,_T_10355}; // @[Cat.scala 29:58]
  wire [45:0] _T_10508 = {_T_10499,_T_10352,_T_10349,_T_10346,_T_10343,_T_10340,_T_10337,_T_10334,_T_10331,_T_10328}; // @[Cat.scala 29:58]
  wire [54:0] _T_10517 = {_T_10508,_T_10325,_T_10322,_T_10319,_T_10316,_T_10313,_T_10310,_T_10307,_T_10304,_T_10301}; // @[Cat.scala 29:58]
  wire [62:0] _T_10525 = {_T_10517,_T_10298,_T_10295,_T_10292,_T_10289,_T_10286,_T_10283,_T_10280,_T_10277}; // @[Cat.scala 29:58]
  wire  _T_10593 = io_multiplicand[0] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10596 = io_multiplicand[1] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10599 = io_multiplicand[2] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10602 = io_multiplicand[3] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10605 = io_multiplicand[4] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10608 = io_multiplicand[5] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10611 = io_multiplicand[6] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10614 = io_multiplicand[7] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10617 = io_multiplicand[8] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10620 = io_multiplicand[9] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10623 = io_multiplicand[10] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10626 = io_multiplicand[11] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10629 = io_multiplicand[12] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10632 = io_multiplicand[13] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10635 = io_multiplicand[14] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10638 = io_multiplicand[15] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10641 = io_multiplicand[16] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10644 = io_multiplicand[17] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10647 = io_multiplicand[18] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10650 = io_multiplicand[19] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10653 = io_multiplicand[20] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10656 = io_multiplicand[21] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10659 = io_multiplicand[22] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10662 = io_multiplicand[23] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10665 = io_multiplicand[24] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10668 = io_multiplicand[25] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10671 = io_multiplicand[26] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10674 = io_multiplicand[27] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10677 = io_multiplicand[28] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10680 = io_multiplicand[29] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10683 = io_multiplicand[30] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10686 = io_multiplicand[31] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10689 = io_multiplicand[32] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10692 = io_multiplicand[33] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10695 = io_multiplicand[34] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10698 = io_multiplicand[35] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10701 = io_multiplicand[36] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10704 = io_multiplicand[37] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10707 = io_multiplicand[38] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10710 = io_multiplicand[39] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10713 = io_multiplicand[40] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10716 = io_multiplicand[41] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10719 = io_multiplicand[42] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10722 = io_multiplicand[43] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10725 = io_multiplicand[44] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10728 = io_multiplicand[45] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10731 = io_multiplicand[46] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10734 = io_multiplicand[47] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10737 = io_multiplicand[48] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10740 = io_multiplicand[49] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10743 = io_multiplicand[50] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10746 = io_multiplicand[51] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10749 = io_multiplicand[52] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10752 = io_multiplicand[53] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10755 = io_multiplicand[54] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10758 = io_multiplicand[55] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10761 = io_multiplicand[56] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10764 = io_multiplicand[57] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10767 = io_multiplicand[58] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10770 = io_multiplicand[59] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10773 = io_multiplicand[60] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10776 = io_multiplicand[61] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10779 = io_multiplicand[62] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire  _T_10782 = io_multiplicand[63] & io_multiplier[33]; // @[partialprod.scala 16:36]
  wire [9:0] _T_10791 = {_T_10782,_T_10779,_T_10776,_T_10773,_T_10770,_T_10767,_T_10764,_T_10761,_T_10758,_T_10755}; // @[Cat.scala 29:58]
  wire [18:0] _T_10800 = {_T_10791,_T_10752,_T_10749,_T_10746,_T_10743,_T_10740,_T_10737,_T_10734,_T_10731,_T_10728}; // @[Cat.scala 29:58]
  wire [27:0] _T_10809 = {_T_10800,_T_10725,_T_10722,_T_10719,_T_10716,_T_10713,_T_10710,_T_10707,_T_10704,_T_10701}; // @[Cat.scala 29:58]
  wire [36:0] _T_10818 = {_T_10809,_T_10698,_T_10695,_T_10692,_T_10689,_T_10686,_T_10683,_T_10680,_T_10677,_T_10674}; // @[Cat.scala 29:58]
  wire [45:0] _T_10827 = {_T_10818,_T_10671,_T_10668,_T_10665,_T_10662,_T_10659,_T_10656,_T_10653,_T_10650,_T_10647}; // @[Cat.scala 29:58]
  wire [54:0] _T_10836 = {_T_10827,_T_10644,_T_10641,_T_10638,_T_10635,_T_10632,_T_10629,_T_10626,_T_10623,_T_10620}; // @[Cat.scala 29:58]
  wire [62:0] _T_10844 = {_T_10836,_T_10617,_T_10614,_T_10611,_T_10608,_T_10605,_T_10602,_T_10599,_T_10596}; // @[Cat.scala 29:58]
  wire  _T_10912 = io_multiplicand[0] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10915 = io_multiplicand[1] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10918 = io_multiplicand[2] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10921 = io_multiplicand[3] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10924 = io_multiplicand[4] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10927 = io_multiplicand[5] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10930 = io_multiplicand[6] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10933 = io_multiplicand[7] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10936 = io_multiplicand[8] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10939 = io_multiplicand[9] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10942 = io_multiplicand[10] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10945 = io_multiplicand[11] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10948 = io_multiplicand[12] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10951 = io_multiplicand[13] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10954 = io_multiplicand[14] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10957 = io_multiplicand[15] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10960 = io_multiplicand[16] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10963 = io_multiplicand[17] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10966 = io_multiplicand[18] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10969 = io_multiplicand[19] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10972 = io_multiplicand[20] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10975 = io_multiplicand[21] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10978 = io_multiplicand[22] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10981 = io_multiplicand[23] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10984 = io_multiplicand[24] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10987 = io_multiplicand[25] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10990 = io_multiplicand[26] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10993 = io_multiplicand[27] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10996 = io_multiplicand[28] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_10999 = io_multiplicand[29] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11002 = io_multiplicand[30] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11005 = io_multiplicand[31] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11008 = io_multiplicand[32] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11011 = io_multiplicand[33] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11014 = io_multiplicand[34] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11017 = io_multiplicand[35] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11020 = io_multiplicand[36] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11023 = io_multiplicand[37] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11026 = io_multiplicand[38] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11029 = io_multiplicand[39] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11032 = io_multiplicand[40] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11035 = io_multiplicand[41] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11038 = io_multiplicand[42] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11041 = io_multiplicand[43] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11044 = io_multiplicand[44] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11047 = io_multiplicand[45] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11050 = io_multiplicand[46] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11053 = io_multiplicand[47] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11056 = io_multiplicand[48] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11059 = io_multiplicand[49] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11062 = io_multiplicand[50] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11065 = io_multiplicand[51] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11068 = io_multiplicand[52] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11071 = io_multiplicand[53] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11074 = io_multiplicand[54] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11077 = io_multiplicand[55] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11080 = io_multiplicand[56] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11083 = io_multiplicand[57] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11086 = io_multiplicand[58] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11089 = io_multiplicand[59] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11092 = io_multiplicand[60] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11095 = io_multiplicand[61] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11098 = io_multiplicand[62] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire  _T_11101 = io_multiplicand[63] & io_multiplier[34]; // @[partialprod.scala 16:36]
  wire [9:0] _T_11110 = {_T_11101,_T_11098,_T_11095,_T_11092,_T_11089,_T_11086,_T_11083,_T_11080,_T_11077,_T_11074}; // @[Cat.scala 29:58]
  wire [18:0] _T_11119 = {_T_11110,_T_11071,_T_11068,_T_11065,_T_11062,_T_11059,_T_11056,_T_11053,_T_11050,_T_11047}; // @[Cat.scala 29:58]
  wire [27:0] _T_11128 = {_T_11119,_T_11044,_T_11041,_T_11038,_T_11035,_T_11032,_T_11029,_T_11026,_T_11023,_T_11020}; // @[Cat.scala 29:58]
  wire [36:0] _T_11137 = {_T_11128,_T_11017,_T_11014,_T_11011,_T_11008,_T_11005,_T_11002,_T_10999,_T_10996,_T_10993}; // @[Cat.scala 29:58]
  wire [45:0] _T_11146 = {_T_11137,_T_10990,_T_10987,_T_10984,_T_10981,_T_10978,_T_10975,_T_10972,_T_10969,_T_10966}; // @[Cat.scala 29:58]
  wire [54:0] _T_11155 = {_T_11146,_T_10963,_T_10960,_T_10957,_T_10954,_T_10951,_T_10948,_T_10945,_T_10942,_T_10939}; // @[Cat.scala 29:58]
  wire [62:0] _T_11163 = {_T_11155,_T_10936,_T_10933,_T_10930,_T_10927,_T_10924,_T_10921,_T_10918,_T_10915}; // @[Cat.scala 29:58]
  wire  _T_11231 = io_multiplicand[0] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11234 = io_multiplicand[1] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11237 = io_multiplicand[2] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11240 = io_multiplicand[3] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11243 = io_multiplicand[4] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11246 = io_multiplicand[5] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11249 = io_multiplicand[6] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11252 = io_multiplicand[7] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11255 = io_multiplicand[8] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11258 = io_multiplicand[9] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11261 = io_multiplicand[10] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11264 = io_multiplicand[11] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11267 = io_multiplicand[12] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11270 = io_multiplicand[13] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11273 = io_multiplicand[14] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11276 = io_multiplicand[15] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11279 = io_multiplicand[16] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11282 = io_multiplicand[17] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11285 = io_multiplicand[18] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11288 = io_multiplicand[19] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11291 = io_multiplicand[20] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11294 = io_multiplicand[21] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11297 = io_multiplicand[22] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11300 = io_multiplicand[23] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11303 = io_multiplicand[24] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11306 = io_multiplicand[25] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11309 = io_multiplicand[26] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11312 = io_multiplicand[27] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11315 = io_multiplicand[28] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11318 = io_multiplicand[29] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11321 = io_multiplicand[30] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11324 = io_multiplicand[31] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11327 = io_multiplicand[32] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11330 = io_multiplicand[33] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11333 = io_multiplicand[34] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11336 = io_multiplicand[35] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11339 = io_multiplicand[36] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11342 = io_multiplicand[37] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11345 = io_multiplicand[38] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11348 = io_multiplicand[39] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11351 = io_multiplicand[40] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11354 = io_multiplicand[41] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11357 = io_multiplicand[42] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11360 = io_multiplicand[43] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11363 = io_multiplicand[44] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11366 = io_multiplicand[45] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11369 = io_multiplicand[46] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11372 = io_multiplicand[47] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11375 = io_multiplicand[48] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11378 = io_multiplicand[49] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11381 = io_multiplicand[50] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11384 = io_multiplicand[51] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11387 = io_multiplicand[52] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11390 = io_multiplicand[53] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11393 = io_multiplicand[54] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11396 = io_multiplicand[55] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11399 = io_multiplicand[56] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11402 = io_multiplicand[57] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11405 = io_multiplicand[58] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11408 = io_multiplicand[59] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11411 = io_multiplicand[60] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11414 = io_multiplicand[61] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11417 = io_multiplicand[62] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire  _T_11420 = io_multiplicand[63] & io_multiplier[35]; // @[partialprod.scala 16:36]
  wire [9:0] _T_11429 = {_T_11420,_T_11417,_T_11414,_T_11411,_T_11408,_T_11405,_T_11402,_T_11399,_T_11396,_T_11393}; // @[Cat.scala 29:58]
  wire [18:0] _T_11438 = {_T_11429,_T_11390,_T_11387,_T_11384,_T_11381,_T_11378,_T_11375,_T_11372,_T_11369,_T_11366}; // @[Cat.scala 29:58]
  wire [27:0] _T_11447 = {_T_11438,_T_11363,_T_11360,_T_11357,_T_11354,_T_11351,_T_11348,_T_11345,_T_11342,_T_11339}; // @[Cat.scala 29:58]
  wire [36:0] _T_11456 = {_T_11447,_T_11336,_T_11333,_T_11330,_T_11327,_T_11324,_T_11321,_T_11318,_T_11315,_T_11312}; // @[Cat.scala 29:58]
  wire [45:0] _T_11465 = {_T_11456,_T_11309,_T_11306,_T_11303,_T_11300,_T_11297,_T_11294,_T_11291,_T_11288,_T_11285}; // @[Cat.scala 29:58]
  wire [54:0] _T_11474 = {_T_11465,_T_11282,_T_11279,_T_11276,_T_11273,_T_11270,_T_11267,_T_11264,_T_11261,_T_11258}; // @[Cat.scala 29:58]
  wire [62:0] _T_11482 = {_T_11474,_T_11255,_T_11252,_T_11249,_T_11246,_T_11243,_T_11240,_T_11237,_T_11234}; // @[Cat.scala 29:58]
  wire  _T_11550 = io_multiplicand[0] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11553 = io_multiplicand[1] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11556 = io_multiplicand[2] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11559 = io_multiplicand[3] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11562 = io_multiplicand[4] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11565 = io_multiplicand[5] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11568 = io_multiplicand[6] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11571 = io_multiplicand[7] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11574 = io_multiplicand[8] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11577 = io_multiplicand[9] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11580 = io_multiplicand[10] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11583 = io_multiplicand[11] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11586 = io_multiplicand[12] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11589 = io_multiplicand[13] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11592 = io_multiplicand[14] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11595 = io_multiplicand[15] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11598 = io_multiplicand[16] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11601 = io_multiplicand[17] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11604 = io_multiplicand[18] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11607 = io_multiplicand[19] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11610 = io_multiplicand[20] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11613 = io_multiplicand[21] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11616 = io_multiplicand[22] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11619 = io_multiplicand[23] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11622 = io_multiplicand[24] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11625 = io_multiplicand[25] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11628 = io_multiplicand[26] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11631 = io_multiplicand[27] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11634 = io_multiplicand[28] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11637 = io_multiplicand[29] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11640 = io_multiplicand[30] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11643 = io_multiplicand[31] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11646 = io_multiplicand[32] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11649 = io_multiplicand[33] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11652 = io_multiplicand[34] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11655 = io_multiplicand[35] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11658 = io_multiplicand[36] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11661 = io_multiplicand[37] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11664 = io_multiplicand[38] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11667 = io_multiplicand[39] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11670 = io_multiplicand[40] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11673 = io_multiplicand[41] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11676 = io_multiplicand[42] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11679 = io_multiplicand[43] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11682 = io_multiplicand[44] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11685 = io_multiplicand[45] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11688 = io_multiplicand[46] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11691 = io_multiplicand[47] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11694 = io_multiplicand[48] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11697 = io_multiplicand[49] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11700 = io_multiplicand[50] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11703 = io_multiplicand[51] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11706 = io_multiplicand[52] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11709 = io_multiplicand[53] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11712 = io_multiplicand[54] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11715 = io_multiplicand[55] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11718 = io_multiplicand[56] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11721 = io_multiplicand[57] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11724 = io_multiplicand[58] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11727 = io_multiplicand[59] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11730 = io_multiplicand[60] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11733 = io_multiplicand[61] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11736 = io_multiplicand[62] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire  _T_11739 = io_multiplicand[63] & io_multiplier[36]; // @[partialprod.scala 16:36]
  wire [9:0] _T_11748 = {_T_11739,_T_11736,_T_11733,_T_11730,_T_11727,_T_11724,_T_11721,_T_11718,_T_11715,_T_11712}; // @[Cat.scala 29:58]
  wire [18:0] _T_11757 = {_T_11748,_T_11709,_T_11706,_T_11703,_T_11700,_T_11697,_T_11694,_T_11691,_T_11688,_T_11685}; // @[Cat.scala 29:58]
  wire [27:0] _T_11766 = {_T_11757,_T_11682,_T_11679,_T_11676,_T_11673,_T_11670,_T_11667,_T_11664,_T_11661,_T_11658}; // @[Cat.scala 29:58]
  wire [36:0] _T_11775 = {_T_11766,_T_11655,_T_11652,_T_11649,_T_11646,_T_11643,_T_11640,_T_11637,_T_11634,_T_11631}; // @[Cat.scala 29:58]
  wire [45:0] _T_11784 = {_T_11775,_T_11628,_T_11625,_T_11622,_T_11619,_T_11616,_T_11613,_T_11610,_T_11607,_T_11604}; // @[Cat.scala 29:58]
  wire [54:0] _T_11793 = {_T_11784,_T_11601,_T_11598,_T_11595,_T_11592,_T_11589,_T_11586,_T_11583,_T_11580,_T_11577}; // @[Cat.scala 29:58]
  wire [62:0] _T_11801 = {_T_11793,_T_11574,_T_11571,_T_11568,_T_11565,_T_11562,_T_11559,_T_11556,_T_11553}; // @[Cat.scala 29:58]
  wire  _T_11869 = io_multiplicand[0] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11872 = io_multiplicand[1] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11875 = io_multiplicand[2] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11878 = io_multiplicand[3] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11881 = io_multiplicand[4] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11884 = io_multiplicand[5] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11887 = io_multiplicand[6] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11890 = io_multiplicand[7] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11893 = io_multiplicand[8] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11896 = io_multiplicand[9] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11899 = io_multiplicand[10] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11902 = io_multiplicand[11] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11905 = io_multiplicand[12] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11908 = io_multiplicand[13] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11911 = io_multiplicand[14] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11914 = io_multiplicand[15] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11917 = io_multiplicand[16] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11920 = io_multiplicand[17] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11923 = io_multiplicand[18] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11926 = io_multiplicand[19] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11929 = io_multiplicand[20] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11932 = io_multiplicand[21] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11935 = io_multiplicand[22] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11938 = io_multiplicand[23] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11941 = io_multiplicand[24] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11944 = io_multiplicand[25] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11947 = io_multiplicand[26] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11950 = io_multiplicand[27] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11953 = io_multiplicand[28] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11956 = io_multiplicand[29] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11959 = io_multiplicand[30] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11962 = io_multiplicand[31] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11965 = io_multiplicand[32] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11968 = io_multiplicand[33] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11971 = io_multiplicand[34] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11974 = io_multiplicand[35] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11977 = io_multiplicand[36] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11980 = io_multiplicand[37] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11983 = io_multiplicand[38] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11986 = io_multiplicand[39] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11989 = io_multiplicand[40] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11992 = io_multiplicand[41] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11995 = io_multiplicand[42] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_11998 = io_multiplicand[43] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12001 = io_multiplicand[44] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12004 = io_multiplicand[45] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12007 = io_multiplicand[46] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12010 = io_multiplicand[47] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12013 = io_multiplicand[48] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12016 = io_multiplicand[49] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12019 = io_multiplicand[50] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12022 = io_multiplicand[51] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12025 = io_multiplicand[52] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12028 = io_multiplicand[53] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12031 = io_multiplicand[54] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12034 = io_multiplicand[55] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12037 = io_multiplicand[56] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12040 = io_multiplicand[57] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12043 = io_multiplicand[58] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12046 = io_multiplicand[59] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12049 = io_multiplicand[60] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12052 = io_multiplicand[61] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12055 = io_multiplicand[62] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire  _T_12058 = io_multiplicand[63] & io_multiplier[37]; // @[partialprod.scala 16:36]
  wire [9:0] _T_12067 = {_T_12058,_T_12055,_T_12052,_T_12049,_T_12046,_T_12043,_T_12040,_T_12037,_T_12034,_T_12031}; // @[Cat.scala 29:58]
  wire [18:0] _T_12076 = {_T_12067,_T_12028,_T_12025,_T_12022,_T_12019,_T_12016,_T_12013,_T_12010,_T_12007,_T_12004}; // @[Cat.scala 29:58]
  wire [27:0] _T_12085 = {_T_12076,_T_12001,_T_11998,_T_11995,_T_11992,_T_11989,_T_11986,_T_11983,_T_11980,_T_11977}; // @[Cat.scala 29:58]
  wire [36:0] _T_12094 = {_T_12085,_T_11974,_T_11971,_T_11968,_T_11965,_T_11962,_T_11959,_T_11956,_T_11953,_T_11950}; // @[Cat.scala 29:58]
  wire [45:0] _T_12103 = {_T_12094,_T_11947,_T_11944,_T_11941,_T_11938,_T_11935,_T_11932,_T_11929,_T_11926,_T_11923}; // @[Cat.scala 29:58]
  wire [54:0] _T_12112 = {_T_12103,_T_11920,_T_11917,_T_11914,_T_11911,_T_11908,_T_11905,_T_11902,_T_11899,_T_11896}; // @[Cat.scala 29:58]
  wire [62:0] _T_12120 = {_T_12112,_T_11893,_T_11890,_T_11887,_T_11884,_T_11881,_T_11878,_T_11875,_T_11872}; // @[Cat.scala 29:58]
  wire  _T_12188 = io_multiplicand[0] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12191 = io_multiplicand[1] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12194 = io_multiplicand[2] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12197 = io_multiplicand[3] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12200 = io_multiplicand[4] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12203 = io_multiplicand[5] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12206 = io_multiplicand[6] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12209 = io_multiplicand[7] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12212 = io_multiplicand[8] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12215 = io_multiplicand[9] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12218 = io_multiplicand[10] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12221 = io_multiplicand[11] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12224 = io_multiplicand[12] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12227 = io_multiplicand[13] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12230 = io_multiplicand[14] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12233 = io_multiplicand[15] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12236 = io_multiplicand[16] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12239 = io_multiplicand[17] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12242 = io_multiplicand[18] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12245 = io_multiplicand[19] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12248 = io_multiplicand[20] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12251 = io_multiplicand[21] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12254 = io_multiplicand[22] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12257 = io_multiplicand[23] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12260 = io_multiplicand[24] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12263 = io_multiplicand[25] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12266 = io_multiplicand[26] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12269 = io_multiplicand[27] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12272 = io_multiplicand[28] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12275 = io_multiplicand[29] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12278 = io_multiplicand[30] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12281 = io_multiplicand[31] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12284 = io_multiplicand[32] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12287 = io_multiplicand[33] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12290 = io_multiplicand[34] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12293 = io_multiplicand[35] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12296 = io_multiplicand[36] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12299 = io_multiplicand[37] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12302 = io_multiplicand[38] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12305 = io_multiplicand[39] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12308 = io_multiplicand[40] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12311 = io_multiplicand[41] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12314 = io_multiplicand[42] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12317 = io_multiplicand[43] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12320 = io_multiplicand[44] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12323 = io_multiplicand[45] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12326 = io_multiplicand[46] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12329 = io_multiplicand[47] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12332 = io_multiplicand[48] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12335 = io_multiplicand[49] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12338 = io_multiplicand[50] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12341 = io_multiplicand[51] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12344 = io_multiplicand[52] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12347 = io_multiplicand[53] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12350 = io_multiplicand[54] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12353 = io_multiplicand[55] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12356 = io_multiplicand[56] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12359 = io_multiplicand[57] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12362 = io_multiplicand[58] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12365 = io_multiplicand[59] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12368 = io_multiplicand[60] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12371 = io_multiplicand[61] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12374 = io_multiplicand[62] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire  _T_12377 = io_multiplicand[63] & io_multiplier[38]; // @[partialprod.scala 16:36]
  wire [9:0] _T_12386 = {_T_12377,_T_12374,_T_12371,_T_12368,_T_12365,_T_12362,_T_12359,_T_12356,_T_12353,_T_12350}; // @[Cat.scala 29:58]
  wire [18:0] _T_12395 = {_T_12386,_T_12347,_T_12344,_T_12341,_T_12338,_T_12335,_T_12332,_T_12329,_T_12326,_T_12323}; // @[Cat.scala 29:58]
  wire [27:0] _T_12404 = {_T_12395,_T_12320,_T_12317,_T_12314,_T_12311,_T_12308,_T_12305,_T_12302,_T_12299,_T_12296}; // @[Cat.scala 29:58]
  wire [36:0] _T_12413 = {_T_12404,_T_12293,_T_12290,_T_12287,_T_12284,_T_12281,_T_12278,_T_12275,_T_12272,_T_12269}; // @[Cat.scala 29:58]
  wire [45:0] _T_12422 = {_T_12413,_T_12266,_T_12263,_T_12260,_T_12257,_T_12254,_T_12251,_T_12248,_T_12245,_T_12242}; // @[Cat.scala 29:58]
  wire [54:0] _T_12431 = {_T_12422,_T_12239,_T_12236,_T_12233,_T_12230,_T_12227,_T_12224,_T_12221,_T_12218,_T_12215}; // @[Cat.scala 29:58]
  wire [62:0] _T_12439 = {_T_12431,_T_12212,_T_12209,_T_12206,_T_12203,_T_12200,_T_12197,_T_12194,_T_12191}; // @[Cat.scala 29:58]
  wire  _T_12507 = io_multiplicand[0] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12510 = io_multiplicand[1] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12513 = io_multiplicand[2] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12516 = io_multiplicand[3] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12519 = io_multiplicand[4] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12522 = io_multiplicand[5] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12525 = io_multiplicand[6] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12528 = io_multiplicand[7] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12531 = io_multiplicand[8] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12534 = io_multiplicand[9] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12537 = io_multiplicand[10] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12540 = io_multiplicand[11] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12543 = io_multiplicand[12] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12546 = io_multiplicand[13] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12549 = io_multiplicand[14] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12552 = io_multiplicand[15] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12555 = io_multiplicand[16] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12558 = io_multiplicand[17] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12561 = io_multiplicand[18] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12564 = io_multiplicand[19] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12567 = io_multiplicand[20] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12570 = io_multiplicand[21] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12573 = io_multiplicand[22] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12576 = io_multiplicand[23] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12579 = io_multiplicand[24] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12582 = io_multiplicand[25] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12585 = io_multiplicand[26] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12588 = io_multiplicand[27] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12591 = io_multiplicand[28] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12594 = io_multiplicand[29] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12597 = io_multiplicand[30] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12600 = io_multiplicand[31] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12603 = io_multiplicand[32] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12606 = io_multiplicand[33] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12609 = io_multiplicand[34] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12612 = io_multiplicand[35] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12615 = io_multiplicand[36] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12618 = io_multiplicand[37] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12621 = io_multiplicand[38] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12624 = io_multiplicand[39] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12627 = io_multiplicand[40] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12630 = io_multiplicand[41] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12633 = io_multiplicand[42] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12636 = io_multiplicand[43] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12639 = io_multiplicand[44] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12642 = io_multiplicand[45] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12645 = io_multiplicand[46] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12648 = io_multiplicand[47] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12651 = io_multiplicand[48] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12654 = io_multiplicand[49] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12657 = io_multiplicand[50] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12660 = io_multiplicand[51] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12663 = io_multiplicand[52] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12666 = io_multiplicand[53] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12669 = io_multiplicand[54] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12672 = io_multiplicand[55] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12675 = io_multiplicand[56] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12678 = io_multiplicand[57] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12681 = io_multiplicand[58] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12684 = io_multiplicand[59] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12687 = io_multiplicand[60] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12690 = io_multiplicand[61] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12693 = io_multiplicand[62] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire  _T_12696 = io_multiplicand[63] & io_multiplier[39]; // @[partialprod.scala 16:36]
  wire [9:0] _T_12705 = {_T_12696,_T_12693,_T_12690,_T_12687,_T_12684,_T_12681,_T_12678,_T_12675,_T_12672,_T_12669}; // @[Cat.scala 29:58]
  wire [18:0] _T_12714 = {_T_12705,_T_12666,_T_12663,_T_12660,_T_12657,_T_12654,_T_12651,_T_12648,_T_12645,_T_12642}; // @[Cat.scala 29:58]
  wire [27:0] _T_12723 = {_T_12714,_T_12639,_T_12636,_T_12633,_T_12630,_T_12627,_T_12624,_T_12621,_T_12618,_T_12615}; // @[Cat.scala 29:58]
  wire [36:0] _T_12732 = {_T_12723,_T_12612,_T_12609,_T_12606,_T_12603,_T_12600,_T_12597,_T_12594,_T_12591,_T_12588}; // @[Cat.scala 29:58]
  wire [45:0] _T_12741 = {_T_12732,_T_12585,_T_12582,_T_12579,_T_12576,_T_12573,_T_12570,_T_12567,_T_12564,_T_12561}; // @[Cat.scala 29:58]
  wire [54:0] _T_12750 = {_T_12741,_T_12558,_T_12555,_T_12552,_T_12549,_T_12546,_T_12543,_T_12540,_T_12537,_T_12534}; // @[Cat.scala 29:58]
  wire [62:0] _T_12758 = {_T_12750,_T_12531,_T_12528,_T_12525,_T_12522,_T_12519,_T_12516,_T_12513,_T_12510}; // @[Cat.scala 29:58]
  wire  _T_12826 = io_multiplicand[0] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12829 = io_multiplicand[1] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12832 = io_multiplicand[2] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12835 = io_multiplicand[3] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12838 = io_multiplicand[4] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12841 = io_multiplicand[5] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12844 = io_multiplicand[6] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12847 = io_multiplicand[7] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12850 = io_multiplicand[8] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12853 = io_multiplicand[9] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12856 = io_multiplicand[10] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12859 = io_multiplicand[11] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12862 = io_multiplicand[12] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12865 = io_multiplicand[13] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12868 = io_multiplicand[14] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12871 = io_multiplicand[15] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12874 = io_multiplicand[16] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12877 = io_multiplicand[17] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12880 = io_multiplicand[18] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12883 = io_multiplicand[19] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12886 = io_multiplicand[20] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12889 = io_multiplicand[21] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12892 = io_multiplicand[22] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12895 = io_multiplicand[23] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12898 = io_multiplicand[24] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12901 = io_multiplicand[25] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12904 = io_multiplicand[26] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12907 = io_multiplicand[27] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12910 = io_multiplicand[28] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12913 = io_multiplicand[29] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12916 = io_multiplicand[30] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12919 = io_multiplicand[31] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12922 = io_multiplicand[32] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12925 = io_multiplicand[33] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12928 = io_multiplicand[34] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12931 = io_multiplicand[35] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12934 = io_multiplicand[36] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12937 = io_multiplicand[37] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12940 = io_multiplicand[38] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12943 = io_multiplicand[39] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12946 = io_multiplicand[40] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12949 = io_multiplicand[41] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12952 = io_multiplicand[42] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12955 = io_multiplicand[43] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12958 = io_multiplicand[44] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12961 = io_multiplicand[45] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12964 = io_multiplicand[46] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12967 = io_multiplicand[47] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12970 = io_multiplicand[48] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12973 = io_multiplicand[49] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12976 = io_multiplicand[50] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12979 = io_multiplicand[51] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12982 = io_multiplicand[52] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12985 = io_multiplicand[53] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12988 = io_multiplicand[54] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12991 = io_multiplicand[55] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12994 = io_multiplicand[56] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_12997 = io_multiplicand[57] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_13000 = io_multiplicand[58] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_13003 = io_multiplicand[59] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_13006 = io_multiplicand[60] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_13009 = io_multiplicand[61] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_13012 = io_multiplicand[62] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire  _T_13015 = io_multiplicand[63] & io_multiplier[40]; // @[partialprod.scala 16:36]
  wire [9:0] _T_13024 = {_T_13015,_T_13012,_T_13009,_T_13006,_T_13003,_T_13000,_T_12997,_T_12994,_T_12991,_T_12988}; // @[Cat.scala 29:58]
  wire [18:0] _T_13033 = {_T_13024,_T_12985,_T_12982,_T_12979,_T_12976,_T_12973,_T_12970,_T_12967,_T_12964,_T_12961}; // @[Cat.scala 29:58]
  wire [27:0] _T_13042 = {_T_13033,_T_12958,_T_12955,_T_12952,_T_12949,_T_12946,_T_12943,_T_12940,_T_12937,_T_12934}; // @[Cat.scala 29:58]
  wire [36:0] _T_13051 = {_T_13042,_T_12931,_T_12928,_T_12925,_T_12922,_T_12919,_T_12916,_T_12913,_T_12910,_T_12907}; // @[Cat.scala 29:58]
  wire [45:0] _T_13060 = {_T_13051,_T_12904,_T_12901,_T_12898,_T_12895,_T_12892,_T_12889,_T_12886,_T_12883,_T_12880}; // @[Cat.scala 29:58]
  wire [54:0] _T_13069 = {_T_13060,_T_12877,_T_12874,_T_12871,_T_12868,_T_12865,_T_12862,_T_12859,_T_12856,_T_12853}; // @[Cat.scala 29:58]
  wire [62:0] _T_13077 = {_T_13069,_T_12850,_T_12847,_T_12844,_T_12841,_T_12838,_T_12835,_T_12832,_T_12829}; // @[Cat.scala 29:58]
  wire  _T_13145 = io_multiplicand[0] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13148 = io_multiplicand[1] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13151 = io_multiplicand[2] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13154 = io_multiplicand[3] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13157 = io_multiplicand[4] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13160 = io_multiplicand[5] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13163 = io_multiplicand[6] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13166 = io_multiplicand[7] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13169 = io_multiplicand[8] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13172 = io_multiplicand[9] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13175 = io_multiplicand[10] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13178 = io_multiplicand[11] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13181 = io_multiplicand[12] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13184 = io_multiplicand[13] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13187 = io_multiplicand[14] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13190 = io_multiplicand[15] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13193 = io_multiplicand[16] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13196 = io_multiplicand[17] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13199 = io_multiplicand[18] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13202 = io_multiplicand[19] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13205 = io_multiplicand[20] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13208 = io_multiplicand[21] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13211 = io_multiplicand[22] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13214 = io_multiplicand[23] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13217 = io_multiplicand[24] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13220 = io_multiplicand[25] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13223 = io_multiplicand[26] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13226 = io_multiplicand[27] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13229 = io_multiplicand[28] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13232 = io_multiplicand[29] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13235 = io_multiplicand[30] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13238 = io_multiplicand[31] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13241 = io_multiplicand[32] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13244 = io_multiplicand[33] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13247 = io_multiplicand[34] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13250 = io_multiplicand[35] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13253 = io_multiplicand[36] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13256 = io_multiplicand[37] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13259 = io_multiplicand[38] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13262 = io_multiplicand[39] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13265 = io_multiplicand[40] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13268 = io_multiplicand[41] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13271 = io_multiplicand[42] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13274 = io_multiplicand[43] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13277 = io_multiplicand[44] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13280 = io_multiplicand[45] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13283 = io_multiplicand[46] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13286 = io_multiplicand[47] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13289 = io_multiplicand[48] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13292 = io_multiplicand[49] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13295 = io_multiplicand[50] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13298 = io_multiplicand[51] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13301 = io_multiplicand[52] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13304 = io_multiplicand[53] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13307 = io_multiplicand[54] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13310 = io_multiplicand[55] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13313 = io_multiplicand[56] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13316 = io_multiplicand[57] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13319 = io_multiplicand[58] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13322 = io_multiplicand[59] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13325 = io_multiplicand[60] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13328 = io_multiplicand[61] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13331 = io_multiplicand[62] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire  _T_13334 = io_multiplicand[63] & io_multiplier[41]; // @[partialprod.scala 16:36]
  wire [9:0] _T_13343 = {_T_13334,_T_13331,_T_13328,_T_13325,_T_13322,_T_13319,_T_13316,_T_13313,_T_13310,_T_13307}; // @[Cat.scala 29:58]
  wire [18:0] _T_13352 = {_T_13343,_T_13304,_T_13301,_T_13298,_T_13295,_T_13292,_T_13289,_T_13286,_T_13283,_T_13280}; // @[Cat.scala 29:58]
  wire [27:0] _T_13361 = {_T_13352,_T_13277,_T_13274,_T_13271,_T_13268,_T_13265,_T_13262,_T_13259,_T_13256,_T_13253}; // @[Cat.scala 29:58]
  wire [36:0] _T_13370 = {_T_13361,_T_13250,_T_13247,_T_13244,_T_13241,_T_13238,_T_13235,_T_13232,_T_13229,_T_13226}; // @[Cat.scala 29:58]
  wire [45:0] _T_13379 = {_T_13370,_T_13223,_T_13220,_T_13217,_T_13214,_T_13211,_T_13208,_T_13205,_T_13202,_T_13199}; // @[Cat.scala 29:58]
  wire [54:0] _T_13388 = {_T_13379,_T_13196,_T_13193,_T_13190,_T_13187,_T_13184,_T_13181,_T_13178,_T_13175,_T_13172}; // @[Cat.scala 29:58]
  wire [62:0] _T_13396 = {_T_13388,_T_13169,_T_13166,_T_13163,_T_13160,_T_13157,_T_13154,_T_13151,_T_13148}; // @[Cat.scala 29:58]
  wire  _T_13464 = io_multiplicand[0] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13467 = io_multiplicand[1] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13470 = io_multiplicand[2] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13473 = io_multiplicand[3] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13476 = io_multiplicand[4] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13479 = io_multiplicand[5] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13482 = io_multiplicand[6] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13485 = io_multiplicand[7] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13488 = io_multiplicand[8] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13491 = io_multiplicand[9] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13494 = io_multiplicand[10] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13497 = io_multiplicand[11] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13500 = io_multiplicand[12] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13503 = io_multiplicand[13] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13506 = io_multiplicand[14] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13509 = io_multiplicand[15] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13512 = io_multiplicand[16] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13515 = io_multiplicand[17] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13518 = io_multiplicand[18] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13521 = io_multiplicand[19] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13524 = io_multiplicand[20] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13527 = io_multiplicand[21] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13530 = io_multiplicand[22] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13533 = io_multiplicand[23] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13536 = io_multiplicand[24] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13539 = io_multiplicand[25] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13542 = io_multiplicand[26] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13545 = io_multiplicand[27] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13548 = io_multiplicand[28] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13551 = io_multiplicand[29] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13554 = io_multiplicand[30] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13557 = io_multiplicand[31] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13560 = io_multiplicand[32] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13563 = io_multiplicand[33] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13566 = io_multiplicand[34] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13569 = io_multiplicand[35] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13572 = io_multiplicand[36] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13575 = io_multiplicand[37] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13578 = io_multiplicand[38] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13581 = io_multiplicand[39] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13584 = io_multiplicand[40] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13587 = io_multiplicand[41] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13590 = io_multiplicand[42] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13593 = io_multiplicand[43] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13596 = io_multiplicand[44] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13599 = io_multiplicand[45] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13602 = io_multiplicand[46] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13605 = io_multiplicand[47] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13608 = io_multiplicand[48] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13611 = io_multiplicand[49] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13614 = io_multiplicand[50] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13617 = io_multiplicand[51] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13620 = io_multiplicand[52] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13623 = io_multiplicand[53] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13626 = io_multiplicand[54] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13629 = io_multiplicand[55] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13632 = io_multiplicand[56] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13635 = io_multiplicand[57] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13638 = io_multiplicand[58] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13641 = io_multiplicand[59] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13644 = io_multiplicand[60] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13647 = io_multiplicand[61] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13650 = io_multiplicand[62] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire  _T_13653 = io_multiplicand[63] & io_multiplier[42]; // @[partialprod.scala 16:36]
  wire [9:0] _T_13662 = {_T_13653,_T_13650,_T_13647,_T_13644,_T_13641,_T_13638,_T_13635,_T_13632,_T_13629,_T_13626}; // @[Cat.scala 29:58]
  wire [18:0] _T_13671 = {_T_13662,_T_13623,_T_13620,_T_13617,_T_13614,_T_13611,_T_13608,_T_13605,_T_13602,_T_13599}; // @[Cat.scala 29:58]
  wire [27:0] _T_13680 = {_T_13671,_T_13596,_T_13593,_T_13590,_T_13587,_T_13584,_T_13581,_T_13578,_T_13575,_T_13572}; // @[Cat.scala 29:58]
  wire [36:0] _T_13689 = {_T_13680,_T_13569,_T_13566,_T_13563,_T_13560,_T_13557,_T_13554,_T_13551,_T_13548,_T_13545}; // @[Cat.scala 29:58]
  wire [45:0] _T_13698 = {_T_13689,_T_13542,_T_13539,_T_13536,_T_13533,_T_13530,_T_13527,_T_13524,_T_13521,_T_13518}; // @[Cat.scala 29:58]
  wire [54:0] _T_13707 = {_T_13698,_T_13515,_T_13512,_T_13509,_T_13506,_T_13503,_T_13500,_T_13497,_T_13494,_T_13491}; // @[Cat.scala 29:58]
  wire [62:0] _T_13715 = {_T_13707,_T_13488,_T_13485,_T_13482,_T_13479,_T_13476,_T_13473,_T_13470,_T_13467}; // @[Cat.scala 29:58]
  wire  _T_13783 = io_multiplicand[0] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13786 = io_multiplicand[1] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13789 = io_multiplicand[2] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13792 = io_multiplicand[3] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13795 = io_multiplicand[4] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13798 = io_multiplicand[5] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13801 = io_multiplicand[6] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13804 = io_multiplicand[7] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13807 = io_multiplicand[8] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13810 = io_multiplicand[9] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13813 = io_multiplicand[10] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13816 = io_multiplicand[11] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13819 = io_multiplicand[12] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13822 = io_multiplicand[13] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13825 = io_multiplicand[14] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13828 = io_multiplicand[15] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13831 = io_multiplicand[16] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13834 = io_multiplicand[17] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13837 = io_multiplicand[18] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13840 = io_multiplicand[19] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13843 = io_multiplicand[20] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13846 = io_multiplicand[21] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13849 = io_multiplicand[22] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13852 = io_multiplicand[23] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13855 = io_multiplicand[24] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13858 = io_multiplicand[25] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13861 = io_multiplicand[26] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13864 = io_multiplicand[27] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13867 = io_multiplicand[28] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13870 = io_multiplicand[29] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13873 = io_multiplicand[30] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13876 = io_multiplicand[31] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13879 = io_multiplicand[32] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13882 = io_multiplicand[33] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13885 = io_multiplicand[34] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13888 = io_multiplicand[35] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13891 = io_multiplicand[36] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13894 = io_multiplicand[37] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13897 = io_multiplicand[38] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13900 = io_multiplicand[39] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13903 = io_multiplicand[40] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13906 = io_multiplicand[41] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13909 = io_multiplicand[42] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13912 = io_multiplicand[43] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13915 = io_multiplicand[44] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13918 = io_multiplicand[45] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13921 = io_multiplicand[46] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13924 = io_multiplicand[47] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13927 = io_multiplicand[48] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13930 = io_multiplicand[49] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13933 = io_multiplicand[50] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13936 = io_multiplicand[51] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13939 = io_multiplicand[52] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13942 = io_multiplicand[53] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13945 = io_multiplicand[54] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13948 = io_multiplicand[55] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13951 = io_multiplicand[56] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13954 = io_multiplicand[57] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13957 = io_multiplicand[58] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13960 = io_multiplicand[59] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13963 = io_multiplicand[60] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13966 = io_multiplicand[61] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13969 = io_multiplicand[62] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire  _T_13972 = io_multiplicand[63] & io_multiplier[43]; // @[partialprod.scala 16:36]
  wire [9:0] _T_13981 = {_T_13972,_T_13969,_T_13966,_T_13963,_T_13960,_T_13957,_T_13954,_T_13951,_T_13948,_T_13945}; // @[Cat.scala 29:58]
  wire [18:0] _T_13990 = {_T_13981,_T_13942,_T_13939,_T_13936,_T_13933,_T_13930,_T_13927,_T_13924,_T_13921,_T_13918}; // @[Cat.scala 29:58]
  wire [27:0] _T_13999 = {_T_13990,_T_13915,_T_13912,_T_13909,_T_13906,_T_13903,_T_13900,_T_13897,_T_13894,_T_13891}; // @[Cat.scala 29:58]
  wire [36:0] _T_14008 = {_T_13999,_T_13888,_T_13885,_T_13882,_T_13879,_T_13876,_T_13873,_T_13870,_T_13867,_T_13864}; // @[Cat.scala 29:58]
  wire [45:0] _T_14017 = {_T_14008,_T_13861,_T_13858,_T_13855,_T_13852,_T_13849,_T_13846,_T_13843,_T_13840,_T_13837}; // @[Cat.scala 29:58]
  wire [54:0] _T_14026 = {_T_14017,_T_13834,_T_13831,_T_13828,_T_13825,_T_13822,_T_13819,_T_13816,_T_13813,_T_13810}; // @[Cat.scala 29:58]
  wire [62:0] _T_14034 = {_T_14026,_T_13807,_T_13804,_T_13801,_T_13798,_T_13795,_T_13792,_T_13789,_T_13786}; // @[Cat.scala 29:58]
  wire  _T_14102 = io_multiplicand[0] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14105 = io_multiplicand[1] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14108 = io_multiplicand[2] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14111 = io_multiplicand[3] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14114 = io_multiplicand[4] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14117 = io_multiplicand[5] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14120 = io_multiplicand[6] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14123 = io_multiplicand[7] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14126 = io_multiplicand[8] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14129 = io_multiplicand[9] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14132 = io_multiplicand[10] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14135 = io_multiplicand[11] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14138 = io_multiplicand[12] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14141 = io_multiplicand[13] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14144 = io_multiplicand[14] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14147 = io_multiplicand[15] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14150 = io_multiplicand[16] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14153 = io_multiplicand[17] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14156 = io_multiplicand[18] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14159 = io_multiplicand[19] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14162 = io_multiplicand[20] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14165 = io_multiplicand[21] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14168 = io_multiplicand[22] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14171 = io_multiplicand[23] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14174 = io_multiplicand[24] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14177 = io_multiplicand[25] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14180 = io_multiplicand[26] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14183 = io_multiplicand[27] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14186 = io_multiplicand[28] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14189 = io_multiplicand[29] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14192 = io_multiplicand[30] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14195 = io_multiplicand[31] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14198 = io_multiplicand[32] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14201 = io_multiplicand[33] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14204 = io_multiplicand[34] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14207 = io_multiplicand[35] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14210 = io_multiplicand[36] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14213 = io_multiplicand[37] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14216 = io_multiplicand[38] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14219 = io_multiplicand[39] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14222 = io_multiplicand[40] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14225 = io_multiplicand[41] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14228 = io_multiplicand[42] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14231 = io_multiplicand[43] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14234 = io_multiplicand[44] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14237 = io_multiplicand[45] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14240 = io_multiplicand[46] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14243 = io_multiplicand[47] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14246 = io_multiplicand[48] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14249 = io_multiplicand[49] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14252 = io_multiplicand[50] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14255 = io_multiplicand[51] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14258 = io_multiplicand[52] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14261 = io_multiplicand[53] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14264 = io_multiplicand[54] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14267 = io_multiplicand[55] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14270 = io_multiplicand[56] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14273 = io_multiplicand[57] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14276 = io_multiplicand[58] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14279 = io_multiplicand[59] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14282 = io_multiplicand[60] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14285 = io_multiplicand[61] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14288 = io_multiplicand[62] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire  _T_14291 = io_multiplicand[63] & io_multiplier[44]; // @[partialprod.scala 16:36]
  wire [9:0] _T_14300 = {_T_14291,_T_14288,_T_14285,_T_14282,_T_14279,_T_14276,_T_14273,_T_14270,_T_14267,_T_14264}; // @[Cat.scala 29:58]
  wire [18:0] _T_14309 = {_T_14300,_T_14261,_T_14258,_T_14255,_T_14252,_T_14249,_T_14246,_T_14243,_T_14240,_T_14237}; // @[Cat.scala 29:58]
  wire [27:0] _T_14318 = {_T_14309,_T_14234,_T_14231,_T_14228,_T_14225,_T_14222,_T_14219,_T_14216,_T_14213,_T_14210}; // @[Cat.scala 29:58]
  wire [36:0] _T_14327 = {_T_14318,_T_14207,_T_14204,_T_14201,_T_14198,_T_14195,_T_14192,_T_14189,_T_14186,_T_14183}; // @[Cat.scala 29:58]
  wire [45:0] _T_14336 = {_T_14327,_T_14180,_T_14177,_T_14174,_T_14171,_T_14168,_T_14165,_T_14162,_T_14159,_T_14156}; // @[Cat.scala 29:58]
  wire [54:0] _T_14345 = {_T_14336,_T_14153,_T_14150,_T_14147,_T_14144,_T_14141,_T_14138,_T_14135,_T_14132,_T_14129}; // @[Cat.scala 29:58]
  wire [62:0] _T_14353 = {_T_14345,_T_14126,_T_14123,_T_14120,_T_14117,_T_14114,_T_14111,_T_14108,_T_14105}; // @[Cat.scala 29:58]
  wire  _T_14421 = io_multiplicand[0] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14424 = io_multiplicand[1] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14427 = io_multiplicand[2] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14430 = io_multiplicand[3] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14433 = io_multiplicand[4] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14436 = io_multiplicand[5] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14439 = io_multiplicand[6] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14442 = io_multiplicand[7] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14445 = io_multiplicand[8] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14448 = io_multiplicand[9] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14451 = io_multiplicand[10] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14454 = io_multiplicand[11] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14457 = io_multiplicand[12] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14460 = io_multiplicand[13] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14463 = io_multiplicand[14] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14466 = io_multiplicand[15] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14469 = io_multiplicand[16] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14472 = io_multiplicand[17] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14475 = io_multiplicand[18] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14478 = io_multiplicand[19] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14481 = io_multiplicand[20] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14484 = io_multiplicand[21] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14487 = io_multiplicand[22] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14490 = io_multiplicand[23] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14493 = io_multiplicand[24] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14496 = io_multiplicand[25] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14499 = io_multiplicand[26] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14502 = io_multiplicand[27] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14505 = io_multiplicand[28] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14508 = io_multiplicand[29] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14511 = io_multiplicand[30] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14514 = io_multiplicand[31] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14517 = io_multiplicand[32] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14520 = io_multiplicand[33] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14523 = io_multiplicand[34] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14526 = io_multiplicand[35] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14529 = io_multiplicand[36] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14532 = io_multiplicand[37] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14535 = io_multiplicand[38] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14538 = io_multiplicand[39] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14541 = io_multiplicand[40] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14544 = io_multiplicand[41] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14547 = io_multiplicand[42] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14550 = io_multiplicand[43] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14553 = io_multiplicand[44] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14556 = io_multiplicand[45] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14559 = io_multiplicand[46] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14562 = io_multiplicand[47] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14565 = io_multiplicand[48] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14568 = io_multiplicand[49] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14571 = io_multiplicand[50] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14574 = io_multiplicand[51] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14577 = io_multiplicand[52] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14580 = io_multiplicand[53] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14583 = io_multiplicand[54] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14586 = io_multiplicand[55] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14589 = io_multiplicand[56] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14592 = io_multiplicand[57] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14595 = io_multiplicand[58] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14598 = io_multiplicand[59] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14601 = io_multiplicand[60] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14604 = io_multiplicand[61] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14607 = io_multiplicand[62] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire  _T_14610 = io_multiplicand[63] & io_multiplier[45]; // @[partialprod.scala 16:36]
  wire [9:0] _T_14619 = {_T_14610,_T_14607,_T_14604,_T_14601,_T_14598,_T_14595,_T_14592,_T_14589,_T_14586,_T_14583}; // @[Cat.scala 29:58]
  wire [18:0] _T_14628 = {_T_14619,_T_14580,_T_14577,_T_14574,_T_14571,_T_14568,_T_14565,_T_14562,_T_14559,_T_14556}; // @[Cat.scala 29:58]
  wire [27:0] _T_14637 = {_T_14628,_T_14553,_T_14550,_T_14547,_T_14544,_T_14541,_T_14538,_T_14535,_T_14532,_T_14529}; // @[Cat.scala 29:58]
  wire [36:0] _T_14646 = {_T_14637,_T_14526,_T_14523,_T_14520,_T_14517,_T_14514,_T_14511,_T_14508,_T_14505,_T_14502}; // @[Cat.scala 29:58]
  wire [45:0] _T_14655 = {_T_14646,_T_14499,_T_14496,_T_14493,_T_14490,_T_14487,_T_14484,_T_14481,_T_14478,_T_14475}; // @[Cat.scala 29:58]
  wire [54:0] _T_14664 = {_T_14655,_T_14472,_T_14469,_T_14466,_T_14463,_T_14460,_T_14457,_T_14454,_T_14451,_T_14448}; // @[Cat.scala 29:58]
  wire [62:0] _T_14672 = {_T_14664,_T_14445,_T_14442,_T_14439,_T_14436,_T_14433,_T_14430,_T_14427,_T_14424}; // @[Cat.scala 29:58]
  wire  _T_14740 = io_multiplicand[0] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14743 = io_multiplicand[1] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14746 = io_multiplicand[2] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14749 = io_multiplicand[3] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14752 = io_multiplicand[4] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14755 = io_multiplicand[5] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14758 = io_multiplicand[6] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14761 = io_multiplicand[7] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14764 = io_multiplicand[8] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14767 = io_multiplicand[9] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14770 = io_multiplicand[10] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14773 = io_multiplicand[11] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14776 = io_multiplicand[12] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14779 = io_multiplicand[13] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14782 = io_multiplicand[14] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14785 = io_multiplicand[15] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14788 = io_multiplicand[16] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14791 = io_multiplicand[17] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14794 = io_multiplicand[18] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14797 = io_multiplicand[19] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14800 = io_multiplicand[20] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14803 = io_multiplicand[21] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14806 = io_multiplicand[22] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14809 = io_multiplicand[23] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14812 = io_multiplicand[24] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14815 = io_multiplicand[25] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14818 = io_multiplicand[26] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14821 = io_multiplicand[27] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14824 = io_multiplicand[28] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14827 = io_multiplicand[29] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14830 = io_multiplicand[30] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14833 = io_multiplicand[31] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14836 = io_multiplicand[32] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14839 = io_multiplicand[33] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14842 = io_multiplicand[34] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14845 = io_multiplicand[35] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14848 = io_multiplicand[36] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14851 = io_multiplicand[37] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14854 = io_multiplicand[38] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14857 = io_multiplicand[39] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14860 = io_multiplicand[40] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14863 = io_multiplicand[41] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14866 = io_multiplicand[42] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14869 = io_multiplicand[43] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14872 = io_multiplicand[44] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14875 = io_multiplicand[45] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14878 = io_multiplicand[46] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14881 = io_multiplicand[47] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14884 = io_multiplicand[48] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14887 = io_multiplicand[49] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14890 = io_multiplicand[50] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14893 = io_multiplicand[51] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14896 = io_multiplicand[52] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14899 = io_multiplicand[53] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14902 = io_multiplicand[54] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14905 = io_multiplicand[55] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14908 = io_multiplicand[56] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14911 = io_multiplicand[57] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14914 = io_multiplicand[58] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14917 = io_multiplicand[59] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14920 = io_multiplicand[60] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14923 = io_multiplicand[61] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14926 = io_multiplicand[62] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire  _T_14929 = io_multiplicand[63] & io_multiplier[46]; // @[partialprod.scala 16:36]
  wire [9:0] _T_14938 = {_T_14929,_T_14926,_T_14923,_T_14920,_T_14917,_T_14914,_T_14911,_T_14908,_T_14905,_T_14902}; // @[Cat.scala 29:58]
  wire [18:0] _T_14947 = {_T_14938,_T_14899,_T_14896,_T_14893,_T_14890,_T_14887,_T_14884,_T_14881,_T_14878,_T_14875}; // @[Cat.scala 29:58]
  wire [27:0] _T_14956 = {_T_14947,_T_14872,_T_14869,_T_14866,_T_14863,_T_14860,_T_14857,_T_14854,_T_14851,_T_14848}; // @[Cat.scala 29:58]
  wire [36:0] _T_14965 = {_T_14956,_T_14845,_T_14842,_T_14839,_T_14836,_T_14833,_T_14830,_T_14827,_T_14824,_T_14821}; // @[Cat.scala 29:58]
  wire [45:0] _T_14974 = {_T_14965,_T_14818,_T_14815,_T_14812,_T_14809,_T_14806,_T_14803,_T_14800,_T_14797,_T_14794}; // @[Cat.scala 29:58]
  wire [54:0] _T_14983 = {_T_14974,_T_14791,_T_14788,_T_14785,_T_14782,_T_14779,_T_14776,_T_14773,_T_14770,_T_14767}; // @[Cat.scala 29:58]
  wire [62:0] _T_14991 = {_T_14983,_T_14764,_T_14761,_T_14758,_T_14755,_T_14752,_T_14749,_T_14746,_T_14743}; // @[Cat.scala 29:58]
  wire  _T_15059 = io_multiplicand[0] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15062 = io_multiplicand[1] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15065 = io_multiplicand[2] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15068 = io_multiplicand[3] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15071 = io_multiplicand[4] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15074 = io_multiplicand[5] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15077 = io_multiplicand[6] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15080 = io_multiplicand[7] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15083 = io_multiplicand[8] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15086 = io_multiplicand[9] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15089 = io_multiplicand[10] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15092 = io_multiplicand[11] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15095 = io_multiplicand[12] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15098 = io_multiplicand[13] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15101 = io_multiplicand[14] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15104 = io_multiplicand[15] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15107 = io_multiplicand[16] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15110 = io_multiplicand[17] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15113 = io_multiplicand[18] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15116 = io_multiplicand[19] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15119 = io_multiplicand[20] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15122 = io_multiplicand[21] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15125 = io_multiplicand[22] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15128 = io_multiplicand[23] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15131 = io_multiplicand[24] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15134 = io_multiplicand[25] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15137 = io_multiplicand[26] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15140 = io_multiplicand[27] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15143 = io_multiplicand[28] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15146 = io_multiplicand[29] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15149 = io_multiplicand[30] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15152 = io_multiplicand[31] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15155 = io_multiplicand[32] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15158 = io_multiplicand[33] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15161 = io_multiplicand[34] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15164 = io_multiplicand[35] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15167 = io_multiplicand[36] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15170 = io_multiplicand[37] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15173 = io_multiplicand[38] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15176 = io_multiplicand[39] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15179 = io_multiplicand[40] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15182 = io_multiplicand[41] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15185 = io_multiplicand[42] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15188 = io_multiplicand[43] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15191 = io_multiplicand[44] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15194 = io_multiplicand[45] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15197 = io_multiplicand[46] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15200 = io_multiplicand[47] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15203 = io_multiplicand[48] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15206 = io_multiplicand[49] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15209 = io_multiplicand[50] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15212 = io_multiplicand[51] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15215 = io_multiplicand[52] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15218 = io_multiplicand[53] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15221 = io_multiplicand[54] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15224 = io_multiplicand[55] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15227 = io_multiplicand[56] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15230 = io_multiplicand[57] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15233 = io_multiplicand[58] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15236 = io_multiplicand[59] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15239 = io_multiplicand[60] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15242 = io_multiplicand[61] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15245 = io_multiplicand[62] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire  _T_15248 = io_multiplicand[63] & io_multiplier[47]; // @[partialprod.scala 16:36]
  wire [9:0] _T_15257 = {_T_15248,_T_15245,_T_15242,_T_15239,_T_15236,_T_15233,_T_15230,_T_15227,_T_15224,_T_15221}; // @[Cat.scala 29:58]
  wire [18:0] _T_15266 = {_T_15257,_T_15218,_T_15215,_T_15212,_T_15209,_T_15206,_T_15203,_T_15200,_T_15197,_T_15194}; // @[Cat.scala 29:58]
  wire [27:0] _T_15275 = {_T_15266,_T_15191,_T_15188,_T_15185,_T_15182,_T_15179,_T_15176,_T_15173,_T_15170,_T_15167}; // @[Cat.scala 29:58]
  wire [36:0] _T_15284 = {_T_15275,_T_15164,_T_15161,_T_15158,_T_15155,_T_15152,_T_15149,_T_15146,_T_15143,_T_15140}; // @[Cat.scala 29:58]
  wire [45:0] _T_15293 = {_T_15284,_T_15137,_T_15134,_T_15131,_T_15128,_T_15125,_T_15122,_T_15119,_T_15116,_T_15113}; // @[Cat.scala 29:58]
  wire [54:0] _T_15302 = {_T_15293,_T_15110,_T_15107,_T_15104,_T_15101,_T_15098,_T_15095,_T_15092,_T_15089,_T_15086}; // @[Cat.scala 29:58]
  wire [62:0] _T_15310 = {_T_15302,_T_15083,_T_15080,_T_15077,_T_15074,_T_15071,_T_15068,_T_15065,_T_15062}; // @[Cat.scala 29:58]
  wire  _T_15378 = io_multiplicand[0] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15381 = io_multiplicand[1] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15384 = io_multiplicand[2] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15387 = io_multiplicand[3] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15390 = io_multiplicand[4] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15393 = io_multiplicand[5] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15396 = io_multiplicand[6] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15399 = io_multiplicand[7] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15402 = io_multiplicand[8] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15405 = io_multiplicand[9] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15408 = io_multiplicand[10] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15411 = io_multiplicand[11] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15414 = io_multiplicand[12] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15417 = io_multiplicand[13] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15420 = io_multiplicand[14] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15423 = io_multiplicand[15] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15426 = io_multiplicand[16] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15429 = io_multiplicand[17] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15432 = io_multiplicand[18] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15435 = io_multiplicand[19] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15438 = io_multiplicand[20] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15441 = io_multiplicand[21] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15444 = io_multiplicand[22] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15447 = io_multiplicand[23] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15450 = io_multiplicand[24] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15453 = io_multiplicand[25] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15456 = io_multiplicand[26] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15459 = io_multiplicand[27] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15462 = io_multiplicand[28] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15465 = io_multiplicand[29] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15468 = io_multiplicand[30] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15471 = io_multiplicand[31] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15474 = io_multiplicand[32] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15477 = io_multiplicand[33] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15480 = io_multiplicand[34] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15483 = io_multiplicand[35] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15486 = io_multiplicand[36] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15489 = io_multiplicand[37] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15492 = io_multiplicand[38] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15495 = io_multiplicand[39] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15498 = io_multiplicand[40] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15501 = io_multiplicand[41] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15504 = io_multiplicand[42] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15507 = io_multiplicand[43] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15510 = io_multiplicand[44] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15513 = io_multiplicand[45] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15516 = io_multiplicand[46] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15519 = io_multiplicand[47] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15522 = io_multiplicand[48] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15525 = io_multiplicand[49] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15528 = io_multiplicand[50] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15531 = io_multiplicand[51] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15534 = io_multiplicand[52] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15537 = io_multiplicand[53] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15540 = io_multiplicand[54] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15543 = io_multiplicand[55] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15546 = io_multiplicand[56] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15549 = io_multiplicand[57] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15552 = io_multiplicand[58] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15555 = io_multiplicand[59] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15558 = io_multiplicand[60] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15561 = io_multiplicand[61] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15564 = io_multiplicand[62] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire  _T_15567 = io_multiplicand[63] & io_multiplier[48]; // @[partialprod.scala 16:36]
  wire [9:0] _T_15576 = {_T_15567,_T_15564,_T_15561,_T_15558,_T_15555,_T_15552,_T_15549,_T_15546,_T_15543,_T_15540}; // @[Cat.scala 29:58]
  wire [18:0] _T_15585 = {_T_15576,_T_15537,_T_15534,_T_15531,_T_15528,_T_15525,_T_15522,_T_15519,_T_15516,_T_15513}; // @[Cat.scala 29:58]
  wire [27:0] _T_15594 = {_T_15585,_T_15510,_T_15507,_T_15504,_T_15501,_T_15498,_T_15495,_T_15492,_T_15489,_T_15486}; // @[Cat.scala 29:58]
  wire [36:0] _T_15603 = {_T_15594,_T_15483,_T_15480,_T_15477,_T_15474,_T_15471,_T_15468,_T_15465,_T_15462,_T_15459}; // @[Cat.scala 29:58]
  wire [45:0] _T_15612 = {_T_15603,_T_15456,_T_15453,_T_15450,_T_15447,_T_15444,_T_15441,_T_15438,_T_15435,_T_15432}; // @[Cat.scala 29:58]
  wire [54:0] _T_15621 = {_T_15612,_T_15429,_T_15426,_T_15423,_T_15420,_T_15417,_T_15414,_T_15411,_T_15408,_T_15405}; // @[Cat.scala 29:58]
  wire [62:0] _T_15629 = {_T_15621,_T_15402,_T_15399,_T_15396,_T_15393,_T_15390,_T_15387,_T_15384,_T_15381}; // @[Cat.scala 29:58]
  wire  _T_15697 = io_multiplicand[0] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15700 = io_multiplicand[1] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15703 = io_multiplicand[2] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15706 = io_multiplicand[3] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15709 = io_multiplicand[4] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15712 = io_multiplicand[5] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15715 = io_multiplicand[6] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15718 = io_multiplicand[7] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15721 = io_multiplicand[8] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15724 = io_multiplicand[9] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15727 = io_multiplicand[10] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15730 = io_multiplicand[11] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15733 = io_multiplicand[12] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15736 = io_multiplicand[13] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15739 = io_multiplicand[14] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15742 = io_multiplicand[15] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15745 = io_multiplicand[16] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15748 = io_multiplicand[17] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15751 = io_multiplicand[18] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15754 = io_multiplicand[19] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15757 = io_multiplicand[20] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15760 = io_multiplicand[21] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15763 = io_multiplicand[22] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15766 = io_multiplicand[23] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15769 = io_multiplicand[24] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15772 = io_multiplicand[25] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15775 = io_multiplicand[26] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15778 = io_multiplicand[27] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15781 = io_multiplicand[28] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15784 = io_multiplicand[29] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15787 = io_multiplicand[30] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15790 = io_multiplicand[31] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15793 = io_multiplicand[32] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15796 = io_multiplicand[33] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15799 = io_multiplicand[34] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15802 = io_multiplicand[35] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15805 = io_multiplicand[36] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15808 = io_multiplicand[37] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15811 = io_multiplicand[38] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15814 = io_multiplicand[39] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15817 = io_multiplicand[40] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15820 = io_multiplicand[41] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15823 = io_multiplicand[42] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15826 = io_multiplicand[43] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15829 = io_multiplicand[44] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15832 = io_multiplicand[45] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15835 = io_multiplicand[46] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15838 = io_multiplicand[47] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15841 = io_multiplicand[48] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15844 = io_multiplicand[49] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15847 = io_multiplicand[50] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15850 = io_multiplicand[51] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15853 = io_multiplicand[52] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15856 = io_multiplicand[53] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15859 = io_multiplicand[54] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15862 = io_multiplicand[55] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15865 = io_multiplicand[56] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15868 = io_multiplicand[57] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15871 = io_multiplicand[58] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15874 = io_multiplicand[59] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15877 = io_multiplicand[60] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15880 = io_multiplicand[61] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15883 = io_multiplicand[62] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire  _T_15886 = io_multiplicand[63] & io_multiplier[49]; // @[partialprod.scala 16:36]
  wire [9:0] _T_15895 = {_T_15886,_T_15883,_T_15880,_T_15877,_T_15874,_T_15871,_T_15868,_T_15865,_T_15862,_T_15859}; // @[Cat.scala 29:58]
  wire [18:0] _T_15904 = {_T_15895,_T_15856,_T_15853,_T_15850,_T_15847,_T_15844,_T_15841,_T_15838,_T_15835,_T_15832}; // @[Cat.scala 29:58]
  wire [27:0] _T_15913 = {_T_15904,_T_15829,_T_15826,_T_15823,_T_15820,_T_15817,_T_15814,_T_15811,_T_15808,_T_15805}; // @[Cat.scala 29:58]
  wire [36:0] _T_15922 = {_T_15913,_T_15802,_T_15799,_T_15796,_T_15793,_T_15790,_T_15787,_T_15784,_T_15781,_T_15778}; // @[Cat.scala 29:58]
  wire [45:0] _T_15931 = {_T_15922,_T_15775,_T_15772,_T_15769,_T_15766,_T_15763,_T_15760,_T_15757,_T_15754,_T_15751}; // @[Cat.scala 29:58]
  wire [54:0] _T_15940 = {_T_15931,_T_15748,_T_15745,_T_15742,_T_15739,_T_15736,_T_15733,_T_15730,_T_15727,_T_15724}; // @[Cat.scala 29:58]
  wire [62:0] _T_15948 = {_T_15940,_T_15721,_T_15718,_T_15715,_T_15712,_T_15709,_T_15706,_T_15703,_T_15700}; // @[Cat.scala 29:58]
  wire  _T_16016 = io_multiplicand[0] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16019 = io_multiplicand[1] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16022 = io_multiplicand[2] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16025 = io_multiplicand[3] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16028 = io_multiplicand[4] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16031 = io_multiplicand[5] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16034 = io_multiplicand[6] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16037 = io_multiplicand[7] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16040 = io_multiplicand[8] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16043 = io_multiplicand[9] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16046 = io_multiplicand[10] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16049 = io_multiplicand[11] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16052 = io_multiplicand[12] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16055 = io_multiplicand[13] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16058 = io_multiplicand[14] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16061 = io_multiplicand[15] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16064 = io_multiplicand[16] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16067 = io_multiplicand[17] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16070 = io_multiplicand[18] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16073 = io_multiplicand[19] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16076 = io_multiplicand[20] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16079 = io_multiplicand[21] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16082 = io_multiplicand[22] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16085 = io_multiplicand[23] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16088 = io_multiplicand[24] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16091 = io_multiplicand[25] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16094 = io_multiplicand[26] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16097 = io_multiplicand[27] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16100 = io_multiplicand[28] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16103 = io_multiplicand[29] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16106 = io_multiplicand[30] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16109 = io_multiplicand[31] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16112 = io_multiplicand[32] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16115 = io_multiplicand[33] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16118 = io_multiplicand[34] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16121 = io_multiplicand[35] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16124 = io_multiplicand[36] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16127 = io_multiplicand[37] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16130 = io_multiplicand[38] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16133 = io_multiplicand[39] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16136 = io_multiplicand[40] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16139 = io_multiplicand[41] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16142 = io_multiplicand[42] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16145 = io_multiplicand[43] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16148 = io_multiplicand[44] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16151 = io_multiplicand[45] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16154 = io_multiplicand[46] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16157 = io_multiplicand[47] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16160 = io_multiplicand[48] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16163 = io_multiplicand[49] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16166 = io_multiplicand[50] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16169 = io_multiplicand[51] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16172 = io_multiplicand[52] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16175 = io_multiplicand[53] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16178 = io_multiplicand[54] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16181 = io_multiplicand[55] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16184 = io_multiplicand[56] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16187 = io_multiplicand[57] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16190 = io_multiplicand[58] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16193 = io_multiplicand[59] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16196 = io_multiplicand[60] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16199 = io_multiplicand[61] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16202 = io_multiplicand[62] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire  _T_16205 = io_multiplicand[63] & io_multiplier[50]; // @[partialprod.scala 16:36]
  wire [9:0] _T_16214 = {_T_16205,_T_16202,_T_16199,_T_16196,_T_16193,_T_16190,_T_16187,_T_16184,_T_16181,_T_16178}; // @[Cat.scala 29:58]
  wire [18:0] _T_16223 = {_T_16214,_T_16175,_T_16172,_T_16169,_T_16166,_T_16163,_T_16160,_T_16157,_T_16154,_T_16151}; // @[Cat.scala 29:58]
  wire [27:0] _T_16232 = {_T_16223,_T_16148,_T_16145,_T_16142,_T_16139,_T_16136,_T_16133,_T_16130,_T_16127,_T_16124}; // @[Cat.scala 29:58]
  wire [36:0] _T_16241 = {_T_16232,_T_16121,_T_16118,_T_16115,_T_16112,_T_16109,_T_16106,_T_16103,_T_16100,_T_16097}; // @[Cat.scala 29:58]
  wire [45:0] _T_16250 = {_T_16241,_T_16094,_T_16091,_T_16088,_T_16085,_T_16082,_T_16079,_T_16076,_T_16073,_T_16070}; // @[Cat.scala 29:58]
  wire [54:0] _T_16259 = {_T_16250,_T_16067,_T_16064,_T_16061,_T_16058,_T_16055,_T_16052,_T_16049,_T_16046,_T_16043}; // @[Cat.scala 29:58]
  wire [62:0] _T_16267 = {_T_16259,_T_16040,_T_16037,_T_16034,_T_16031,_T_16028,_T_16025,_T_16022,_T_16019}; // @[Cat.scala 29:58]
  wire  _T_16335 = io_multiplicand[0] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16338 = io_multiplicand[1] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16341 = io_multiplicand[2] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16344 = io_multiplicand[3] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16347 = io_multiplicand[4] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16350 = io_multiplicand[5] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16353 = io_multiplicand[6] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16356 = io_multiplicand[7] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16359 = io_multiplicand[8] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16362 = io_multiplicand[9] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16365 = io_multiplicand[10] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16368 = io_multiplicand[11] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16371 = io_multiplicand[12] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16374 = io_multiplicand[13] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16377 = io_multiplicand[14] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16380 = io_multiplicand[15] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16383 = io_multiplicand[16] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16386 = io_multiplicand[17] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16389 = io_multiplicand[18] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16392 = io_multiplicand[19] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16395 = io_multiplicand[20] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16398 = io_multiplicand[21] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16401 = io_multiplicand[22] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16404 = io_multiplicand[23] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16407 = io_multiplicand[24] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16410 = io_multiplicand[25] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16413 = io_multiplicand[26] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16416 = io_multiplicand[27] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16419 = io_multiplicand[28] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16422 = io_multiplicand[29] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16425 = io_multiplicand[30] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16428 = io_multiplicand[31] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16431 = io_multiplicand[32] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16434 = io_multiplicand[33] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16437 = io_multiplicand[34] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16440 = io_multiplicand[35] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16443 = io_multiplicand[36] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16446 = io_multiplicand[37] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16449 = io_multiplicand[38] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16452 = io_multiplicand[39] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16455 = io_multiplicand[40] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16458 = io_multiplicand[41] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16461 = io_multiplicand[42] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16464 = io_multiplicand[43] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16467 = io_multiplicand[44] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16470 = io_multiplicand[45] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16473 = io_multiplicand[46] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16476 = io_multiplicand[47] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16479 = io_multiplicand[48] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16482 = io_multiplicand[49] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16485 = io_multiplicand[50] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16488 = io_multiplicand[51] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16491 = io_multiplicand[52] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16494 = io_multiplicand[53] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16497 = io_multiplicand[54] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16500 = io_multiplicand[55] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16503 = io_multiplicand[56] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16506 = io_multiplicand[57] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16509 = io_multiplicand[58] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16512 = io_multiplicand[59] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16515 = io_multiplicand[60] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16518 = io_multiplicand[61] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16521 = io_multiplicand[62] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire  _T_16524 = io_multiplicand[63] & io_multiplier[51]; // @[partialprod.scala 16:36]
  wire [9:0] _T_16533 = {_T_16524,_T_16521,_T_16518,_T_16515,_T_16512,_T_16509,_T_16506,_T_16503,_T_16500,_T_16497}; // @[Cat.scala 29:58]
  wire [18:0] _T_16542 = {_T_16533,_T_16494,_T_16491,_T_16488,_T_16485,_T_16482,_T_16479,_T_16476,_T_16473,_T_16470}; // @[Cat.scala 29:58]
  wire [27:0] _T_16551 = {_T_16542,_T_16467,_T_16464,_T_16461,_T_16458,_T_16455,_T_16452,_T_16449,_T_16446,_T_16443}; // @[Cat.scala 29:58]
  wire [36:0] _T_16560 = {_T_16551,_T_16440,_T_16437,_T_16434,_T_16431,_T_16428,_T_16425,_T_16422,_T_16419,_T_16416}; // @[Cat.scala 29:58]
  wire [45:0] _T_16569 = {_T_16560,_T_16413,_T_16410,_T_16407,_T_16404,_T_16401,_T_16398,_T_16395,_T_16392,_T_16389}; // @[Cat.scala 29:58]
  wire [54:0] _T_16578 = {_T_16569,_T_16386,_T_16383,_T_16380,_T_16377,_T_16374,_T_16371,_T_16368,_T_16365,_T_16362}; // @[Cat.scala 29:58]
  wire [62:0] _T_16586 = {_T_16578,_T_16359,_T_16356,_T_16353,_T_16350,_T_16347,_T_16344,_T_16341,_T_16338}; // @[Cat.scala 29:58]
  wire  _T_16654 = io_multiplicand[0] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16657 = io_multiplicand[1] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16660 = io_multiplicand[2] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16663 = io_multiplicand[3] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16666 = io_multiplicand[4] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16669 = io_multiplicand[5] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16672 = io_multiplicand[6] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16675 = io_multiplicand[7] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16678 = io_multiplicand[8] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16681 = io_multiplicand[9] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16684 = io_multiplicand[10] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16687 = io_multiplicand[11] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16690 = io_multiplicand[12] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16693 = io_multiplicand[13] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16696 = io_multiplicand[14] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16699 = io_multiplicand[15] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16702 = io_multiplicand[16] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16705 = io_multiplicand[17] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16708 = io_multiplicand[18] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16711 = io_multiplicand[19] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16714 = io_multiplicand[20] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16717 = io_multiplicand[21] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16720 = io_multiplicand[22] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16723 = io_multiplicand[23] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16726 = io_multiplicand[24] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16729 = io_multiplicand[25] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16732 = io_multiplicand[26] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16735 = io_multiplicand[27] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16738 = io_multiplicand[28] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16741 = io_multiplicand[29] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16744 = io_multiplicand[30] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16747 = io_multiplicand[31] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16750 = io_multiplicand[32] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16753 = io_multiplicand[33] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16756 = io_multiplicand[34] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16759 = io_multiplicand[35] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16762 = io_multiplicand[36] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16765 = io_multiplicand[37] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16768 = io_multiplicand[38] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16771 = io_multiplicand[39] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16774 = io_multiplicand[40] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16777 = io_multiplicand[41] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16780 = io_multiplicand[42] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16783 = io_multiplicand[43] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16786 = io_multiplicand[44] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16789 = io_multiplicand[45] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16792 = io_multiplicand[46] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16795 = io_multiplicand[47] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16798 = io_multiplicand[48] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16801 = io_multiplicand[49] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16804 = io_multiplicand[50] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16807 = io_multiplicand[51] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16810 = io_multiplicand[52] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16813 = io_multiplicand[53] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16816 = io_multiplicand[54] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16819 = io_multiplicand[55] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16822 = io_multiplicand[56] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16825 = io_multiplicand[57] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16828 = io_multiplicand[58] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16831 = io_multiplicand[59] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16834 = io_multiplicand[60] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16837 = io_multiplicand[61] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16840 = io_multiplicand[62] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire  _T_16843 = io_multiplicand[63] & io_multiplier[52]; // @[partialprod.scala 16:36]
  wire [9:0] _T_16852 = {_T_16843,_T_16840,_T_16837,_T_16834,_T_16831,_T_16828,_T_16825,_T_16822,_T_16819,_T_16816}; // @[Cat.scala 29:58]
  wire [18:0] _T_16861 = {_T_16852,_T_16813,_T_16810,_T_16807,_T_16804,_T_16801,_T_16798,_T_16795,_T_16792,_T_16789}; // @[Cat.scala 29:58]
  wire [27:0] _T_16870 = {_T_16861,_T_16786,_T_16783,_T_16780,_T_16777,_T_16774,_T_16771,_T_16768,_T_16765,_T_16762}; // @[Cat.scala 29:58]
  wire [36:0] _T_16879 = {_T_16870,_T_16759,_T_16756,_T_16753,_T_16750,_T_16747,_T_16744,_T_16741,_T_16738,_T_16735}; // @[Cat.scala 29:58]
  wire [45:0] _T_16888 = {_T_16879,_T_16732,_T_16729,_T_16726,_T_16723,_T_16720,_T_16717,_T_16714,_T_16711,_T_16708}; // @[Cat.scala 29:58]
  wire [54:0] _T_16897 = {_T_16888,_T_16705,_T_16702,_T_16699,_T_16696,_T_16693,_T_16690,_T_16687,_T_16684,_T_16681}; // @[Cat.scala 29:58]
  wire [62:0] _T_16905 = {_T_16897,_T_16678,_T_16675,_T_16672,_T_16669,_T_16666,_T_16663,_T_16660,_T_16657}; // @[Cat.scala 29:58]
  wire  _T_16973 = io_multiplicand[0] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_16976 = io_multiplicand[1] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_16979 = io_multiplicand[2] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_16982 = io_multiplicand[3] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_16985 = io_multiplicand[4] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_16988 = io_multiplicand[5] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_16991 = io_multiplicand[6] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_16994 = io_multiplicand[7] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_16997 = io_multiplicand[8] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17000 = io_multiplicand[9] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17003 = io_multiplicand[10] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17006 = io_multiplicand[11] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17009 = io_multiplicand[12] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17012 = io_multiplicand[13] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17015 = io_multiplicand[14] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17018 = io_multiplicand[15] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17021 = io_multiplicand[16] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17024 = io_multiplicand[17] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17027 = io_multiplicand[18] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17030 = io_multiplicand[19] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17033 = io_multiplicand[20] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17036 = io_multiplicand[21] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17039 = io_multiplicand[22] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17042 = io_multiplicand[23] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17045 = io_multiplicand[24] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17048 = io_multiplicand[25] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17051 = io_multiplicand[26] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17054 = io_multiplicand[27] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17057 = io_multiplicand[28] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17060 = io_multiplicand[29] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17063 = io_multiplicand[30] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17066 = io_multiplicand[31] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17069 = io_multiplicand[32] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17072 = io_multiplicand[33] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17075 = io_multiplicand[34] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17078 = io_multiplicand[35] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17081 = io_multiplicand[36] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17084 = io_multiplicand[37] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17087 = io_multiplicand[38] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17090 = io_multiplicand[39] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17093 = io_multiplicand[40] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17096 = io_multiplicand[41] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17099 = io_multiplicand[42] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17102 = io_multiplicand[43] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17105 = io_multiplicand[44] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17108 = io_multiplicand[45] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17111 = io_multiplicand[46] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17114 = io_multiplicand[47] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17117 = io_multiplicand[48] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17120 = io_multiplicand[49] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17123 = io_multiplicand[50] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17126 = io_multiplicand[51] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17129 = io_multiplicand[52] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17132 = io_multiplicand[53] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17135 = io_multiplicand[54] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17138 = io_multiplicand[55] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17141 = io_multiplicand[56] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17144 = io_multiplicand[57] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17147 = io_multiplicand[58] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17150 = io_multiplicand[59] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17153 = io_multiplicand[60] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17156 = io_multiplicand[61] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17159 = io_multiplicand[62] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire  _T_17162 = io_multiplicand[63] & io_multiplier[53]; // @[partialprod.scala 16:36]
  wire [9:0] _T_17171 = {_T_17162,_T_17159,_T_17156,_T_17153,_T_17150,_T_17147,_T_17144,_T_17141,_T_17138,_T_17135}; // @[Cat.scala 29:58]
  wire [18:0] _T_17180 = {_T_17171,_T_17132,_T_17129,_T_17126,_T_17123,_T_17120,_T_17117,_T_17114,_T_17111,_T_17108}; // @[Cat.scala 29:58]
  wire [27:0] _T_17189 = {_T_17180,_T_17105,_T_17102,_T_17099,_T_17096,_T_17093,_T_17090,_T_17087,_T_17084,_T_17081}; // @[Cat.scala 29:58]
  wire [36:0] _T_17198 = {_T_17189,_T_17078,_T_17075,_T_17072,_T_17069,_T_17066,_T_17063,_T_17060,_T_17057,_T_17054}; // @[Cat.scala 29:58]
  wire [45:0] _T_17207 = {_T_17198,_T_17051,_T_17048,_T_17045,_T_17042,_T_17039,_T_17036,_T_17033,_T_17030,_T_17027}; // @[Cat.scala 29:58]
  wire [54:0] _T_17216 = {_T_17207,_T_17024,_T_17021,_T_17018,_T_17015,_T_17012,_T_17009,_T_17006,_T_17003,_T_17000}; // @[Cat.scala 29:58]
  wire [62:0] _T_17224 = {_T_17216,_T_16997,_T_16994,_T_16991,_T_16988,_T_16985,_T_16982,_T_16979,_T_16976}; // @[Cat.scala 29:58]
  wire  _T_17292 = io_multiplicand[0] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17295 = io_multiplicand[1] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17298 = io_multiplicand[2] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17301 = io_multiplicand[3] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17304 = io_multiplicand[4] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17307 = io_multiplicand[5] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17310 = io_multiplicand[6] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17313 = io_multiplicand[7] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17316 = io_multiplicand[8] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17319 = io_multiplicand[9] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17322 = io_multiplicand[10] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17325 = io_multiplicand[11] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17328 = io_multiplicand[12] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17331 = io_multiplicand[13] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17334 = io_multiplicand[14] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17337 = io_multiplicand[15] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17340 = io_multiplicand[16] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17343 = io_multiplicand[17] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17346 = io_multiplicand[18] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17349 = io_multiplicand[19] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17352 = io_multiplicand[20] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17355 = io_multiplicand[21] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17358 = io_multiplicand[22] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17361 = io_multiplicand[23] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17364 = io_multiplicand[24] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17367 = io_multiplicand[25] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17370 = io_multiplicand[26] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17373 = io_multiplicand[27] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17376 = io_multiplicand[28] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17379 = io_multiplicand[29] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17382 = io_multiplicand[30] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17385 = io_multiplicand[31] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17388 = io_multiplicand[32] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17391 = io_multiplicand[33] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17394 = io_multiplicand[34] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17397 = io_multiplicand[35] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17400 = io_multiplicand[36] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17403 = io_multiplicand[37] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17406 = io_multiplicand[38] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17409 = io_multiplicand[39] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17412 = io_multiplicand[40] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17415 = io_multiplicand[41] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17418 = io_multiplicand[42] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17421 = io_multiplicand[43] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17424 = io_multiplicand[44] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17427 = io_multiplicand[45] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17430 = io_multiplicand[46] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17433 = io_multiplicand[47] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17436 = io_multiplicand[48] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17439 = io_multiplicand[49] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17442 = io_multiplicand[50] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17445 = io_multiplicand[51] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17448 = io_multiplicand[52] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17451 = io_multiplicand[53] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17454 = io_multiplicand[54] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17457 = io_multiplicand[55] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17460 = io_multiplicand[56] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17463 = io_multiplicand[57] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17466 = io_multiplicand[58] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17469 = io_multiplicand[59] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17472 = io_multiplicand[60] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17475 = io_multiplicand[61] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17478 = io_multiplicand[62] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire  _T_17481 = io_multiplicand[63] & io_multiplier[54]; // @[partialprod.scala 16:36]
  wire [9:0] _T_17490 = {_T_17481,_T_17478,_T_17475,_T_17472,_T_17469,_T_17466,_T_17463,_T_17460,_T_17457,_T_17454}; // @[Cat.scala 29:58]
  wire [18:0] _T_17499 = {_T_17490,_T_17451,_T_17448,_T_17445,_T_17442,_T_17439,_T_17436,_T_17433,_T_17430,_T_17427}; // @[Cat.scala 29:58]
  wire [27:0] _T_17508 = {_T_17499,_T_17424,_T_17421,_T_17418,_T_17415,_T_17412,_T_17409,_T_17406,_T_17403,_T_17400}; // @[Cat.scala 29:58]
  wire [36:0] _T_17517 = {_T_17508,_T_17397,_T_17394,_T_17391,_T_17388,_T_17385,_T_17382,_T_17379,_T_17376,_T_17373}; // @[Cat.scala 29:58]
  wire [45:0] _T_17526 = {_T_17517,_T_17370,_T_17367,_T_17364,_T_17361,_T_17358,_T_17355,_T_17352,_T_17349,_T_17346}; // @[Cat.scala 29:58]
  wire [54:0] _T_17535 = {_T_17526,_T_17343,_T_17340,_T_17337,_T_17334,_T_17331,_T_17328,_T_17325,_T_17322,_T_17319}; // @[Cat.scala 29:58]
  wire [62:0] _T_17543 = {_T_17535,_T_17316,_T_17313,_T_17310,_T_17307,_T_17304,_T_17301,_T_17298,_T_17295}; // @[Cat.scala 29:58]
  wire  _T_17611 = io_multiplicand[0] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17614 = io_multiplicand[1] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17617 = io_multiplicand[2] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17620 = io_multiplicand[3] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17623 = io_multiplicand[4] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17626 = io_multiplicand[5] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17629 = io_multiplicand[6] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17632 = io_multiplicand[7] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17635 = io_multiplicand[8] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17638 = io_multiplicand[9] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17641 = io_multiplicand[10] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17644 = io_multiplicand[11] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17647 = io_multiplicand[12] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17650 = io_multiplicand[13] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17653 = io_multiplicand[14] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17656 = io_multiplicand[15] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17659 = io_multiplicand[16] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17662 = io_multiplicand[17] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17665 = io_multiplicand[18] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17668 = io_multiplicand[19] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17671 = io_multiplicand[20] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17674 = io_multiplicand[21] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17677 = io_multiplicand[22] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17680 = io_multiplicand[23] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17683 = io_multiplicand[24] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17686 = io_multiplicand[25] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17689 = io_multiplicand[26] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17692 = io_multiplicand[27] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17695 = io_multiplicand[28] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17698 = io_multiplicand[29] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17701 = io_multiplicand[30] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17704 = io_multiplicand[31] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17707 = io_multiplicand[32] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17710 = io_multiplicand[33] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17713 = io_multiplicand[34] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17716 = io_multiplicand[35] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17719 = io_multiplicand[36] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17722 = io_multiplicand[37] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17725 = io_multiplicand[38] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17728 = io_multiplicand[39] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17731 = io_multiplicand[40] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17734 = io_multiplicand[41] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17737 = io_multiplicand[42] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17740 = io_multiplicand[43] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17743 = io_multiplicand[44] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17746 = io_multiplicand[45] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17749 = io_multiplicand[46] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17752 = io_multiplicand[47] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17755 = io_multiplicand[48] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17758 = io_multiplicand[49] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17761 = io_multiplicand[50] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17764 = io_multiplicand[51] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17767 = io_multiplicand[52] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17770 = io_multiplicand[53] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17773 = io_multiplicand[54] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17776 = io_multiplicand[55] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17779 = io_multiplicand[56] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17782 = io_multiplicand[57] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17785 = io_multiplicand[58] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17788 = io_multiplicand[59] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17791 = io_multiplicand[60] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17794 = io_multiplicand[61] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17797 = io_multiplicand[62] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire  _T_17800 = io_multiplicand[63] & io_multiplier[55]; // @[partialprod.scala 16:36]
  wire [9:0] _T_17809 = {_T_17800,_T_17797,_T_17794,_T_17791,_T_17788,_T_17785,_T_17782,_T_17779,_T_17776,_T_17773}; // @[Cat.scala 29:58]
  wire [18:0] _T_17818 = {_T_17809,_T_17770,_T_17767,_T_17764,_T_17761,_T_17758,_T_17755,_T_17752,_T_17749,_T_17746}; // @[Cat.scala 29:58]
  wire [27:0] _T_17827 = {_T_17818,_T_17743,_T_17740,_T_17737,_T_17734,_T_17731,_T_17728,_T_17725,_T_17722,_T_17719}; // @[Cat.scala 29:58]
  wire [36:0] _T_17836 = {_T_17827,_T_17716,_T_17713,_T_17710,_T_17707,_T_17704,_T_17701,_T_17698,_T_17695,_T_17692}; // @[Cat.scala 29:58]
  wire [45:0] _T_17845 = {_T_17836,_T_17689,_T_17686,_T_17683,_T_17680,_T_17677,_T_17674,_T_17671,_T_17668,_T_17665}; // @[Cat.scala 29:58]
  wire [54:0] _T_17854 = {_T_17845,_T_17662,_T_17659,_T_17656,_T_17653,_T_17650,_T_17647,_T_17644,_T_17641,_T_17638}; // @[Cat.scala 29:58]
  wire [62:0] _T_17862 = {_T_17854,_T_17635,_T_17632,_T_17629,_T_17626,_T_17623,_T_17620,_T_17617,_T_17614}; // @[Cat.scala 29:58]
  wire  _T_17930 = io_multiplicand[0] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17933 = io_multiplicand[1] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17936 = io_multiplicand[2] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17939 = io_multiplicand[3] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17942 = io_multiplicand[4] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17945 = io_multiplicand[5] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17948 = io_multiplicand[6] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17951 = io_multiplicand[7] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17954 = io_multiplicand[8] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17957 = io_multiplicand[9] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17960 = io_multiplicand[10] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17963 = io_multiplicand[11] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17966 = io_multiplicand[12] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17969 = io_multiplicand[13] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17972 = io_multiplicand[14] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17975 = io_multiplicand[15] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17978 = io_multiplicand[16] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17981 = io_multiplicand[17] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17984 = io_multiplicand[18] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17987 = io_multiplicand[19] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17990 = io_multiplicand[20] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17993 = io_multiplicand[21] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17996 = io_multiplicand[22] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_17999 = io_multiplicand[23] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18002 = io_multiplicand[24] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18005 = io_multiplicand[25] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18008 = io_multiplicand[26] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18011 = io_multiplicand[27] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18014 = io_multiplicand[28] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18017 = io_multiplicand[29] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18020 = io_multiplicand[30] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18023 = io_multiplicand[31] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18026 = io_multiplicand[32] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18029 = io_multiplicand[33] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18032 = io_multiplicand[34] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18035 = io_multiplicand[35] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18038 = io_multiplicand[36] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18041 = io_multiplicand[37] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18044 = io_multiplicand[38] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18047 = io_multiplicand[39] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18050 = io_multiplicand[40] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18053 = io_multiplicand[41] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18056 = io_multiplicand[42] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18059 = io_multiplicand[43] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18062 = io_multiplicand[44] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18065 = io_multiplicand[45] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18068 = io_multiplicand[46] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18071 = io_multiplicand[47] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18074 = io_multiplicand[48] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18077 = io_multiplicand[49] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18080 = io_multiplicand[50] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18083 = io_multiplicand[51] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18086 = io_multiplicand[52] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18089 = io_multiplicand[53] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18092 = io_multiplicand[54] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18095 = io_multiplicand[55] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18098 = io_multiplicand[56] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18101 = io_multiplicand[57] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18104 = io_multiplicand[58] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18107 = io_multiplicand[59] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18110 = io_multiplicand[60] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18113 = io_multiplicand[61] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18116 = io_multiplicand[62] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire  _T_18119 = io_multiplicand[63] & io_multiplier[56]; // @[partialprod.scala 16:36]
  wire [9:0] _T_18128 = {_T_18119,_T_18116,_T_18113,_T_18110,_T_18107,_T_18104,_T_18101,_T_18098,_T_18095,_T_18092}; // @[Cat.scala 29:58]
  wire [18:0] _T_18137 = {_T_18128,_T_18089,_T_18086,_T_18083,_T_18080,_T_18077,_T_18074,_T_18071,_T_18068,_T_18065}; // @[Cat.scala 29:58]
  wire [27:0] _T_18146 = {_T_18137,_T_18062,_T_18059,_T_18056,_T_18053,_T_18050,_T_18047,_T_18044,_T_18041,_T_18038}; // @[Cat.scala 29:58]
  wire [36:0] _T_18155 = {_T_18146,_T_18035,_T_18032,_T_18029,_T_18026,_T_18023,_T_18020,_T_18017,_T_18014,_T_18011}; // @[Cat.scala 29:58]
  wire [45:0] _T_18164 = {_T_18155,_T_18008,_T_18005,_T_18002,_T_17999,_T_17996,_T_17993,_T_17990,_T_17987,_T_17984}; // @[Cat.scala 29:58]
  wire [54:0] _T_18173 = {_T_18164,_T_17981,_T_17978,_T_17975,_T_17972,_T_17969,_T_17966,_T_17963,_T_17960,_T_17957}; // @[Cat.scala 29:58]
  wire [62:0] _T_18181 = {_T_18173,_T_17954,_T_17951,_T_17948,_T_17945,_T_17942,_T_17939,_T_17936,_T_17933}; // @[Cat.scala 29:58]
  wire  _T_18249 = io_multiplicand[0] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18252 = io_multiplicand[1] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18255 = io_multiplicand[2] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18258 = io_multiplicand[3] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18261 = io_multiplicand[4] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18264 = io_multiplicand[5] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18267 = io_multiplicand[6] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18270 = io_multiplicand[7] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18273 = io_multiplicand[8] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18276 = io_multiplicand[9] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18279 = io_multiplicand[10] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18282 = io_multiplicand[11] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18285 = io_multiplicand[12] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18288 = io_multiplicand[13] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18291 = io_multiplicand[14] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18294 = io_multiplicand[15] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18297 = io_multiplicand[16] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18300 = io_multiplicand[17] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18303 = io_multiplicand[18] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18306 = io_multiplicand[19] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18309 = io_multiplicand[20] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18312 = io_multiplicand[21] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18315 = io_multiplicand[22] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18318 = io_multiplicand[23] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18321 = io_multiplicand[24] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18324 = io_multiplicand[25] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18327 = io_multiplicand[26] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18330 = io_multiplicand[27] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18333 = io_multiplicand[28] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18336 = io_multiplicand[29] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18339 = io_multiplicand[30] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18342 = io_multiplicand[31] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18345 = io_multiplicand[32] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18348 = io_multiplicand[33] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18351 = io_multiplicand[34] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18354 = io_multiplicand[35] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18357 = io_multiplicand[36] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18360 = io_multiplicand[37] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18363 = io_multiplicand[38] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18366 = io_multiplicand[39] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18369 = io_multiplicand[40] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18372 = io_multiplicand[41] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18375 = io_multiplicand[42] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18378 = io_multiplicand[43] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18381 = io_multiplicand[44] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18384 = io_multiplicand[45] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18387 = io_multiplicand[46] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18390 = io_multiplicand[47] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18393 = io_multiplicand[48] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18396 = io_multiplicand[49] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18399 = io_multiplicand[50] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18402 = io_multiplicand[51] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18405 = io_multiplicand[52] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18408 = io_multiplicand[53] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18411 = io_multiplicand[54] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18414 = io_multiplicand[55] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18417 = io_multiplicand[56] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18420 = io_multiplicand[57] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18423 = io_multiplicand[58] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18426 = io_multiplicand[59] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18429 = io_multiplicand[60] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18432 = io_multiplicand[61] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18435 = io_multiplicand[62] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire  _T_18438 = io_multiplicand[63] & io_multiplier[57]; // @[partialprod.scala 16:36]
  wire [9:0] _T_18447 = {_T_18438,_T_18435,_T_18432,_T_18429,_T_18426,_T_18423,_T_18420,_T_18417,_T_18414,_T_18411}; // @[Cat.scala 29:58]
  wire [18:0] _T_18456 = {_T_18447,_T_18408,_T_18405,_T_18402,_T_18399,_T_18396,_T_18393,_T_18390,_T_18387,_T_18384}; // @[Cat.scala 29:58]
  wire [27:0] _T_18465 = {_T_18456,_T_18381,_T_18378,_T_18375,_T_18372,_T_18369,_T_18366,_T_18363,_T_18360,_T_18357}; // @[Cat.scala 29:58]
  wire [36:0] _T_18474 = {_T_18465,_T_18354,_T_18351,_T_18348,_T_18345,_T_18342,_T_18339,_T_18336,_T_18333,_T_18330}; // @[Cat.scala 29:58]
  wire [45:0] _T_18483 = {_T_18474,_T_18327,_T_18324,_T_18321,_T_18318,_T_18315,_T_18312,_T_18309,_T_18306,_T_18303}; // @[Cat.scala 29:58]
  wire [54:0] _T_18492 = {_T_18483,_T_18300,_T_18297,_T_18294,_T_18291,_T_18288,_T_18285,_T_18282,_T_18279,_T_18276}; // @[Cat.scala 29:58]
  wire [62:0] _T_18500 = {_T_18492,_T_18273,_T_18270,_T_18267,_T_18264,_T_18261,_T_18258,_T_18255,_T_18252}; // @[Cat.scala 29:58]
  wire  _T_18568 = io_multiplicand[0] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18571 = io_multiplicand[1] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18574 = io_multiplicand[2] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18577 = io_multiplicand[3] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18580 = io_multiplicand[4] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18583 = io_multiplicand[5] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18586 = io_multiplicand[6] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18589 = io_multiplicand[7] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18592 = io_multiplicand[8] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18595 = io_multiplicand[9] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18598 = io_multiplicand[10] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18601 = io_multiplicand[11] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18604 = io_multiplicand[12] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18607 = io_multiplicand[13] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18610 = io_multiplicand[14] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18613 = io_multiplicand[15] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18616 = io_multiplicand[16] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18619 = io_multiplicand[17] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18622 = io_multiplicand[18] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18625 = io_multiplicand[19] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18628 = io_multiplicand[20] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18631 = io_multiplicand[21] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18634 = io_multiplicand[22] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18637 = io_multiplicand[23] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18640 = io_multiplicand[24] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18643 = io_multiplicand[25] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18646 = io_multiplicand[26] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18649 = io_multiplicand[27] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18652 = io_multiplicand[28] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18655 = io_multiplicand[29] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18658 = io_multiplicand[30] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18661 = io_multiplicand[31] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18664 = io_multiplicand[32] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18667 = io_multiplicand[33] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18670 = io_multiplicand[34] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18673 = io_multiplicand[35] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18676 = io_multiplicand[36] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18679 = io_multiplicand[37] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18682 = io_multiplicand[38] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18685 = io_multiplicand[39] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18688 = io_multiplicand[40] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18691 = io_multiplicand[41] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18694 = io_multiplicand[42] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18697 = io_multiplicand[43] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18700 = io_multiplicand[44] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18703 = io_multiplicand[45] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18706 = io_multiplicand[46] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18709 = io_multiplicand[47] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18712 = io_multiplicand[48] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18715 = io_multiplicand[49] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18718 = io_multiplicand[50] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18721 = io_multiplicand[51] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18724 = io_multiplicand[52] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18727 = io_multiplicand[53] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18730 = io_multiplicand[54] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18733 = io_multiplicand[55] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18736 = io_multiplicand[56] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18739 = io_multiplicand[57] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18742 = io_multiplicand[58] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18745 = io_multiplicand[59] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18748 = io_multiplicand[60] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18751 = io_multiplicand[61] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18754 = io_multiplicand[62] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire  _T_18757 = io_multiplicand[63] & io_multiplier[58]; // @[partialprod.scala 16:36]
  wire [9:0] _T_18766 = {_T_18757,_T_18754,_T_18751,_T_18748,_T_18745,_T_18742,_T_18739,_T_18736,_T_18733,_T_18730}; // @[Cat.scala 29:58]
  wire [18:0] _T_18775 = {_T_18766,_T_18727,_T_18724,_T_18721,_T_18718,_T_18715,_T_18712,_T_18709,_T_18706,_T_18703}; // @[Cat.scala 29:58]
  wire [27:0] _T_18784 = {_T_18775,_T_18700,_T_18697,_T_18694,_T_18691,_T_18688,_T_18685,_T_18682,_T_18679,_T_18676}; // @[Cat.scala 29:58]
  wire [36:0] _T_18793 = {_T_18784,_T_18673,_T_18670,_T_18667,_T_18664,_T_18661,_T_18658,_T_18655,_T_18652,_T_18649}; // @[Cat.scala 29:58]
  wire [45:0] _T_18802 = {_T_18793,_T_18646,_T_18643,_T_18640,_T_18637,_T_18634,_T_18631,_T_18628,_T_18625,_T_18622}; // @[Cat.scala 29:58]
  wire [54:0] _T_18811 = {_T_18802,_T_18619,_T_18616,_T_18613,_T_18610,_T_18607,_T_18604,_T_18601,_T_18598,_T_18595}; // @[Cat.scala 29:58]
  wire [62:0] _T_18819 = {_T_18811,_T_18592,_T_18589,_T_18586,_T_18583,_T_18580,_T_18577,_T_18574,_T_18571}; // @[Cat.scala 29:58]
  wire  _T_18887 = io_multiplicand[0] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18890 = io_multiplicand[1] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18893 = io_multiplicand[2] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18896 = io_multiplicand[3] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18899 = io_multiplicand[4] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18902 = io_multiplicand[5] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18905 = io_multiplicand[6] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18908 = io_multiplicand[7] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18911 = io_multiplicand[8] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18914 = io_multiplicand[9] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18917 = io_multiplicand[10] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18920 = io_multiplicand[11] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18923 = io_multiplicand[12] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18926 = io_multiplicand[13] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18929 = io_multiplicand[14] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18932 = io_multiplicand[15] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18935 = io_multiplicand[16] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18938 = io_multiplicand[17] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18941 = io_multiplicand[18] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18944 = io_multiplicand[19] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18947 = io_multiplicand[20] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18950 = io_multiplicand[21] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18953 = io_multiplicand[22] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18956 = io_multiplicand[23] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18959 = io_multiplicand[24] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18962 = io_multiplicand[25] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18965 = io_multiplicand[26] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18968 = io_multiplicand[27] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18971 = io_multiplicand[28] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18974 = io_multiplicand[29] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18977 = io_multiplicand[30] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18980 = io_multiplicand[31] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18983 = io_multiplicand[32] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18986 = io_multiplicand[33] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18989 = io_multiplicand[34] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18992 = io_multiplicand[35] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18995 = io_multiplicand[36] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_18998 = io_multiplicand[37] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19001 = io_multiplicand[38] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19004 = io_multiplicand[39] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19007 = io_multiplicand[40] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19010 = io_multiplicand[41] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19013 = io_multiplicand[42] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19016 = io_multiplicand[43] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19019 = io_multiplicand[44] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19022 = io_multiplicand[45] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19025 = io_multiplicand[46] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19028 = io_multiplicand[47] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19031 = io_multiplicand[48] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19034 = io_multiplicand[49] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19037 = io_multiplicand[50] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19040 = io_multiplicand[51] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19043 = io_multiplicand[52] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19046 = io_multiplicand[53] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19049 = io_multiplicand[54] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19052 = io_multiplicand[55] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19055 = io_multiplicand[56] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19058 = io_multiplicand[57] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19061 = io_multiplicand[58] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19064 = io_multiplicand[59] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19067 = io_multiplicand[60] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19070 = io_multiplicand[61] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19073 = io_multiplicand[62] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire  _T_19076 = io_multiplicand[63] & io_multiplier[59]; // @[partialprod.scala 16:36]
  wire [9:0] _T_19085 = {_T_19076,_T_19073,_T_19070,_T_19067,_T_19064,_T_19061,_T_19058,_T_19055,_T_19052,_T_19049}; // @[Cat.scala 29:58]
  wire [18:0] _T_19094 = {_T_19085,_T_19046,_T_19043,_T_19040,_T_19037,_T_19034,_T_19031,_T_19028,_T_19025,_T_19022}; // @[Cat.scala 29:58]
  wire [27:0] _T_19103 = {_T_19094,_T_19019,_T_19016,_T_19013,_T_19010,_T_19007,_T_19004,_T_19001,_T_18998,_T_18995}; // @[Cat.scala 29:58]
  wire [36:0] _T_19112 = {_T_19103,_T_18992,_T_18989,_T_18986,_T_18983,_T_18980,_T_18977,_T_18974,_T_18971,_T_18968}; // @[Cat.scala 29:58]
  wire [45:0] _T_19121 = {_T_19112,_T_18965,_T_18962,_T_18959,_T_18956,_T_18953,_T_18950,_T_18947,_T_18944,_T_18941}; // @[Cat.scala 29:58]
  wire [54:0] _T_19130 = {_T_19121,_T_18938,_T_18935,_T_18932,_T_18929,_T_18926,_T_18923,_T_18920,_T_18917,_T_18914}; // @[Cat.scala 29:58]
  wire [62:0] _T_19138 = {_T_19130,_T_18911,_T_18908,_T_18905,_T_18902,_T_18899,_T_18896,_T_18893,_T_18890}; // @[Cat.scala 29:58]
  wire  _T_19206 = io_multiplicand[0] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19209 = io_multiplicand[1] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19212 = io_multiplicand[2] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19215 = io_multiplicand[3] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19218 = io_multiplicand[4] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19221 = io_multiplicand[5] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19224 = io_multiplicand[6] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19227 = io_multiplicand[7] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19230 = io_multiplicand[8] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19233 = io_multiplicand[9] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19236 = io_multiplicand[10] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19239 = io_multiplicand[11] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19242 = io_multiplicand[12] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19245 = io_multiplicand[13] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19248 = io_multiplicand[14] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19251 = io_multiplicand[15] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19254 = io_multiplicand[16] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19257 = io_multiplicand[17] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19260 = io_multiplicand[18] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19263 = io_multiplicand[19] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19266 = io_multiplicand[20] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19269 = io_multiplicand[21] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19272 = io_multiplicand[22] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19275 = io_multiplicand[23] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19278 = io_multiplicand[24] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19281 = io_multiplicand[25] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19284 = io_multiplicand[26] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19287 = io_multiplicand[27] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19290 = io_multiplicand[28] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19293 = io_multiplicand[29] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19296 = io_multiplicand[30] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19299 = io_multiplicand[31] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19302 = io_multiplicand[32] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19305 = io_multiplicand[33] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19308 = io_multiplicand[34] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19311 = io_multiplicand[35] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19314 = io_multiplicand[36] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19317 = io_multiplicand[37] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19320 = io_multiplicand[38] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19323 = io_multiplicand[39] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19326 = io_multiplicand[40] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19329 = io_multiplicand[41] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19332 = io_multiplicand[42] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19335 = io_multiplicand[43] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19338 = io_multiplicand[44] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19341 = io_multiplicand[45] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19344 = io_multiplicand[46] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19347 = io_multiplicand[47] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19350 = io_multiplicand[48] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19353 = io_multiplicand[49] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19356 = io_multiplicand[50] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19359 = io_multiplicand[51] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19362 = io_multiplicand[52] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19365 = io_multiplicand[53] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19368 = io_multiplicand[54] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19371 = io_multiplicand[55] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19374 = io_multiplicand[56] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19377 = io_multiplicand[57] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19380 = io_multiplicand[58] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19383 = io_multiplicand[59] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19386 = io_multiplicand[60] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19389 = io_multiplicand[61] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19392 = io_multiplicand[62] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire  _T_19395 = io_multiplicand[63] & io_multiplier[60]; // @[partialprod.scala 16:36]
  wire [9:0] _T_19404 = {_T_19395,_T_19392,_T_19389,_T_19386,_T_19383,_T_19380,_T_19377,_T_19374,_T_19371,_T_19368}; // @[Cat.scala 29:58]
  wire [18:0] _T_19413 = {_T_19404,_T_19365,_T_19362,_T_19359,_T_19356,_T_19353,_T_19350,_T_19347,_T_19344,_T_19341}; // @[Cat.scala 29:58]
  wire [27:0] _T_19422 = {_T_19413,_T_19338,_T_19335,_T_19332,_T_19329,_T_19326,_T_19323,_T_19320,_T_19317,_T_19314}; // @[Cat.scala 29:58]
  wire [36:0] _T_19431 = {_T_19422,_T_19311,_T_19308,_T_19305,_T_19302,_T_19299,_T_19296,_T_19293,_T_19290,_T_19287}; // @[Cat.scala 29:58]
  wire [45:0] _T_19440 = {_T_19431,_T_19284,_T_19281,_T_19278,_T_19275,_T_19272,_T_19269,_T_19266,_T_19263,_T_19260}; // @[Cat.scala 29:58]
  wire [54:0] _T_19449 = {_T_19440,_T_19257,_T_19254,_T_19251,_T_19248,_T_19245,_T_19242,_T_19239,_T_19236,_T_19233}; // @[Cat.scala 29:58]
  wire [62:0] _T_19457 = {_T_19449,_T_19230,_T_19227,_T_19224,_T_19221,_T_19218,_T_19215,_T_19212,_T_19209}; // @[Cat.scala 29:58]
  wire  _T_19525 = io_multiplicand[0] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19528 = io_multiplicand[1] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19531 = io_multiplicand[2] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19534 = io_multiplicand[3] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19537 = io_multiplicand[4] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19540 = io_multiplicand[5] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19543 = io_multiplicand[6] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19546 = io_multiplicand[7] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19549 = io_multiplicand[8] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19552 = io_multiplicand[9] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19555 = io_multiplicand[10] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19558 = io_multiplicand[11] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19561 = io_multiplicand[12] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19564 = io_multiplicand[13] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19567 = io_multiplicand[14] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19570 = io_multiplicand[15] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19573 = io_multiplicand[16] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19576 = io_multiplicand[17] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19579 = io_multiplicand[18] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19582 = io_multiplicand[19] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19585 = io_multiplicand[20] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19588 = io_multiplicand[21] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19591 = io_multiplicand[22] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19594 = io_multiplicand[23] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19597 = io_multiplicand[24] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19600 = io_multiplicand[25] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19603 = io_multiplicand[26] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19606 = io_multiplicand[27] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19609 = io_multiplicand[28] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19612 = io_multiplicand[29] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19615 = io_multiplicand[30] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19618 = io_multiplicand[31] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19621 = io_multiplicand[32] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19624 = io_multiplicand[33] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19627 = io_multiplicand[34] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19630 = io_multiplicand[35] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19633 = io_multiplicand[36] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19636 = io_multiplicand[37] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19639 = io_multiplicand[38] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19642 = io_multiplicand[39] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19645 = io_multiplicand[40] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19648 = io_multiplicand[41] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19651 = io_multiplicand[42] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19654 = io_multiplicand[43] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19657 = io_multiplicand[44] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19660 = io_multiplicand[45] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19663 = io_multiplicand[46] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19666 = io_multiplicand[47] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19669 = io_multiplicand[48] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19672 = io_multiplicand[49] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19675 = io_multiplicand[50] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19678 = io_multiplicand[51] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19681 = io_multiplicand[52] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19684 = io_multiplicand[53] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19687 = io_multiplicand[54] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19690 = io_multiplicand[55] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19693 = io_multiplicand[56] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19696 = io_multiplicand[57] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19699 = io_multiplicand[58] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19702 = io_multiplicand[59] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19705 = io_multiplicand[60] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19708 = io_multiplicand[61] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19711 = io_multiplicand[62] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire  _T_19714 = io_multiplicand[63] & io_multiplier[61]; // @[partialprod.scala 16:36]
  wire [9:0] _T_19723 = {_T_19714,_T_19711,_T_19708,_T_19705,_T_19702,_T_19699,_T_19696,_T_19693,_T_19690,_T_19687}; // @[Cat.scala 29:58]
  wire [18:0] _T_19732 = {_T_19723,_T_19684,_T_19681,_T_19678,_T_19675,_T_19672,_T_19669,_T_19666,_T_19663,_T_19660}; // @[Cat.scala 29:58]
  wire [27:0] _T_19741 = {_T_19732,_T_19657,_T_19654,_T_19651,_T_19648,_T_19645,_T_19642,_T_19639,_T_19636,_T_19633}; // @[Cat.scala 29:58]
  wire [36:0] _T_19750 = {_T_19741,_T_19630,_T_19627,_T_19624,_T_19621,_T_19618,_T_19615,_T_19612,_T_19609,_T_19606}; // @[Cat.scala 29:58]
  wire [45:0] _T_19759 = {_T_19750,_T_19603,_T_19600,_T_19597,_T_19594,_T_19591,_T_19588,_T_19585,_T_19582,_T_19579}; // @[Cat.scala 29:58]
  wire [54:0] _T_19768 = {_T_19759,_T_19576,_T_19573,_T_19570,_T_19567,_T_19564,_T_19561,_T_19558,_T_19555,_T_19552}; // @[Cat.scala 29:58]
  wire [62:0] _T_19776 = {_T_19768,_T_19549,_T_19546,_T_19543,_T_19540,_T_19537,_T_19534,_T_19531,_T_19528}; // @[Cat.scala 29:58]
  wire  _T_19844 = io_multiplicand[0] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19847 = io_multiplicand[1] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19850 = io_multiplicand[2] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19853 = io_multiplicand[3] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19856 = io_multiplicand[4] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19859 = io_multiplicand[5] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19862 = io_multiplicand[6] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19865 = io_multiplicand[7] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19868 = io_multiplicand[8] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19871 = io_multiplicand[9] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19874 = io_multiplicand[10] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19877 = io_multiplicand[11] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19880 = io_multiplicand[12] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19883 = io_multiplicand[13] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19886 = io_multiplicand[14] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19889 = io_multiplicand[15] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19892 = io_multiplicand[16] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19895 = io_multiplicand[17] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19898 = io_multiplicand[18] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19901 = io_multiplicand[19] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19904 = io_multiplicand[20] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19907 = io_multiplicand[21] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19910 = io_multiplicand[22] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19913 = io_multiplicand[23] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19916 = io_multiplicand[24] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19919 = io_multiplicand[25] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19922 = io_multiplicand[26] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19925 = io_multiplicand[27] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19928 = io_multiplicand[28] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19931 = io_multiplicand[29] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19934 = io_multiplicand[30] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19937 = io_multiplicand[31] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19940 = io_multiplicand[32] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19943 = io_multiplicand[33] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19946 = io_multiplicand[34] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19949 = io_multiplicand[35] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19952 = io_multiplicand[36] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19955 = io_multiplicand[37] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19958 = io_multiplicand[38] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19961 = io_multiplicand[39] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19964 = io_multiplicand[40] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19967 = io_multiplicand[41] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19970 = io_multiplicand[42] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19973 = io_multiplicand[43] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19976 = io_multiplicand[44] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19979 = io_multiplicand[45] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19982 = io_multiplicand[46] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19985 = io_multiplicand[47] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19988 = io_multiplicand[48] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19991 = io_multiplicand[49] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19994 = io_multiplicand[50] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_19997 = io_multiplicand[51] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_20000 = io_multiplicand[52] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_20003 = io_multiplicand[53] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_20006 = io_multiplicand[54] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_20009 = io_multiplicand[55] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_20012 = io_multiplicand[56] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_20015 = io_multiplicand[57] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_20018 = io_multiplicand[58] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_20021 = io_multiplicand[59] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_20024 = io_multiplicand[60] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_20027 = io_multiplicand[61] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_20030 = io_multiplicand[62] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire  _T_20033 = io_multiplicand[63] & io_multiplier[62]; // @[partialprod.scala 16:36]
  wire [9:0] _T_20042 = {_T_20033,_T_20030,_T_20027,_T_20024,_T_20021,_T_20018,_T_20015,_T_20012,_T_20009,_T_20006}; // @[Cat.scala 29:58]
  wire [18:0] _T_20051 = {_T_20042,_T_20003,_T_20000,_T_19997,_T_19994,_T_19991,_T_19988,_T_19985,_T_19982,_T_19979}; // @[Cat.scala 29:58]
  wire [27:0] _T_20060 = {_T_20051,_T_19976,_T_19973,_T_19970,_T_19967,_T_19964,_T_19961,_T_19958,_T_19955,_T_19952}; // @[Cat.scala 29:58]
  wire [36:0] _T_20069 = {_T_20060,_T_19949,_T_19946,_T_19943,_T_19940,_T_19937,_T_19934,_T_19931,_T_19928,_T_19925}; // @[Cat.scala 29:58]
  wire [45:0] _T_20078 = {_T_20069,_T_19922,_T_19919,_T_19916,_T_19913,_T_19910,_T_19907,_T_19904,_T_19901,_T_19898}; // @[Cat.scala 29:58]
  wire [54:0] _T_20087 = {_T_20078,_T_19895,_T_19892,_T_19889,_T_19886,_T_19883,_T_19880,_T_19877,_T_19874,_T_19871}; // @[Cat.scala 29:58]
  wire [62:0] _T_20095 = {_T_20087,_T_19868,_T_19865,_T_19862,_T_19859,_T_19856,_T_19853,_T_19850,_T_19847}; // @[Cat.scala 29:58]
  wire  _T_20163 = io_multiplicand[0] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20166 = io_multiplicand[1] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20169 = io_multiplicand[2] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20172 = io_multiplicand[3] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20175 = io_multiplicand[4] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20178 = io_multiplicand[5] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20181 = io_multiplicand[6] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20184 = io_multiplicand[7] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20187 = io_multiplicand[8] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20190 = io_multiplicand[9] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20193 = io_multiplicand[10] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20196 = io_multiplicand[11] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20199 = io_multiplicand[12] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20202 = io_multiplicand[13] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20205 = io_multiplicand[14] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20208 = io_multiplicand[15] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20211 = io_multiplicand[16] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20214 = io_multiplicand[17] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20217 = io_multiplicand[18] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20220 = io_multiplicand[19] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20223 = io_multiplicand[20] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20226 = io_multiplicand[21] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20229 = io_multiplicand[22] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20232 = io_multiplicand[23] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20235 = io_multiplicand[24] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20238 = io_multiplicand[25] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20241 = io_multiplicand[26] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20244 = io_multiplicand[27] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20247 = io_multiplicand[28] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20250 = io_multiplicand[29] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20253 = io_multiplicand[30] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20256 = io_multiplicand[31] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20259 = io_multiplicand[32] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20262 = io_multiplicand[33] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20265 = io_multiplicand[34] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20268 = io_multiplicand[35] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20271 = io_multiplicand[36] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20274 = io_multiplicand[37] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20277 = io_multiplicand[38] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20280 = io_multiplicand[39] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20283 = io_multiplicand[40] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20286 = io_multiplicand[41] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20289 = io_multiplicand[42] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20292 = io_multiplicand[43] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20295 = io_multiplicand[44] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20298 = io_multiplicand[45] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20301 = io_multiplicand[46] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20304 = io_multiplicand[47] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20307 = io_multiplicand[48] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20310 = io_multiplicand[49] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20313 = io_multiplicand[50] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20316 = io_multiplicand[51] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20319 = io_multiplicand[52] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20322 = io_multiplicand[53] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20325 = io_multiplicand[54] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20328 = io_multiplicand[55] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20331 = io_multiplicand[56] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20334 = io_multiplicand[57] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20337 = io_multiplicand[58] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20340 = io_multiplicand[59] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20343 = io_multiplicand[60] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20346 = io_multiplicand[61] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20349 = io_multiplicand[62] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire  _T_20352 = io_multiplicand[63] & io_multiplier[63]; // @[partialprod.scala 16:36]
  wire [9:0] _T_20361 = {_T_20352,_T_20349,_T_20346,_T_20343,_T_20340,_T_20337,_T_20334,_T_20331,_T_20328,_T_20325}; // @[Cat.scala 29:58]
  wire [18:0] _T_20370 = {_T_20361,_T_20322,_T_20319,_T_20316,_T_20313,_T_20310,_T_20307,_T_20304,_T_20301,_T_20298}; // @[Cat.scala 29:58]
  wire [27:0] _T_20379 = {_T_20370,_T_20295,_T_20292,_T_20289,_T_20286,_T_20283,_T_20280,_T_20277,_T_20274,_T_20271}; // @[Cat.scala 29:58]
  wire [36:0] _T_20388 = {_T_20379,_T_20268,_T_20265,_T_20262,_T_20259,_T_20256,_T_20253,_T_20250,_T_20247,_T_20244}; // @[Cat.scala 29:58]
  wire [45:0] _T_20397 = {_T_20388,_T_20241,_T_20238,_T_20235,_T_20232,_T_20229,_T_20226,_T_20223,_T_20220,_T_20217}; // @[Cat.scala 29:58]
  wire [54:0] _T_20406 = {_T_20397,_T_20214,_T_20211,_T_20208,_T_20205,_T_20202,_T_20199,_T_20196,_T_20193,_T_20190}; // @[Cat.scala 29:58]
  wire [62:0] _T_20414 = {_T_20406,_T_20187,_T_20184,_T_20181,_T_20178,_T_20175,_T_20172,_T_20169,_T_20166}; // @[Cat.scala 29:58]
  assign io_outs_0 = {_T_317,_T_66}; // @[partialprod.scala 18:16]
  assign io_outs_1 = {_T_636,_T_385}; // @[partialprod.scala 18:16]
  assign io_outs_2 = {_T_955,_T_704}; // @[partialprod.scala 18:16]
  assign io_outs_3 = {_T_1274,_T_1023}; // @[partialprod.scala 18:16]
  assign io_outs_4 = {_T_1593,_T_1342}; // @[partialprod.scala 18:16]
  assign io_outs_5 = {_T_1912,_T_1661}; // @[partialprod.scala 18:16]
  assign io_outs_6 = {_T_2231,_T_1980}; // @[partialprod.scala 18:16]
  assign io_outs_7 = {_T_2550,_T_2299}; // @[partialprod.scala 18:16]
  assign io_outs_8 = {_T_2869,_T_2618}; // @[partialprod.scala 18:16]
  assign io_outs_9 = {_T_3188,_T_2937}; // @[partialprod.scala 18:16]
  assign io_outs_10 = {_T_3507,_T_3256}; // @[partialprod.scala 18:16]
  assign io_outs_11 = {_T_3826,_T_3575}; // @[partialprod.scala 18:16]
  assign io_outs_12 = {_T_4145,_T_3894}; // @[partialprod.scala 18:16]
  assign io_outs_13 = {_T_4464,_T_4213}; // @[partialprod.scala 18:16]
  assign io_outs_14 = {_T_4783,_T_4532}; // @[partialprod.scala 18:16]
  assign io_outs_15 = {_T_5102,_T_4851}; // @[partialprod.scala 18:16]
  assign io_outs_16 = {_T_5421,_T_5170}; // @[partialprod.scala 18:16]
  assign io_outs_17 = {_T_5740,_T_5489}; // @[partialprod.scala 18:16]
  assign io_outs_18 = {_T_6059,_T_5808}; // @[partialprod.scala 18:16]
  assign io_outs_19 = {_T_6378,_T_6127}; // @[partialprod.scala 18:16]
  assign io_outs_20 = {_T_6697,_T_6446}; // @[partialprod.scala 18:16]
  assign io_outs_21 = {_T_7016,_T_6765}; // @[partialprod.scala 18:16]
  assign io_outs_22 = {_T_7335,_T_7084}; // @[partialprod.scala 18:16]
  assign io_outs_23 = {_T_7654,_T_7403}; // @[partialprod.scala 18:16]
  assign io_outs_24 = {_T_7973,_T_7722}; // @[partialprod.scala 18:16]
  assign io_outs_25 = {_T_8292,_T_8041}; // @[partialprod.scala 18:16]
  assign io_outs_26 = {_T_8611,_T_8360}; // @[partialprod.scala 18:16]
  assign io_outs_27 = {_T_8930,_T_8679}; // @[partialprod.scala 18:16]
  assign io_outs_28 = {_T_9249,_T_8998}; // @[partialprod.scala 18:16]
  assign io_outs_29 = {_T_9568,_T_9317}; // @[partialprod.scala 18:16]
  assign io_outs_30 = {_T_9887,_T_9636}; // @[partialprod.scala 18:16]
  assign io_outs_31 = {_T_10206,_T_9955}; // @[partialprod.scala 18:16]
  assign io_outs_32 = {_T_10525,_T_10274}; // @[partialprod.scala 18:16]
  assign io_outs_33 = {_T_10844,_T_10593}; // @[partialprod.scala 18:16]
  assign io_outs_34 = {_T_11163,_T_10912}; // @[partialprod.scala 18:16]
  assign io_outs_35 = {_T_11482,_T_11231}; // @[partialprod.scala 18:16]
  assign io_outs_36 = {_T_11801,_T_11550}; // @[partialprod.scala 18:16]
  assign io_outs_37 = {_T_12120,_T_11869}; // @[partialprod.scala 18:16]
  assign io_outs_38 = {_T_12439,_T_12188}; // @[partialprod.scala 18:16]
  assign io_outs_39 = {_T_12758,_T_12507}; // @[partialprod.scala 18:16]
  assign io_outs_40 = {_T_13077,_T_12826}; // @[partialprod.scala 18:16]
  assign io_outs_41 = {_T_13396,_T_13145}; // @[partialprod.scala 18:16]
  assign io_outs_42 = {_T_13715,_T_13464}; // @[partialprod.scala 18:16]
  assign io_outs_43 = {_T_14034,_T_13783}; // @[partialprod.scala 18:16]
  assign io_outs_44 = {_T_14353,_T_14102}; // @[partialprod.scala 18:16]
  assign io_outs_45 = {_T_14672,_T_14421}; // @[partialprod.scala 18:16]
  assign io_outs_46 = {_T_14991,_T_14740}; // @[partialprod.scala 18:16]
  assign io_outs_47 = {_T_15310,_T_15059}; // @[partialprod.scala 18:16]
  assign io_outs_48 = {_T_15629,_T_15378}; // @[partialprod.scala 18:16]
  assign io_outs_49 = {_T_15948,_T_15697}; // @[partialprod.scala 18:16]
  assign io_outs_50 = {_T_16267,_T_16016}; // @[partialprod.scala 18:16]
  assign io_outs_51 = {_T_16586,_T_16335}; // @[partialprod.scala 18:16]
  assign io_outs_52 = {_T_16905,_T_16654}; // @[partialprod.scala 18:16]
  assign io_outs_53 = {_T_17224,_T_16973}; // @[partialprod.scala 18:16]
  assign io_outs_54 = {_T_17543,_T_17292}; // @[partialprod.scala 18:16]
  assign io_outs_55 = {_T_17862,_T_17611}; // @[partialprod.scala 18:16]
  assign io_outs_56 = {_T_18181,_T_17930}; // @[partialprod.scala 18:16]
  assign io_outs_57 = {_T_18500,_T_18249}; // @[partialprod.scala 18:16]
  assign io_outs_58 = {_T_18819,_T_18568}; // @[partialprod.scala 18:16]
  assign io_outs_59 = {_T_19138,_T_18887}; // @[partialprod.scala 18:16]
  assign io_outs_60 = {_T_19457,_T_19206}; // @[partialprod.scala 18:16]
  assign io_outs_61 = {_T_19776,_T_19525}; // @[partialprod.scala 18:16]
  assign io_outs_62 = {_T_20095,_T_19844}; // @[partialprod.scala 18:16]
  assign io_outs_63 = {_T_20414,_T_20163}; // @[partialprod.scala 18:16]
endmodule
module HalfAdder(
  input   io_a,
  input   io_b,
  output  io_s,
  output  io_co
);
  assign io_s = io_a ^ io_b; // @[comp.scala 15:8]
  assign io_co = io_a & io_b; // @[comp.scala 16:9]
endmodule
module FullAdder(
  input   io_a,
  input   io_b,
  input   io_ci,
  output  io_s,
  output  io_co
);
  wire  a_xor_b = io_a ^ io_b; // @[comp.scala 28:22]
  wire  a_and_b = io_a & io_b; // @[comp.scala 31:22]
  wire  a_and_cin = io_a & io_ci; // @[comp.scala 32:24]
  wire  b_and_cin = io_b & io_ci; // @[comp.scala 33:24]
  wire  _T_1 = a_and_b | b_and_cin; // @[comp.scala 34:20]
  assign io_s = a_xor_b ^ io_ci; // @[comp.scala 29:8]
  assign io_co = _T_1 | a_and_cin; // @[comp.scala 34:9]
endmodule
module Wallace(
  input  [63:0]  io_pp_0,
  input  [63:0]  io_pp_1,
  input  [63:0]  io_pp_2,
  input  [63:0]  io_pp_3,
  input  [63:0]  io_pp_4,
  input  [63:0]  io_pp_5,
  input  [63:0]  io_pp_6,
  input  [63:0]  io_pp_7,
  input  [63:0]  io_pp_8,
  input  [63:0]  io_pp_9,
  input  [63:0]  io_pp_10,
  input  [63:0]  io_pp_11,
  input  [63:0]  io_pp_12,
  input  [63:0]  io_pp_13,
  input  [63:0]  io_pp_14,
  input  [63:0]  io_pp_15,
  input  [63:0]  io_pp_16,
  input  [63:0]  io_pp_17,
  input  [63:0]  io_pp_18,
  input  [63:0]  io_pp_19,
  input  [63:0]  io_pp_20,
  input  [63:0]  io_pp_21,
  input  [63:0]  io_pp_22,
  input  [63:0]  io_pp_23,
  input  [63:0]  io_pp_24,
  input  [63:0]  io_pp_25,
  input  [63:0]  io_pp_26,
  input  [63:0]  io_pp_27,
  input  [63:0]  io_pp_28,
  input  [63:0]  io_pp_29,
  input  [63:0]  io_pp_30,
  input  [63:0]  io_pp_31,
  input  [63:0]  io_pp_32,
  input  [63:0]  io_pp_33,
  input  [63:0]  io_pp_34,
  input  [63:0]  io_pp_35,
  input  [63:0]  io_pp_36,
  input  [63:0]  io_pp_37,
  input  [63:0]  io_pp_38,
  input  [63:0]  io_pp_39,
  input  [63:0]  io_pp_40,
  input  [63:0]  io_pp_41,
  input  [63:0]  io_pp_42,
  input  [63:0]  io_pp_43,
  input  [63:0]  io_pp_44,
  input  [63:0]  io_pp_45,
  input  [63:0]  io_pp_46,
  input  [63:0]  io_pp_47,
  input  [63:0]  io_pp_48,
  input  [63:0]  io_pp_49,
  input  [63:0]  io_pp_50,
  input  [63:0]  io_pp_51,
  input  [63:0]  io_pp_52,
  input  [63:0]  io_pp_53,
  input  [63:0]  io_pp_54,
  input  [63:0]  io_pp_55,
  input  [63:0]  io_pp_56,
  input  [63:0]  io_pp_57,
  input  [63:0]  io_pp_58,
  input  [63:0]  io_pp_59,
  input  [63:0]  io_pp_60,
  input  [63:0]  io_pp_61,
  input  [63:0]  io_pp_62,
  input  [63:0]  io_pp_63,
  output [127:0] io_augend,
  output [127:0] io_addend
);
  wire  HalfAdder_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_1_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_1_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_1_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_1_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_4_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_4_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_4_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_4_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_4_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_5_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_5_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_5_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_5_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_5_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_6_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_6_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_6_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_6_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_6_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_7_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_7_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_7_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_7_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_7_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_8_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_8_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_8_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_8_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_8_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_2_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_2_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_2_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_2_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_9_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_9_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_9_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_9_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_9_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_10_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_10_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_10_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_10_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_10_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_11_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_11_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_11_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_11_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_11_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_12_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_12_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_12_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_12_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_12_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_13_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_13_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_13_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_13_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_13_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_14_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_14_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_14_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_14_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_14_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_15_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_15_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_15_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_15_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_15_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_16_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_16_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_16_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_16_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_16_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_17_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_17_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_17_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_17_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_17_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_3_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_3_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_3_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_3_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_18_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_18_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_18_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_18_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_18_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_19_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_19_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_19_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_19_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_19_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_20_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_20_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_20_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_20_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_20_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_21_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_21_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_21_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_21_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_21_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_22_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_22_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_22_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_22_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_22_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_23_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_23_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_23_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_23_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_23_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_24_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_24_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_24_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_24_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_24_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_25_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_25_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_25_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_25_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_25_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_26_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_26_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_26_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_26_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_26_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_27_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_27_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_27_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_27_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_27_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_28_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_28_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_28_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_28_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_28_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_29_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_29_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_29_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_29_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_29_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_30_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_30_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_30_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_30_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_30_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_31_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_31_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_31_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_31_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_31_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_32_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_32_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_32_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_32_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_32_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_33_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_33_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_33_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_33_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_33_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_34_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_34_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_34_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_34_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_34_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_35_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_35_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_35_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_35_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_35_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_36_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_36_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_36_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_36_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_36_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_37_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_37_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_37_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_37_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_37_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_38_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_38_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_38_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_38_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_38_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_39_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_39_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_39_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_39_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_39_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_40_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_40_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_40_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_40_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_40_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_41_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_41_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_41_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_41_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_41_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_42_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_42_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_42_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_42_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_42_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_43_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_43_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_43_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_43_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_43_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_44_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_44_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_44_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_44_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_44_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_4_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_4_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_4_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_4_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_45_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_45_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_45_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_45_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_45_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_46_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_46_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_46_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_46_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_46_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_47_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_47_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_47_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_47_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_47_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_48_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_48_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_48_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_48_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_48_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_49_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_49_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_49_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_49_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_49_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_50_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_50_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_50_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_50_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_50_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_51_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_51_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_51_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_51_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_51_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_52_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_52_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_52_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_52_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_52_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_53_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_53_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_53_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_53_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_53_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_54_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_54_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_54_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_54_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_54_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_55_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_55_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_55_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_55_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_55_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_56_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_56_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_56_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_56_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_56_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_57_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_57_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_57_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_57_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_57_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_58_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_58_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_58_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_58_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_58_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_59_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_59_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_59_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_59_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_59_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_60_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_60_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_60_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_60_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_60_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_61_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_61_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_61_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_61_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_61_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_62_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_62_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_62_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_62_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_62_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_5_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_5_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_5_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_5_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_63_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_63_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_63_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_63_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_63_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_64_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_64_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_64_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_64_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_64_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_65_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_65_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_65_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_65_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_65_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_66_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_66_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_66_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_66_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_66_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_67_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_67_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_67_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_67_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_67_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_68_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_68_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_68_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_68_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_68_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_69_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_69_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_69_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_69_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_69_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_70_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_70_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_70_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_70_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_70_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_71_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_71_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_71_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_71_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_71_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_72_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_72_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_72_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_72_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_72_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_73_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_73_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_73_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_73_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_73_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_74_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_74_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_74_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_74_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_74_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_75_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_75_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_75_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_75_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_75_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_76_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_76_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_76_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_76_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_76_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_77_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_77_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_77_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_77_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_77_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_78_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_78_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_78_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_78_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_78_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_79_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_79_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_79_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_79_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_79_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_80_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_80_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_80_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_80_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_80_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_81_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_81_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_81_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_81_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_81_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_82_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_82_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_82_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_82_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_82_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_83_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_83_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_83_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_83_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_83_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_6_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_6_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_6_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_6_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_84_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_84_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_84_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_84_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_84_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_85_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_85_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_85_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_85_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_85_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_86_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_86_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_86_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_86_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_86_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_87_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_87_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_87_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_87_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_87_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_88_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_88_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_88_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_88_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_88_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_89_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_89_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_89_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_89_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_89_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_90_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_90_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_90_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_90_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_90_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_91_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_91_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_91_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_91_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_91_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_92_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_92_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_92_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_92_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_92_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_93_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_93_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_93_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_93_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_93_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_94_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_94_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_94_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_94_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_94_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_95_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_95_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_95_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_95_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_95_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_96_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_96_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_96_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_96_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_96_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_97_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_97_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_97_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_97_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_97_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_98_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_98_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_98_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_98_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_98_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_99_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_99_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_99_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_99_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_99_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_100_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_100_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_100_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_100_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_100_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_101_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_101_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_101_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_101_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_101_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_102_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_102_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_102_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_102_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_102_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_103_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_103_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_103_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_103_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_103_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_104_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_104_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_104_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_104_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_104_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_105_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_105_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_105_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_105_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_105_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_106_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_106_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_106_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_106_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_106_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_107_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_107_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_107_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_107_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_107_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_108_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_108_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_108_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_108_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_108_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_109_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_109_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_109_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_109_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_109_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_110_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_110_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_110_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_110_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_110_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_111_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_111_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_111_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_111_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_111_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_112_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_112_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_112_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_112_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_112_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_113_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_113_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_113_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_113_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_113_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_114_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_114_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_114_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_114_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_114_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_115_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_115_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_115_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_115_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_115_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_116_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_116_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_116_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_116_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_116_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_117_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_117_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_117_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_117_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_117_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_118_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_118_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_118_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_118_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_118_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_119_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_119_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_119_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_119_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_119_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_120_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_120_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_120_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_120_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_120_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_121_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_121_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_121_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_121_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_121_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_122_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_122_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_122_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_122_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_122_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_123_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_123_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_123_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_123_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_123_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_124_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_124_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_124_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_124_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_124_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_125_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_125_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_125_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_125_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_125_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_126_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_126_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_126_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_126_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_126_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_127_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_127_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_127_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_127_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_127_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_128_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_128_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_128_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_128_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_128_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_129_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_129_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_129_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_129_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_129_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_130_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_130_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_130_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_130_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_130_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_131_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_131_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_131_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_131_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_131_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_132_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_132_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_132_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_132_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_132_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_133_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_133_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_133_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_133_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_133_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_134_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_134_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_134_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_134_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_134_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_135_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_135_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_135_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_135_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_135_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_136_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_136_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_136_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_136_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_136_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_137_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_137_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_137_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_137_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_137_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_138_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_138_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_138_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_138_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_138_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_139_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_139_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_139_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_139_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_139_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_140_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_140_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_140_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_140_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_140_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_141_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_141_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_141_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_141_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_141_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_142_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_142_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_142_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_142_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_142_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_143_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_143_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_143_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_143_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_143_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_144_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_144_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_144_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_144_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_144_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_145_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_145_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_145_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_145_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_145_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_146_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_146_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_146_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_146_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_146_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_147_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_147_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_147_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_147_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_147_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_148_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_148_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_148_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_148_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_148_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_149_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_149_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_149_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_149_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_149_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_150_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_150_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_150_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_150_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_150_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_151_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_151_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_151_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_151_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_151_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_152_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_152_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_152_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_152_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_152_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_153_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_153_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_153_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_153_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_153_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_154_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_154_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_154_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_154_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_154_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_155_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_155_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_155_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_155_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_155_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_156_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_156_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_156_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_156_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_156_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_157_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_157_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_157_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_157_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_157_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_158_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_158_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_158_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_158_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_158_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_159_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_159_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_159_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_159_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_159_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_160_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_160_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_160_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_160_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_160_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_161_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_161_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_161_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_161_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_161_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_162_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_162_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_162_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_162_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_162_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_163_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_163_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_163_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_163_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_163_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_164_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_164_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_164_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_164_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_164_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_7_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_7_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_7_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_7_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_165_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_165_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_165_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_165_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_165_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_166_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_166_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_166_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_166_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_166_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_167_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_167_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_167_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_167_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_167_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_168_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_168_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_168_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_168_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_168_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_169_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_169_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_169_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_169_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_169_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_170_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_170_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_170_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_170_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_170_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_171_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_171_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_171_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_171_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_171_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_172_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_172_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_172_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_172_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_172_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_173_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_173_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_173_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_173_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_173_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_174_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_174_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_174_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_174_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_174_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_175_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_175_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_175_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_175_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_175_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_176_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_176_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_176_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_176_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_176_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_177_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_177_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_177_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_177_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_177_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_178_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_178_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_178_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_178_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_178_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_179_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_179_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_179_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_179_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_179_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_180_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_180_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_180_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_180_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_180_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_181_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_181_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_181_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_181_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_181_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_182_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_182_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_182_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_182_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_182_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_183_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_183_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_183_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_183_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_183_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_184_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_184_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_184_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_184_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_184_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_185_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_185_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_185_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_185_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_185_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_186_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_186_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_186_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_186_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_186_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_187_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_187_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_187_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_187_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_187_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_188_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_188_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_188_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_188_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_188_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_189_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_189_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_189_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_189_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_189_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_190_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_190_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_190_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_190_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_190_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_191_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_191_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_191_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_191_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_191_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_192_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_192_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_192_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_192_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_192_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_193_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_193_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_193_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_193_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_193_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_194_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_194_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_194_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_194_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_194_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_195_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_195_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_195_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_195_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_195_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_196_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_196_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_196_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_196_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_196_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_197_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_197_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_197_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_197_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_197_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_8_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_8_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_8_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_8_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_198_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_198_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_198_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_198_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_198_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_199_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_199_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_199_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_199_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_199_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_200_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_200_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_200_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_200_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_200_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_201_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_201_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_201_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_201_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_201_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_202_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_202_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_202_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_202_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_202_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_203_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_203_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_203_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_203_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_203_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_204_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_204_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_204_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_204_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_204_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_205_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_205_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_205_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_205_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_205_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_206_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_206_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_206_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_206_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_206_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_207_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_207_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_207_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_207_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_207_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_208_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_208_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_208_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_208_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_208_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_209_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_209_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_209_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_209_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_209_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_210_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_210_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_210_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_210_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_210_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_211_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_211_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_211_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_211_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_211_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_212_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_212_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_212_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_212_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_212_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_213_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_213_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_213_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_213_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_213_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_214_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_214_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_214_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_214_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_214_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_215_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_215_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_215_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_215_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_215_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_216_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_216_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_216_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_216_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_216_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_217_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_217_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_217_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_217_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_217_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_218_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_218_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_218_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_218_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_218_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_219_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_219_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_219_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_219_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_219_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_220_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_220_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_220_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_220_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_220_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_221_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_221_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_221_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_221_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_221_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_222_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_222_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_222_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_222_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_222_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_223_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_223_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_223_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_223_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_223_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_224_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_224_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_224_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_224_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_224_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_225_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_225_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_225_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_225_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_225_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_226_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_226_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_226_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_226_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_226_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_227_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_227_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_227_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_227_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_227_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_228_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_228_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_228_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_228_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_228_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_229_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_229_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_229_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_229_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_229_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_230_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_230_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_230_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_230_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_230_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_231_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_231_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_231_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_231_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_231_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_232_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_232_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_232_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_232_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_232_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_233_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_233_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_233_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_233_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_233_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_9_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_9_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_9_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_9_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_234_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_234_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_234_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_234_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_234_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_235_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_235_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_235_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_235_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_235_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_236_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_236_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_236_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_236_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_236_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_237_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_237_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_237_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_237_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_237_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_238_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_238_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_238_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_238_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_238_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_239_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_239_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_239_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_239_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_239_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_240_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_240_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_240_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_240_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_240_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_241_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_241_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_241_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_241_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_241_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_242_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_242_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_242_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_242_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_242_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_243_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_243_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_243_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_243_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_243_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_244_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_244_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_244_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_244_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_244_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_245_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_245_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_245_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_245_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_245_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_246_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_246_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_246_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_246_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_246_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_247_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_247_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_247_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_247_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_247_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_248_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_248_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_248_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_248_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_248_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_249_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_249_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_249_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_249_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_249_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_250_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_250_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_250_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_250_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_250_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_251_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_251_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_251_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_251_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_251_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_252_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_252_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_252_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_252_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_252_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_253_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_253_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_253_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_253_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_253_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_254_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_254_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_254_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_254_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_254_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_255_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_255_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_255_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_255_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_255_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_256_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_256_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_256_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_256_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_256_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_257_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_257_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_257_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_257_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_257_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_258_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_258_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_258_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_258_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_258_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_259_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_259_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_259_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_259_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_259_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_260_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_260_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_260_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_260_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_260_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_261_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_261_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_261_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_261_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_261_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_262_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_262_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_262_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_262_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_262_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_263_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_263_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_263_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_263_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_263_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_264_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_264_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_264_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_264_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_264_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_265_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_265_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_265_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_265_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_265_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_266_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_266_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_266_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_266_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_266_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_267_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_267_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_267_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_267_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_267_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_268_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_268_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_268_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_268_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_268_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_269_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_269_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_269_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_269_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_269_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_270_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_270_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_270_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_270_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_270_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_271_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_271_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_271_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_271_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_271_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_272_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_272_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_272_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_272_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_272_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_10_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_10_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_10_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_10_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_273_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_273_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_273_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_273_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_273_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_274_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_274_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_274_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_274_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_274_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_275_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_275_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_275_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_275_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_275_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_276_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_276_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_276_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_276_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_276_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_277_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_277_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_277_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_277_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_277_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_278_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_278_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_278_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_278_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_278_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_279_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_279_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_279_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_279_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_279_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_280_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_280_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_280_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_280_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_280_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_281_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_281_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_281_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_281_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_281_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_282_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_282_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_282_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_282_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_282_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_283_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_283_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_283_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_283_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_283_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_284_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_284_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_284_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_284_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_284_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_285_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_285_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_285_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_285_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_285_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_286_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_286_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_286_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_286_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_286_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_287_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_287_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_287_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_287_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_287_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_288_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_288_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_288_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_288_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_288_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_289_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_289_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_289_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_289_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_289_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_290_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_290_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_290_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_290_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_290_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_291_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_291_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_291_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_291_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_291_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_292_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_292_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_292_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_292_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_292_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_293_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_293_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_293_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_293_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_293_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_294_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_294_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_294_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_294_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_294_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_295_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_295_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_295_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_295_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_295_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_296_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_296_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_296_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_296_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_296_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_297_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_297_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_297_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_297_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_297_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_298_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_298_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_298_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_298_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_298_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_299_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_299_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_299_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_299_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_299_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_300_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_300_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_300_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_300_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_300_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_301_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_301_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_301_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_301_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_301_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_302_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_302_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_302_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_302_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_302_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_303_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_303_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_303_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_303_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_303_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_304_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_304_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_304_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_304_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_304_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_305_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_305_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_305_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_305_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_305_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_306_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_306_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_306_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_306_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_306_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_307_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_307_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_307_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_307_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_307_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_308_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_308_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_308_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_308_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_308_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_309_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_309_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_309_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_309_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_309_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_310_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_310_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_310_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_310_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_310_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_311_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_311_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_311_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_311_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_311_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_312_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_312_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_312_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_312_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_312_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_313_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_313_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_313_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_313_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_313_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_314_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_314_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_314_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_314_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_314_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_11_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_11_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_11_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_11_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_315_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_315_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_315_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_315_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_315_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_316_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_316_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_316_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_316_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_316_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_317_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_317_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_317_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_317_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_317_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_318_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_318_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_318_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_318_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_318_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_319_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_319_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_319_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_319_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_319_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_320_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_320_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_320_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_320_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_320_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_321_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_321_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_321_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_321_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_321_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_322_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_322_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_322_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_322_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_322_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_323_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_323_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_323_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_323_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_323_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_324_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_324_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_324_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_324_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_324_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_325_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_325_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_325_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_325_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_325_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_326_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_326_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_326_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_326_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_326_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_327_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_327_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_327_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_327_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_327_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_328_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_328_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_328_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_328_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_328_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_329_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_329_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_329_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_329_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_329_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_330_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_330_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_330_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_330_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_330_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_331_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_331_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_331_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_331_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_331_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_332_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_332_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_332_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_332_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_332_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_333_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_333_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_333_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_333_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_333_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_334_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_334_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_334_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_334_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_334_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_335_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_335_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_335_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_335_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_335_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_336_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_336_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_336_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_336_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_336_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_337_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_337_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_337_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_337_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_337_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_338_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_338_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_338_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_338_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_338_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_339_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_339_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_339_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_339_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_339_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_340_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_340_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_340_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_340_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_340_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_341_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_341_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_341_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_341_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_341_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_342_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_342_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_342_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_342_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_342_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_343_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_343_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_343_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_343_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_343_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_344_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_344_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_344_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_344_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_344_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_345_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_345_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_345_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_345_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_345_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_346_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_346_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_346_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_346_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_346_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_347_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_347_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_347_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_347_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_347_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_348_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_348_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_348_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_348_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_348_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_349_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_349_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_349_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_349_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_349_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_350_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_350_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_350_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_350_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_350_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_351_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_351_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_351_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_351_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_351_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_352_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_352_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_352_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_352_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_352_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_353_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_353_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_353_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_353_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_353_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_354_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_354_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_354_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_354_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_354_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_355_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_355_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_355_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_355_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_355_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_356_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_356_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_356_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_356_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_356_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_357_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_357_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_357_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_357_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_357_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_358_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_358_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_358_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_358_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_358_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_359_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_359_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_359_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_359_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_359_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_12_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_12_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_12_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_12_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_360_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_360_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_360_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_360_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_360_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_361_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_361_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_361_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_361_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_361_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_362_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_362_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_362_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_362_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_362_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_363_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_363_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_363_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_363_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_363_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_364_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_364_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_364_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_364_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_364_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_365_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_365_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_365_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_365_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_365_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_366_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_366_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_366_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_366_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_366_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_367_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_367_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_367_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_367_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_367_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_368_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_368_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_368_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_368_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_368_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_369_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_369_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_369_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_369_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_369_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_370_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_370_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_370_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_370_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_370_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_371_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_371_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_371_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_371_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_371_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_372_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_372_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_372_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_372_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_372_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_373_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_373_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_373_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_373_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_373_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_374_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_374_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_374_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_374_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_374_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_375_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_375_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_375_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_375_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_375_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_376_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_376_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_376_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_376_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_376_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_377_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_377_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_377_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_377_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_377_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_378_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_378_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_378_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_378_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_378_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_379_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_379_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_379_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_379_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_379_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_380_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_380_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_380_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_380_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_380_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_381_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_381_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_381_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_381_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_381_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_382_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_382_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_382_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_382_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_382_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_383_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_383_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_383_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_383_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_383_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_384_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_384_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_384_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_384_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_384_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_385_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_385_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_385_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_385_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_385_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_386_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_386_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_386_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_386_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_386_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_387_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_387_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_387_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_387_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_387_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_388_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_388_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_388_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_388_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_388_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_389_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_389_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_389_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_389_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_389_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_390_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_390_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_390_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_390_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_390_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_391_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_391_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_391_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_391_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_391_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_392_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_392_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_392_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_392_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_392_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_393_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_393_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_393_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_393_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_393_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_394_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_394_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_394_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_394_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_394_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_395_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_395_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_395_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_395_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_395_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_396_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_396_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_396_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_396_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_396_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_397_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_397_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_397_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_397_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_397_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_398_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_398_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_398_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_398_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_398_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_399_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_399_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_399_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_399_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_399_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_400_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_400_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_400_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_400_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_400_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_401_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_401_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_401_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_401_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_401_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_402_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_402_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_402_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_402_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_402_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_403_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_403_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_403_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_403_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_403_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_404_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_404_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_404_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_404_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_404_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_405_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_405_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_405_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_405_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_405_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_406_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_406_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_406_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_406_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_406_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_407_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_407_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_407_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_407_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_407_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_13_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_13_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_13_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_13_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_408_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_408_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_408_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_408_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_408_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_409_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_409_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_409_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_409_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_409_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_410_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_410_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_410_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_410_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_410_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_411_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_411_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_411_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_411_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_411_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_412_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_412_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_412_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_412_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_412_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_413_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_413_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_413_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_413_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_413_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_414_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_414_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_414_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_414_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_414_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_415_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_415_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_415_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_415_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_415_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_416_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_416_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_416_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_416_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_416_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_417_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_417_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_417_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_417_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_417_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_418_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_418_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_418_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_418_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_418_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_419_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_419_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_419_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_419_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_419_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_420_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_420_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_420_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_420_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_420_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_421_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_421_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_421_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_421_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_421_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_422_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_422_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_422_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_422_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_422_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_423_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_423_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_423_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_423_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_423_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_424_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_424_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_424_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_424_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_424_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_425_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_425_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_425_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_425_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_425_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_426_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_426_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_426_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_426_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_426_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_427_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_427_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_427_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_427_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_427_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_428_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_428_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_428_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_428_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_428_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_429_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_429_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_429_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_429_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_429_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_430_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_430_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_430_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_430_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_430_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_431_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_431_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_431_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_431_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_431_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_432_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_432_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_432_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_432_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_432_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_433_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_433_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_433_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_433_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_433_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_434_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_434_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_434_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_434_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_434_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_435_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_435_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_435_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_435_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_435_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_436_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_436_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_436_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_436_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_436_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_437_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_437_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_437_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_437_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_437_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_438_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_438_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_438_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_438_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_438_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_439_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_439_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_439_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_439_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_439_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_440_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_440_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_440_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_440_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_440_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_441_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_441_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_441_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_441_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_441_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_442_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_442_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_442_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_442_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_442_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_443_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_443_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_443_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_443_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_443_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_444_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_444_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_444_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_444_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_444_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_445_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_445_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_445_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_445_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_445_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_446_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_446_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_446_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_446_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_446_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_447_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_447_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_447_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_447_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_447_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_448_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_448_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_448_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_448_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_448_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_449_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_449_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_449_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_449_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_449_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_450_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_450_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_450_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_450_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_450_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_451_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_451_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_451_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_451_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_451_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_452_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_452_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_452_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_452_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_452_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_453_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_453_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_453_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_453_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_453_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_454_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_454_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_454_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_454_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_454_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_455_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_455_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_455_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_455_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_455_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_456_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_456_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_456_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_456_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_456_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_457_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_457_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_457_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_457_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_457_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_458_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_458_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_458_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_458_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_458_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_14_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_14_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_14_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_14_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_459_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_459_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_459_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_459_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_459_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_460_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_460_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_460_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_460_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_460_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_461_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_461_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_461_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_461_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_461_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_462_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_462_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_462_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_462_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_462_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_463_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_463_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_463_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_463_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_463_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_464_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_464_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_464_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_464_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_464_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_465_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_465_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_465_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_465_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_465_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_466_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_466_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_466_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_466_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_466_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_467_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_467_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_467_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_467_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_467_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_468_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_468_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_468_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_468_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_468_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_469_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_469_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_469_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_469_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_469_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_470_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_470_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_470_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_470_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_470_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_471_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_471_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_471_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_471_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_471_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_472_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_472_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_472_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_472_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_472_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_473_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_473_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_473_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_473_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_473_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_474_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_474_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_474_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_474_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_474_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_475_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_475_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_475_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_475_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_475_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_476_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_476_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_476_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_476_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_476_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_477_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_477_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_477_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_477_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_477_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_478_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_478_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_478_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_478_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_478_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_479_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_479_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_479_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_479_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_479_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_480_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_480_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_480_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_480_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_480_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_481_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_481_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_481_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_481_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_481_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_482_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_482_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_482_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_482_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_482_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_483_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_483_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_483_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_483_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_483_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_484_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_484_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_484_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_484_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_484_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_485_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_485_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_485_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_485_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_485_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_486_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_486_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_486_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_486_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_486_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_487_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_487_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_487_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_487_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_487_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_488_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_488_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_488_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_488_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_488_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_489_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_489_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_489_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_489_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_489_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_490_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_490_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_490_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_490_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_490_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_491_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_491_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_491_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_491_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_491_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_492_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_492_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_492_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_492_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_492_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_493_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_493_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_493_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_493_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_493_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_494_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_494_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_494_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_494_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_494_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_495_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_495_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_495_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_495_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_495_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_496_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_496_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_496_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_496_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_496_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_497_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_497_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_497_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_497_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_497_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_498_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_498_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_498_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_498_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_498_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_499_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_499_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_499_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_499_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_499_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_500_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_500_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_500_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_500_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_500_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_501_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_501_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_501_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_501_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_501_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_502_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_502_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_502_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_502_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_502_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_503_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_503_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_503_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_503_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_503_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_504_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_504_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_504_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_504_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_504_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_505_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_505_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_505_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_505_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_505_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_506_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_506_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_506_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_506_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_506_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_507_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_507_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_507_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_507_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_507_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_508_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_508_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_508_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_508_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_508_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_509_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_509_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_509_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_509_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_509_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_510_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_510_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_510_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_510_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_510_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_511_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_511_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_511_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_511_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_511_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_512_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_512_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_512_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_512_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_512_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_15_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_15_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_15_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_15_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_513_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_513_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_513_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_513_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_513_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_514_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_514_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_514_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_514_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_514_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_515_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_515_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_515_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_515_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_515_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_516_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_516_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_516_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_516_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_516_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_517_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_517_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_517_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_517_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_517_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_518_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_518_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_518_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_518_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_518_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_519_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_519_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_519_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_519_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_519_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_520_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_520_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_520_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_520_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_520_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_521_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_521_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_521_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_521_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_521_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_522_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_522_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_522_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_522_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_522_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_523_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_523_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_523_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_523_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_523_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_524_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_524_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_524_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_524_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_524_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_525_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_525_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_525_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_525_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_525_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_526_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_526_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_526_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_526_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_526_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_527_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_527_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_527_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_527_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_527_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_528_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_528_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_528_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_528_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_528_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_529_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_529_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_529_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_529_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_529_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_530_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_530_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_530_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_530_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_530_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_531_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_531_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_531_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_531_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_531_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_532_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_532_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_532_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_532_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_532_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_533_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_533_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_533_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_533_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_533_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_534_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_534_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_534_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_534_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_534_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_535_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_535_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_535_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_535_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_535_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_536_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_536_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_536_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_536_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_536_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_537_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_537_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_537_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_537_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_537_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_538_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_538_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_538_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_538_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_538_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_539_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_539_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_539_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_539_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_539_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_540_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_540_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_540_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_540_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_540_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_541_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_541_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_541_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_541_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_541_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_542_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_542_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_542_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_542_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_542_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_543_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_543_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_543_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_543_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_543_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_544_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_544_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_544_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_544_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_544_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_545_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_545_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_545_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_545_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_545_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_546_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_546_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_546_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_546_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_546_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_547_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_547_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_547_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_547_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_547_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_548_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_548_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_548_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_548_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_548_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_549_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_549_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_549_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_549_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_549_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_550_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_550_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_550_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_550_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_550_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_551_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_551_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_551_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_551_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_551_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_552_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_552_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_552_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_552_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_552_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_553_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_553_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_553_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_553_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_553_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_554_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_554_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_554_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_554_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_554_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_555_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_555_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_555_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_555_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_555_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_556_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_556_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_556_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_556_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_556_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_557_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_557_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_557_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_557_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_557_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_558_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_558_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_558_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_558_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_558_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_559_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_559_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_559_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_559_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_559_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_560_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_560_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_560_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_560_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_560_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_561_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_561_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_561_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_561_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_561_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_562_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_562_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_562_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_562_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_562_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_563_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_563_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_563_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_563_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_563_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_564_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_564_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_564_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_564_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_564_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_565_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_565_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_565_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_565_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_565_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_566_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_566_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_566_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_566_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_566_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_567_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_567_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_567_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_567_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_567_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_568_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_568_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_568_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_568_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_568_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_569_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_569_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_569_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_569_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_569_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_16_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_16_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_16_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_16_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_570_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_570_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_570_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_570_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_570_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_571_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_571_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_571_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_571_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_571_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_572_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_572_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_572_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_572_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_572_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_573_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_573_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_573_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_573_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_573_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_574_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_574_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_574_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_574_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_574_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_575_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_575_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_575_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_575_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_575_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_576_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_576_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_576_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_576_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_576_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_577_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_577_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_577_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_577_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_577_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_578_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_578_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_578_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_578_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_578_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_579_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_579_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_579_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_579_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_579_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_580_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_580_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_580_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_580_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_580_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_581_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_581_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_581_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_581_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_581_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_582_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_582_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_582_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_582_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_582_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_583_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_583_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_583_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_583_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_583_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_584_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_584_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_584_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_584_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_584_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_585_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_585_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_585_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_585_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_585_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_586_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_586_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_586_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_586_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_586_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_587_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_587_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_587_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_587_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_587_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_588_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_588_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_588_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_588_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_588_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_589_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_589_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_589_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_589_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_589_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_590_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_590_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_590_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_590_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_590_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_591_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_591_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_591_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_591_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_591_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_592_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_592_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_592_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_592_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_592_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_593_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_593_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_593_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_593_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_593_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_594_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_594_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_594_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_594_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_594_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_595_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_595_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_595_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_595_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_595_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_596_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_596_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_596_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_596_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_596_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_597_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_597_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_597_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_597_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_597_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_598_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_598_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_598_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_598_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_598_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_599_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_599_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_599_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_599_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_599_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_600_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_600_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_600_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_600_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_600_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_601_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_601_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_601_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_601_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_601_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_602_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_602_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_602_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_602_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_602_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_603_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_603_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_603_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_603_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_603_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_604_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_604_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_604_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_604_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_604_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_605_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_605_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_605_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_605_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_605_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_606_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_606_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_606_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_606_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_606_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_607_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_607_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_607_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_607_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_607_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_608_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_608_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_608_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_608_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_608_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_609_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_609_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_609_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_609_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_609_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_610_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_610_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_610_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_610_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_610_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_611_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_611_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_611_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_611_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_611_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_612_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_612_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_612_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_612_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_612_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_613_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_613_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_613_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_613_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_613_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_614_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_614_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_614_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_614_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_614_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_615_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_615_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_615_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_615_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_615_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_616_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_616_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_616_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_616_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_616_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_617_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_617_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_617_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_617_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_617_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_618_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_618_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_618_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_618_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_618_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_619_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_619_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_619_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_619_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_619_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_620_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_620_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_620_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_620_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_620_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_621_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_621_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_621_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_621_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_621_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_622_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_622_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_622_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_622_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_622_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_623_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_623_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_623_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_623_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_623_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_624_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_624_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_624_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_624_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_624_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_625_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_625_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_625_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_625_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_625_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_626_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_626_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_626_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_626_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_626_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_627_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_627_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_627_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_627_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_627_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_628_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_628_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_628_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_628_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_628_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_629_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_629_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_629_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_629_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_629_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_17_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_17_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_17_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_17_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_630_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_630_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_630_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_630_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_630_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_631_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_631_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_631_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_631_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_631_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_632_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_632_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_632_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_632_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_632_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_633_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_633_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_633_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_633_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_633_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_634_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_634_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_634_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_634_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_634_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_635_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_635_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_635_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_635_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_635_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_636_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_636_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_636_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_636_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_636_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_637_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_637_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_637_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_637_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_637_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_638_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_638_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_638_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_638_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_638_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_639_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_639_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_639_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_639_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_639_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_640_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_640_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_640_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_640_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_640_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_641_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_641_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_641_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_641_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_641_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_642_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_642_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_642_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_642_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_642_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_643_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_643_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_643_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_643_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_643_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_644_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_644_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_644_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_644_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_644_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_645_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_645_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_645_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_645_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_645_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_646_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_646_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_646_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_646_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_646_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_647_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_647_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_647_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_647_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_647_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_648_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_648_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_648_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_648_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_648_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_649_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_649_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_649_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_649_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_649_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_650_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_650_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_650_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_650_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_650_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_651_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_651_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_651_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_651_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_651_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_652_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_652_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_652_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_652_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_652_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_653_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_653_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_653_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_653_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_653_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_654_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_654_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_654_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_654_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_654_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_655_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_655_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_655_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_655_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_655_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_656_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_656_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_656_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_656_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_656_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_657_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_657_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_657_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_657_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_657_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_658_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_658_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_658_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_658_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_658_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_659_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_659_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_659_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_659_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_659_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_660_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_660_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_660_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_660_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_660_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_661_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_661_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_661_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_661_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_661_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_662_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_662_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_662_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_662_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_662_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_663_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_663_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_663_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_663_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_663_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_664_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_664_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_664_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_664_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_664_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_665_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_665_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_665_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_665_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_665_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_666_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_666_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_666_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_666_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_666_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_667_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_667_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_667_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_667_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_667_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_668_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_668_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_668_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_668_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_668_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_669_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_669_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_669_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_669_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_669_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_670_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_670_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_670_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_670_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_670_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_671_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_671_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_671_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_671_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_671_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_672_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_672_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_672_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_672_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_672_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_673_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_673_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_673_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_673_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_673_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_674_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_674_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_674_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_674_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_674_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_675_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_675_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_675_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_675_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_675_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_676_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_676_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_676_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_676_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_676_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_677_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_677_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_677_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_677_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_677_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_678_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_678_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_678_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_678_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_678_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_679_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_679_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_679_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_679_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_679_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_680_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_680_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_680_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_680_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_680_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_681_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_681_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_681_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_681_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_681_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_682_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_682_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_682_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_682_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_682_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_683_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_683_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_683_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_683_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_683_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_684_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_684_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_684_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_684_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_684_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_685_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_685_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_685_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_685_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_685_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_686_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_686_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_686_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_686_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_686_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_687_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_687_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_687_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_687_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_687_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_688_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_688_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_688_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_688_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_688_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_689_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_689_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_689_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_689_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_689_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_690_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_690_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_690_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_690_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_690_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_691_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_691_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_691_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_691_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_691_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_692_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_692_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_692_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_692_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_692_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_693_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_693_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_693_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_693_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_693_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_694_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_694_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_694_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_694_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_694_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_695_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_695_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_695_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_695_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_695_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_696_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_696_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_696_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_696_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_696_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_697_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_697_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_697_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_697_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_697_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_698_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_698_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_698_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_698_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_698_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_699_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_699_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_699_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_699_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_699_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_700_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_700_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_700_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_700_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_700_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_701_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_701_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_701_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_701_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_701_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_702_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_702_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_702_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_702_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_702_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_703_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_703_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_703_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_703_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_703_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_704_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_704_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_704_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_704_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_704_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_705_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_705_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_705_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_705_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_705_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_706_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_706_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_706_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_706_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_706_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_707_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_707_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_707_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_707_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_707_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_708_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_708_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_708_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_708_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_708_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_709_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_709_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_709_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_709_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_709_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_710_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_710_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_710_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_710_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_710_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_711_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_711_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_711_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_711_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_711_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_712_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_712_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_712_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_712_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_712_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_18_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_18_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_18_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_18_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_713_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_713_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_713_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_713_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_713_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_714_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_714_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_714_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_714_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_714_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_715_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_715_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_715_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_715_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_715_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_716_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_716_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_716_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_716_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_716_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_717_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_717_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_717_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_717_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_717_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_718_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_718_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_718_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_718_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_718_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_719_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_719_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_719_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_719_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_719_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_720_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_720_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_720_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_720_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_720_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_721_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_721_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_721_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_721_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_721_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_722_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_722_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_722_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_722_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_722_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_723_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_723_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_723_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_723_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_723_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_724_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_724_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_724_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_724_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_724_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_725_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_725_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_725_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_725_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_725_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_726_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_726_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_726_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_726_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_726_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_727_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_727_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_727_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_727_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_727_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_728_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_728_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_728_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_728_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_728_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_729_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_729_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_729_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_729_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_729_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_730_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_730_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_730_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_730_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_730_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_731_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_731_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_731_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_731_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_731_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_732_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_732_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_732_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_732_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_732_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_733_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_733_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_733_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_733_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_733_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_734_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_734_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_734_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_734_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_734_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_735_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_735_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_735_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_735_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_735_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_736_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_736_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_736_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_736_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_736_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_737_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_737_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_737_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_737_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_737_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_738_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_738_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_738_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_738_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_738_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_739_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_739_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_739_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_739_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_739_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_740_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_740_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_740_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_740_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_740_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_741_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_741_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_741_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_741_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_741_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_742_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_742_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_742_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_742_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_742_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_743_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_743_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_743_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_743_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_743_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_744_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_744_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_744_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_744_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_744_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_745_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_745_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_745_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_745_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_745_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_746_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_746_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_746_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_746_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_746_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_747_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_747_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_747_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_747_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_747_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_748_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_748_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_748_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_748_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_748_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_749_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_749_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_749_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_749_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_749_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_750_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_750_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_750_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_750_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_750_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_751_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_751_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_751_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_751_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_751_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_752_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_752_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_752_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_752_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_752_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_753_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_753_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_753_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_753_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_753_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_754_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_754_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_754_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_754_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_754_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_755_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_755_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_755_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_755_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_755_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_756_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_756_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_756_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_756_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_756_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_757_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_757_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_757_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_757_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_757_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_758_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_758_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_758_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_758_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_758_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_759_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_759_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_759_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_759_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_759_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_760_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_760_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_760_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_760_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_760_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_761_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_761_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_761_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_761_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_761_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_762_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_762_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_762_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_762_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_762_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_763_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_763_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_763_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_763_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_763_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_764_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_764_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_764_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_764_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_764_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_765_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_765_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_765_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_765_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_765_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_766_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_766_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_766_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_766_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_766_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_767_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_767_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_767_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_767_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_767_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_768_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_768_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_768_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_768_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_768_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_769_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_769_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_769_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_769_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_769_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_770_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_770_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_770_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_770_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_770_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_771_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_771_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_771_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_771_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_771_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_19_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_19_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_19_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_19_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_772_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_772_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_772_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_772_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_772_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_773_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_773_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_773_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_773_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_773_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_774_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_774_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_774_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_774_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_774_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_775_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_775_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_775_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_775_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_775_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_776_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_776_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_776_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_776_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_776_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_777_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_777_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_777_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_777_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_777_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_778_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_778_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_778_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_778_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_778_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_779_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_779_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_779_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_779_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_779_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_780_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_780_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_780_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_780_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_780_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_781_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_781_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_781_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_781_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_781_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_782_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_782_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_782_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_782_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_782_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_783_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_783_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_783_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_783_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_783_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_784_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_784_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_784_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_784_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_784_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_785_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_785_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_785_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_785_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_785_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_786_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_786_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_786_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_786_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_786_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_787_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_787_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_787_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_787_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_787_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_788_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_788_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_788_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_788_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_788_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_789_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_789_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_789_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_789_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_789_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_790_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_790_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_790_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_790_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_790_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_791_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_791_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_791_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_791_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_791_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_792_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_792_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_792_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_792_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_792_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_793_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_793_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_793_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_793_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_793_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_794_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_794_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_794_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_794_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_794_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_795_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_795_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_795_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_795_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_795_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_796_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_796_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_796_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_796_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_796_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_797_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_797_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_797_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_797_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_797_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_798_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_798_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_798_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_798_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_798_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_799_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_799_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_799_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_799_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_799_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_800_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_800_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_800_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_800_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_800_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_801_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_801_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_801_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_801_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_801_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_802_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_802_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_802_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_802_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_802_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_803_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_803_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_803_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_803_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_803_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_804_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_804_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_804_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_804_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_804_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_805_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_805_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_805_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_805_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_805_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_806_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_806_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_806_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_806_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_806_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_807_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_807_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_807_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_807_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_807_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_808_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_808_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_808_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_808_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_808_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_809_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_809_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_809_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_809_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_809_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_810_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_810_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_810_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_810_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_810_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_811_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_811_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_811_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_811_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_811_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_812_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_812_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_812_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_812_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_812_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_813_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_813_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_813_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_813_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_813_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_814_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_814_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_814_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_814_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_814_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_815_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_815_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_815_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_815_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_815_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_816_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_816_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_816_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_816_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_816_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_817_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_817_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_817_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_817_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_817_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_818_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_818_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_818_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_818_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_818_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_819_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_819_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_819_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_819_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_819_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_820_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_820_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_820_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_820_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_820_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_821_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_821_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_821_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_821_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_821_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_822_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_822_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_822_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_822_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_822_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_823_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_823_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_823_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_823_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_823_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_824_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_824_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_824_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_824_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_824_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_825_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_825_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_825_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_825_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_825_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_826_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_826_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_826_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_826_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_826_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_827_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_827_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_827_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_827_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_827_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_828_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_828_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_828_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_828_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_828_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_829_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_829_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_829_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_829_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_829_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_830_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_830_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_830_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_830_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_830_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_831_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_831_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_831_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_831_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_831_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_832_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_832_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_832_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_832_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_832_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_833_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_833_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_833_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_833_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_833_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_834_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_834_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_834_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_834_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_834_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_835_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_835_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_835_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_835_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_835_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_836_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_836_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_836_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_836_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_836_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_837_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_837_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_837_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_837_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_837_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_838_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_838_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_838_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_838_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_838_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_839_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_839_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_839_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_839_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_839_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_840_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_840_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_840_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_840_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_840_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_841_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_841_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_841_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_841_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_841_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_842_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_842_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_842_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_842_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_842_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_843_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_843_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_843_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_843_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_843_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_844_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_844_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_844_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_844_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_844_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_845_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_845_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_845_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_845_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_845_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_846_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_846_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_846_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_846_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_846_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_847_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_847_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_847_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_847_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_847_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_848_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_848_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_848_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_848_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_848_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_849_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_849_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_849_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_849_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_849_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_850_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_850_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_850_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_850_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_850_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_851_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_851_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_851_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_851_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_851_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_852_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_852_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_852_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_852_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_852_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_853_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_853_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_853_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_853_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_853_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_854_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_854_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_854_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_854_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_854_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_855_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_855_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_855_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_855_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_855_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_856_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_856_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_856_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_856_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_856_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_857_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_857_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_857_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_857_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_857_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_858_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_858_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_858_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_858_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_858_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_859_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_859_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_859_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_859_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_859_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_860_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_860_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_860_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_860_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_860_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_861_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_861_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_861_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_861_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_861_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_862_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_862_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_862_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_862_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_862_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_863_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_863_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_863_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_863_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_863_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_864_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_864_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_864_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_864_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_864_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_865_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_865_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_865_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_865_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_865_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_866_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_866_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_866_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_866_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_866_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_867_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_867_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_867_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_867_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_867_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_868_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_868_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_868_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_868_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_868_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_869_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_869_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_869_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_869_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_869_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_870_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_870_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_870_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_870_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_870_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_871_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_871_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_871_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_871_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_871_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_872_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_872_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_872_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_872_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_872_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_873_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_873_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_873_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_873_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_873_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_874_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_874_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_874_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_874_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_874_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_875_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_875_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_875_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_875_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_875_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_876_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_876_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_876_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_876_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_876_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_877_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_877_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_877_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_877_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_877_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_878_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_878_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_878_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_878_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_878_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_879_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_879_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_879_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_879_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_879_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_880_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_880_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_880_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_880_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_880_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_20_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_20_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_20_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_20_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_881_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_881_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_881_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_881_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_881_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_882_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_882_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_882_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_882_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_882_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_883_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_883_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_883_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_883_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_883_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_884_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_884_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_884_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_884_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_884_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_885_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_885_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_885_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_885_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_885_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_886_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_886_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_886_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_886_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_886_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_887_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_887_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_887_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_887_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_887_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_888_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_888_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_888_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_888_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_888_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_889_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_889_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_889_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_889_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_889_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_890_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_890_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_890_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_890_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_890_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_891_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_891_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_891_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_891_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_891_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_892_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_892_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_892_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_892_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_892_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_893_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_893_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_893_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_893_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_893_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_894_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_894_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_894_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_894_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_894_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_895_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_895_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_895_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_895_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_895_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_896_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_896_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_896_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_896_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_896_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_897_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_897_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_897_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_897_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_897_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_898_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_898_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_898_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_898_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_898_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_899_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_899_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_899_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_899_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_899_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_900_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_900_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_900_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_900_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_900_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_901_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_901_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_901_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_901_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_901_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_902_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_902_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_902_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_902_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_902_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_903_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_903_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_903_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_903_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_903_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_904_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_904_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_904_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_904_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_904_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_905_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_905_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_905_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_905_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_905_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_906_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_906_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_906_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_906_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_906_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_907_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_907_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_907_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_907_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_907_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_908_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_908_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_908_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_908_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_908_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_909_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_909_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_909_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_909_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_909_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_910_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_910_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_910_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_910_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_910_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_911_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_911_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_911_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_911_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_911_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_912_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_912_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_912_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_912_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_912_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_913_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_913_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_913_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_913_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_913_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_914_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_914_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_914_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_914_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_914_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_915_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_915_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_915_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_915_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_915_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_916_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_916_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_916_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_916_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_916_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_917_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_917_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_917_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_917_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_917_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_918_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_918_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_918_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_918_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_918_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_919_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_919_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_919_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_919_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_919_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_920_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_920_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_920_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_920_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_920_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_921_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_921_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_921_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_921_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_921_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_922_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_922_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_922_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_922_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_922_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_923_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_923_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_923_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_923_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_923_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_924_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_924_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_924_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_924_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_924_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_925_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_925_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_925_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_925_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_925_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_926_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_926_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_926_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_926_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_926_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_927_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_927_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_927_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_927_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_927_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_928_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_928_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_928_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_928_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_928_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_929_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_929_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_929_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_929_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_929_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_930_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_930_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_930_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_930_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_930_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_931_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_931_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_931_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_931_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_931_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_932_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_932_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_932_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_932_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_932_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_933_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_933_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_933_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_933_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_933_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_934_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_934_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_934_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_934_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_934_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_935_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_935_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_935_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_935_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_935_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_936_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_936_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_936_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_936_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_936_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_937_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_937_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_937_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_937_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_937_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_938_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_938_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_938_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_938_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_938_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_939_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_939_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_939_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_939_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_939_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_940_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_940_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_940_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_940_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_940_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_941_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_941_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_941_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_941_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_941_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_942_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_942_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_942_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_942_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_942_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_943_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_943_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_943_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_943_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_943_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_944_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_944_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_944_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_944_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_944_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_945_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_945_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_945_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_945_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_945_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_946_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_946_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_946_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_946_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_946_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_947_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_947_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_947_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_947_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_947_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_948_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_948_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_948_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_948_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_948_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_949_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_949_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_949_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_949_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_949_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_950_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_950_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_950_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_950_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_950_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_951_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_951_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_951_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_951_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_951_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_952_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_952_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_952_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_952_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_952_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_953_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_953_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_953_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_953_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_953_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_954_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_954_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_954_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_954_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_954_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_955_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_955_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_955_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_955_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_955_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_956_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_956_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_956_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_956_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_956_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_957_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_957_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_957_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_957_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_957_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_958_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_958_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_958_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_958_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_958_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_959_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_959_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_959_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_959_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_959_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_960_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_960_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_960_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_960_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_960_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_961_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_961_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_961_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_961_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_961_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_962_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_962_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_962_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_962_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_962_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_963_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_963_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_963_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_963_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_963_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_964_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_964_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_964_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_964_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_964_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_965_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_965_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_965_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_965_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_965_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_966_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_966_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_966_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_966_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_966_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_967_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_967_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_967_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_967_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_967_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_968_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_968_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_968_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_968_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_968_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_969_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_969_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_969_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_969_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_969_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_970_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_970_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_970_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_970_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_970_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_971_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_971_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_971_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_971_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_971_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_972_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_972_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_972_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_972_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_972_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_973_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_973_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_973_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_973_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_973_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_974_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_974_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_974_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_974_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_974_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_975_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_975_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_975_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_975_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_975_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_976_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_976_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_976_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_976_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_976_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_977_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_977_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_977_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_977_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_977_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_21_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_21_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_21_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_21_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_978_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_978_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_978_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_978_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_978_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_979_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_979_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_979_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_979_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_979_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_980_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_980_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_980_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_980_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_980_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_981_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_981_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_981_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_981_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_981_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_982_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_982_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_982_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_982_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_982_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_983_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_983_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_983_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_983_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_983_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_984_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_984_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_984_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_984_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_984_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_985_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_985_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_985_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_985_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_985_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_986_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_986_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_986_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_986_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_986_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_987_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_987_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_987_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_987_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_987_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_988_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_988_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_988_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_988_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_988_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_989_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_989_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_989_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_989_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_989_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_990_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_990_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_990_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_990_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_990_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_991_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_991_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_991_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_991_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_991_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_992_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_992_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_992_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_992_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_992_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_993_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_993_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_993_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_993_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_993_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_994_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_994_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_994_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_994_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_994_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_995_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_995_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_995_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_995_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_995_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_996_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_996_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_996_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_996_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_996_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_997_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_997_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_997_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_997_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_997_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_998_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_998_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_998_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_998_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_998_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_999_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_999_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_999_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_999_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_999_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1000_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1000_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1000_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1000_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1000_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1001_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1001_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1001_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1001_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1001_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1002_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1002_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1002_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1002_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1002_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1003_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1003_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1003_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1003_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1003_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1004_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1004_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1004_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1004_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1004_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1005_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1005_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1005_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1005_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1005_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1006_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1006_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1006_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1006_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1006_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1007_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1007_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1007_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1007_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1007_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1008_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1008_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1008_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1008_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1008_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1009_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1009_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1009_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1009_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1009_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1010_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1010_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1010_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1010_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1010_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1011_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1011_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1011_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1011_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1011_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1012_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1012_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1012_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1012_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1012_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1013_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1013_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1013_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1013_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1013_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1014_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1014_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1014_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1014_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1014_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1015_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1015_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1015_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1015_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1015_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1016_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1016_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1016_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1016_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1016_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1017_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1017_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1017_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1017_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1017_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1018_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1018_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1018_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1018_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1018_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1019_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1019_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1019_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1019_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1019_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1020_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1020_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1020_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1020_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1020_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1021_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1021_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1021_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1021_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1021_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1022_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1022_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1022_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1022_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1022_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1023_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1023_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1023_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1023_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1023_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1024_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1024_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1024_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1024_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1024_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1025_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1025_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1025_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1025_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1025_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1026_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1026_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1026_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1026_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1026_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1027_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1027_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1027_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1027_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1027_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1028_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1028_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1028_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1028_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1028_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1029_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1029_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1029_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1029_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1029_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1030_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1030_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1030_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1030_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1030_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1031_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1031_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1031_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1031_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1031_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1032_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1032_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1032_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1032_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1032_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1033_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1033_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1033_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1033_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1033_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1034_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1034_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1034_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1034_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1034_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1035_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1035_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1035_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1035_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1035_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1036_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1036_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1036_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1036_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1036_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1037_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1037_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1037_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1037_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1037_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1038_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1038_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1038_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1038_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1038_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1039_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1039_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1039_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1039_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1039_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1040_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1040_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1040_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1040_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1040_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1041_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1041_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1041_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1041_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1041_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1042_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1042_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1042_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1042_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1042_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1043_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1043_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1043_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1043_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1043_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1044_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1044_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1044_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1044_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1044_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1045_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1045_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1045_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1045_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1045_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1046_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1046_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1046_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1046_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1046_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1047_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1047_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1047_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1047_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1047_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1048_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1048_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1048_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1048_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1048_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1049_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1049_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1049_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1049_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1049_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1050_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1050_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1050_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1050_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1050_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1051_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1051_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1051_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1051_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1051_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1052_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1052_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1052_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1052_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1052_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1053_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1053_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1053_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1053_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1053_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1054_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1054_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1054_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1054_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1054_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1055_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1055_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1055_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1055_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1055_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1056_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1056_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1056_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1056_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1056_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1057_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1057_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1057_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1057_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1057_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1058_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1058_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1058_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1058_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1058_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1059_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1059_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1059_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1059_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1059_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1060_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1060_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1060_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1060_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1060_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1061_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1061_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1061_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1061_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1061_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1062_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1062_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1062_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1062_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1062_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1063_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1063_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1063_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1063_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1063_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1064_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1064_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1064_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1064_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1064_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1065_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1065_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1065_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1065_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1065_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1066_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1066_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1066_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1066_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1066_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1067_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1067_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1067_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1067_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1067_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1068_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1068_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1068_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1068_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1068_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1069_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1069_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1069_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1069_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1069_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1070_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1070_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1070_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1070_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1070_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1071_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1071_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1071_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1071_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1071_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1072_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1072_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1072_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1072_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1072_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1073_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1073_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1073_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1073_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1073_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1074_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1074_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1074_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1074_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1074_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1075_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1075_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1075_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1075_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1075_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1076_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1076_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1076_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1076_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1076_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1077_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1077_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1077_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1077_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1077_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1078_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1078_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1078_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1078_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1078_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1079_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1079_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1079_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1079_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1079_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1080_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1080_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1080_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1080_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1080_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1081_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1081_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1081_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1081_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1081_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1082_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1082_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1082_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1082_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1082_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1083_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1083_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1083_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1083_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1083_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1084_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1084_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1084_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1084_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1084_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1085_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1085_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1085_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1085_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1085_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1086_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1086_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1086_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1086_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1086_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1087_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1087_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1087_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1087_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1087_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1088_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1088_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1088_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1088_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1088_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1089_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1089_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1089_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1089_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1089_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1090_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1090_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1090_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1090_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1090_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1091_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1091_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1091_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1091_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1091_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1092_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1092_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1092_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1092_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1092_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1093_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1093_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1093_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1093_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1093_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1094_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1094_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1094_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1094_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1094_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1095_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1095_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1095_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1095_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1095_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1096_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1096_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1096_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1096_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1096_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1097_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1097_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1097_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1097_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1097_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1098_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1098_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1098_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1098_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1098_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1099_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1099_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1099_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1099_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1099_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1100_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1100_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1100_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1100_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1100_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_22_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_22_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_22_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_22_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1101_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1101_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1101_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1101_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1101_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1102_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1102_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1102_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1102_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1102_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1103_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1103_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1103_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1103_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1103_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1104_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1104_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1104_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1104_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1104_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1105_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1105_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1105_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1105_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1105_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1106_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1106_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1106_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1106_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1106_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1107_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1107_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1107_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1107_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1107_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1108_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1108_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1108_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1108_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1108_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1109_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1109_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1109_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1109_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1109_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1110_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1110_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1110_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1110_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1110_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1111_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1111_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1111_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1111_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1111_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1112_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1112_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1112_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1112_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1112_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1113_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1113_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1113_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1113_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1113_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1114_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1114_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1114_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1114_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1114_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1115_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1115_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1115_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1115_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1115_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1116_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1116_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1116_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1116_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1116_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1117_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1117_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1117_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1117_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1117_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1118_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1118_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1118_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1118_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1118_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1119_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1119_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1119_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1119_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1119_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1120_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1120_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1120_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1120_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1120_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1121_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1121_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1121_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1121_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1121_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1122_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1122_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1122_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1122_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1122_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1123_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1123_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1123_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1123_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1123_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1124_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1124_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1124_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1124_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1124_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1125_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1125_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1125_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1125_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1125_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1126_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1126_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1126_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1126_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1126_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1127_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1127_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1127_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1127_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1127_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1128_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1128_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1128_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1128_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1128_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1129_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1129_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1129_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1129_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1129_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1130_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1130_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1130_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1130_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1130_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1131_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1131_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1131_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1131_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1131_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1132_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1132_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1132_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1132_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1132_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1133_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1133_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1133_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1133_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1133_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1134_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1134_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1134_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1134_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1134_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1135_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1135_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1135_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1135_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1135_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_23_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_23_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_23_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_23_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1136_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1136_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1136_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1136_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1136_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1137_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1137_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1137_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1137_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1137_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1138_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1138_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1138_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1138_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1138_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1139_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1139_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1139_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1139_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1139_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1140_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1140_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1140_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1140_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1140_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1141_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1141_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1141_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1141_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1141_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1142_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1142_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1142_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1142_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1142_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1143_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1143_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1143_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1143_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1143_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1144_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1144_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1144_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1144_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1144_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1145_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1145_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1145_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1145_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1145_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1146_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1146_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1146_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1146_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1146_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1147_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1147_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1147_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1147_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1147_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1148_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1148_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1148_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1148_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1148_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1149_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1149_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1149_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1149_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1149_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1150_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1150_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1150_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1150_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1150_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1151_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1151_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1151_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1151_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1151_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1152_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1152_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1152_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1152_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1152_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1153_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1153_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1153_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1153_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1153_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1154_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1154_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1154_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1154_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1154_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1155_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1155_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1155_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1155_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1155_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1156_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1156_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1156_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1156_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1156_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1157_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1157_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1157_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1157_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1157_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1158_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1158_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1158_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1158_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1158_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1159_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1159_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1159_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1159_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1159_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1160_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1160_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1160_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1160_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1160_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1161_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1161_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1161_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1161_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1161_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1162_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1162_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1162_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1162_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1162_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1163_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1163_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1163_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1163_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1163_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1164_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1164_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1164_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1164_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1164_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1165_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1165_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1165_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1165_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1165_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1166_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1166_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1166_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1166_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1166_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1167_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1167_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1167_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1167_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1167_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_24_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_24_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_24_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_24_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1168_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1168_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1168_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1168_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1168_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1169_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1169_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1169_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1169_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1169_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1170_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1170_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1170_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1170_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1170_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1171_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1171_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1171_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1171_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1171_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1172_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1172_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1172_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1172_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1172_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1173_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1173_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1173_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1173_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1173_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1174_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1174_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1174_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1174_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1174_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1175_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1175_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1175_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1175_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1175_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1176_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1176_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1176_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1176_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1176_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1177_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1177_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1177_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1177_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1177_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1178_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1178_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1178_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1178_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1178_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1179_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1179_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1179_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1179_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1179_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1180_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1180_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1180_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1180_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1180_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1181_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1181_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1181_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1181_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1181_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1182_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1182_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1182_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1182_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1182_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1183_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1183_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1183_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1183_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1183_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1184_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1184_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1184_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1184_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1184_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1185_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1185_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1185_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1185_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1185_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1186_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1186_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1186_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1186_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1186_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1187_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1187_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1187_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1187_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1187_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1188_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1188_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1188_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1188_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1188_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1189_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1189_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1189_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1189_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1189_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1190_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1190_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1190_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1190_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1190_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1191_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1191_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1191_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1191_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1191_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1192_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1192_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1192_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1192_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1192_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1193_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1193_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1193_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1193_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1193_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1194_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1194_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1194_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1194_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1194_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1195_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1195_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1195_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1195_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1195_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1196_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1196_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1196_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1196_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1196_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_25_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_25_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_25_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_25_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1197_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1197_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1197_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1197_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1197_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1198_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1198_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1198_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1198_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1198_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1199_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1199_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1199_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1199_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1199_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1200_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1200_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1200_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1200_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1200_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1201_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1201_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1201_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1201_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1201_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1202_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1202_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1202_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1202_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1202_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1203_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1203_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1203_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1203_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1203_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1204_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1204_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1204_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1204_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1204_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1205_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1205_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1205_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1205_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1205_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1206_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1206_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1206_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1206_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1206_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1207_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1207_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1207_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1207_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1207_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1208_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1208_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1208_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1208_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1208_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1209_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1209_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1209_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1209_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1209_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1210_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1210_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1210_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1210_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1210_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1211_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1211_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1211_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1211_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1211_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1212_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1212_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1212_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1212_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1212_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1213_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1213_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1213_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1213_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1213_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1214_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1214_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1214_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1214_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1214_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1215_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1215_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1215_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1215_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1215_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1216_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1216_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1216_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1216_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1216_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1217_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1217_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1217_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1217_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1217_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1218_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1218_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1218_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1218_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1218_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1219_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1219_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1219_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1219_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1219_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1220_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1220_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1220_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1220_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1220_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1221_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1221_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1221_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1221_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1221_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1222_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1222_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1222_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1222_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1222_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1223_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1223_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1223_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1223_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1223_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1224_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1224_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1224_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1224_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1224_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1225_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1225_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1225_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1225_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1225_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1226_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1226_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1226_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1226_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1226_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1227_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1227_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1227_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1227_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1227_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1228_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1228_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1228_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1228_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1228_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1229_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1229_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1229_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1229_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1229_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1230_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1230_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1230_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1230_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1230_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1231_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1231_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1231_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1231_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1231_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1232_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1232_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1232_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1232_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1232_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1233_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1233_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1233_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1233_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1233_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1234_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1234_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1234_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1234_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1234_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1235_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1235_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1235_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1235_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1235_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1236_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1236_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1236_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1236_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1236_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1237_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1237_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1237_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1237_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1237_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1238_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1238_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1238_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1238_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1238_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1239_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1239_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1239_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1239_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1239_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1240_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1240_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1240_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1240_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1240_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1241_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1241_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1241_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1241_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1241_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1242_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1242_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1242_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1242_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1242_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1243_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1243_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1243_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1243_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1243_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1244_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1244_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1244_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1244_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1244_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1245_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1245_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1245_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1245_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1245_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_26_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_26_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_26_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_26_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1246_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1246_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1246_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1246_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1246_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1247_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1247_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1247_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1247_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1247_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1248_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1248_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1248_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1248_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1248_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1249_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1249_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1249_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1249_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1249_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1250_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1250_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1250_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1250_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1250_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1251_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1251_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1251_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1251_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1251_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1252_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1252_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1252_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1252_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1252_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1253_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1253_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1253_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1253_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1253_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1254_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1254_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1254_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1254_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1254_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1255_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1255_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1255_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1255_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1255_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1256_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1256_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1256_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1256_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1256_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1257_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1257_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1257_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1257_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1257_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1258_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1258_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1258_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1258_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1258_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1259_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1259_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1259_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1259_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1259_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1260_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1260_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1260_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1260_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1260_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1261_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1261_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1261_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1261_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1261_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1262_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1262_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1262_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1262_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1262_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1263_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1263_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1263_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1263_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1263_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1264_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1264_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1264_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1264_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1264_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1265_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1265_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1265_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1265_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1265_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_27_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_27_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_27_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_27_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1266_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1266_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1266_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1266_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1266_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1267_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1267_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1267_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1267_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1267_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1268_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1268_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1268_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1268_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1268_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1269_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1269_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1269_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1269_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1269_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1270_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1270_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1270_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1270_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1270_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1271_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1271_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1271_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1271_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1271_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1272_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1272_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1272_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1272_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1272_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1273_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1273_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1273_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1273_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1273_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1274_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1274_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1274_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1274_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1274_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1275_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1275_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1275_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1275_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1275_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1276_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1276_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1276_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1276_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1276_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1277_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1277_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1277_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1277_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1277_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1278_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1278_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1278_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1278_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1278_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1279_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1279_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1279_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1279_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1279_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1280_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1280_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1280_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1280_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1280_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1281_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1281_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1281_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1281_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1281_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1282_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1282_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1282_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1282_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1282_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_28_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_28_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_28_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_28_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1283_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1283_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1283_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1283_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1283_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1284_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1284_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1284_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1284_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1284_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1285_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1285_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1285_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1285_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1285_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1286_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1286_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1286_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1286_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1286_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1287_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1287_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1287_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1287_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1287_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1288_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1288_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1288_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1288_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1288_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1289_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1289_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1289_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1289_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1289_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1290_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1290_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1290_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1290_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1290_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1291_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1291_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1291_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1291_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1291_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1292_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1292_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1292_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1292_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1292_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1293_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1293_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1293_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1293_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1293_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1294_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1294_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1294_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1294_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1294_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1295_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1295_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1295_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1295_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1295_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1296_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1296_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1296_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1296_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1296_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_29_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_29_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_29_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_29_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1297_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1297_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1297_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1297_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1297_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1298_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1298_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1298_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1298_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1298_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1299_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1299_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1299_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1299_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1299_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1300_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1300_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1300_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1300_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1300_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1301_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1301_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1301_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1301_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1301_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1302_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1302_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1302_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1302_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1302_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1303_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1303_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1303_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1303_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1303_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1304_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1304_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1304_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1304_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1304_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1305_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1305_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1305_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1305_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1305_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1306_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1306_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1306_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1306_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1306_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1307_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1307_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1307_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1307_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1307_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_30_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_30_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_30_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_30_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1308_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1308_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1308_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1308_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1308_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1309_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1309_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1309_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1309_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1309_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1310_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1310_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1310_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1310_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1310_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1311_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1311_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1311_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1311_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1311_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1312_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1312_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1312_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1312_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1312_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1313_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1313_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1313_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1313_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1313_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1314_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1314_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1314_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1314_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1314_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1315_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1315_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1315_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1315_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1315_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_31_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_31_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_31_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_31_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1316_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1316_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1316_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1316_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1316_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1317_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1317_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1317_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1317_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1317_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1318_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1318_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1318_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1318_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1318_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1319_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1319_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1319_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1319_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1319_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1320_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1320_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1320_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1320_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1320_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_32_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_32_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_32_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_32_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1321_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1321_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1321_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1321_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1321_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_33_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_33_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_33_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_33_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_34_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_34_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_34_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_34_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_35_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_35_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_35_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_35_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_36_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_36_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_36_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_36_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1322_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1322_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1322_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1322_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1322_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1323_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1323_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1323_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1323_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1323_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1324_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1324_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1324_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1324_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1324_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1325_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1325_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1325_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1325_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1325_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1326_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1326_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1326_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1326_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1326_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1327_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1327_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1327_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1327_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1327_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1328_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1328_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1328_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1328_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1328_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1329_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1329_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1329_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1329_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1329_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1330_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1330_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1330_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1330_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1330_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1331_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1331_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1331_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1331_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1331_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1332_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1332_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1332_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1332_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1332_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1333_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1333_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1333_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1333_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1333_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1334_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1334_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1334_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1334_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1334_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_37_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_37_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_37_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_37_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1335_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1335_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1335_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1335_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1335_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1336_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1336_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1336_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1336_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1336_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_38_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_38_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_38_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_38_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1337_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1337_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1337_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1337_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1337_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1338_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1338_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1338_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1338_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1338_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1339_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1339_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1339_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1339_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1339_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1340_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1340_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1340_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1340_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1340_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1341_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1341_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1341_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1341_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1341_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1342_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1342_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1342_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1342_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1342_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1343_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1343_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1343_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1343_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1343_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1344_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1344_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1344_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1344_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1344_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1345_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1345_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1345_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1345_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1345_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1346_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1346_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1346_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1346_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1346_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1347_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1347_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1347_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1347_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1347_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1348_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1348_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1348_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1348_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1348_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1349_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1349_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1349_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1349_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1349_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1350_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1350_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1350_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1350_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1350_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1351_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1351_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1351_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1351_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1351_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1352_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1352_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1352_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1352_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1352_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1353_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1353_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1353_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1353_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1353_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1354_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1354_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1354_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1354_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1354_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1355_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1355_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1355_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1355_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1355_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1356_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1356_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1356_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1356_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1356_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1357_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1357_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1357_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1357_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1357_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1358_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1358_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1358_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1358_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1358_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1359_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1359_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1359_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1359_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1359_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1360_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1360_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1360_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1360_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1360_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1361_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1361_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1361_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1361_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1361_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_39_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_39_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_39_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_39_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1362_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1362_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1362_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1362_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1362_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1363_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1363_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1363_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1363_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1363_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1364_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1364_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1364_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1364_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1364_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1365_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1365_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1365_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1365_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1365_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_40_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_40_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_40_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_40_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1366_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1366_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1366_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1366_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1366_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1367_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1367_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1367_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1367_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1367_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1368_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1368_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1368_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1368_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1368_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1369_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1369_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1369_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1369_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1369_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_41_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_41_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_41_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_41_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1370_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1370_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1370_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1370_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1370_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1371_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1371_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1371_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1371_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1371_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1372_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1372_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1372_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1372_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1372_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1373_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1373_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1373_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1373_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1373_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1374_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1374_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1374_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1374_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1374_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1375_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1375_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1375_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1375_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1375_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1376_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1376_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1376_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1376_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1376_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1377_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1377_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1377_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1377_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1377_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1378_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1378_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1378_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1378_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1378_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1379_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1379_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1379_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1379_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1379_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1380_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1380_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1380_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1380_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1380_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1381_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1381_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1381_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1381_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1381_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1382_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1382_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1382_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1382_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1382_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1383_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1383_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1383_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1383_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1383_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1384_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1384_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1384_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1384_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1384_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1385_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1385_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1385_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1385_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1385_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1386_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1386_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1386_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1386_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1386_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1387_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1387_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1387_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1387_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1387_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1388_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1388_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1388_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1388_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1388_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1389_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1389_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1389_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1389_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1389_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1390_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1390_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1390_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1390_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1390_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1391_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1391_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1391_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1391_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1391_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1392_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1392_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1392_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1392_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1392_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1393_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1393_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1393_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1393_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1393_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1394_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1394_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1394_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1394_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1394_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1395_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1395_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1395_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1395_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1395_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1396_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1396_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1396_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1396_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1396_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1397_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1397_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1397_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1397_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1397_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1398_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1398_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1398_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1398_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1398_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1399_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1399_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1399_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1399_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1399_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1400_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1400_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1400_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1400_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1400_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1401_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1401_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1401_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1401_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1401_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1402_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1402_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1402_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1402_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1402_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1403_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1403_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1403_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1403_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1403_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1404_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1404_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1404_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1404_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1404_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1405_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1405_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1405_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1405_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1405_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1406_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1406_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1406_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1406_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1406_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1407_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1407_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1407_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1407_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1407_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1408_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1408_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1408_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1408_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1408_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1409_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1409_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1409_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1409_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1409_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1410_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1410_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1410_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1410_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1410_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1411_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1411_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1411_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1411_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1411_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1412_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1412_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1412_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1412_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1412_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1413_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1413_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1413_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1413_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1413_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1414_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1414_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1414_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1414_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1414_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1415_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1415_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1415_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1415_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1415_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1416_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1416_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1416_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1416_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1416_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1417_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1417_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1417_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1417_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1417_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1418_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1418_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1418_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1418_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1418_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1419_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1419_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1419_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1419_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1419_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1420_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1420_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1420_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1420_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1420_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_42_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_42_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_42_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_42_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1421_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1421_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1421_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1421_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1421_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1422_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1422_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1422_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1422_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1422_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1423_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1423_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1423_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1423_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1423_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1424_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1424_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1424_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1424_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1424_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1425_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1425_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1425_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1425_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1425_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1426_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1426_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1426_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1426_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1426_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1427_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1427_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1427_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1427_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1427_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1428_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1428_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1428_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1428_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1428_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1429_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1429_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1429_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1429_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1429_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1430_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1430_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1430_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1430_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1430_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1431_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1431_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1431_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1431_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1431_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1432_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1432_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1432_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1432_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1432_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1433_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1433_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1433_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1433_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1433_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1434_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1434_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1434_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1434_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1434_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1435_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1435_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1435_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1435_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1435_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1436_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1436_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1436_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1436_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1436_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1437_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1437_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1437_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1437_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1437_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1438_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1438_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1438_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1438_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1438_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1439_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1439_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1439_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1439_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1439_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1440_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1440_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1440_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1440_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1440_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1441_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1441_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1441_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1441_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1441_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1442_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1442_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1442_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1442_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1442_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1443_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1443_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1443_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1443_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1443_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1444_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1444_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1444_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1444_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1444_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1445_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1445_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1445_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1445_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1445_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1446_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1446_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1446_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1446_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1446_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1447_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1447_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1447_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1447_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1447_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1448_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1448_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1448_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1448_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1448_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1449_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1449_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1449_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1449_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1449_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1450_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1450_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1450_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1450_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1450_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1451_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1451_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1451_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1451_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1451_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1452_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1452_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1452_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1452_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1452_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1453_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1453_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1453_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1453_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1453_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1454_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1454_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1454_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1454_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1454_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1455_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1455_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1455_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1455_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1455_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1456_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1456_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1456_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1456_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1456_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1457_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1457_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1457_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1457_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1457_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1458_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1458_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1458_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1458_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1458_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1459_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1459_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1459_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1459_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1459_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1460_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1460_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1460_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1460_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1460_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1461_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1461_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1461_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1461_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1461_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1462_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1462_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1462_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1462_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1462_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1463_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1463_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1463_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1463_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1463_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1464_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1464_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1464_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1464_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1464_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1465_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1465_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1465_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1465_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1465_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1466_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1466_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1466_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1466_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1466_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1467_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1467_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1467_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1467_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1467_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1468_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1468_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1468_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1468_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1468_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1469_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1469_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1469_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1469_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1469_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1470_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1470_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1470_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1470_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1470_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1471_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1471_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1471_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1471_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1471_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1472_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1472_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1472_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1472_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1472_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1473_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1473_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1473_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1473_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1473_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_43_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_43_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_43_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_43_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1474_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1474_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1474_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1474_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1474_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1475_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1475_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1475_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1475_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1475_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1476_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1476_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1476_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1476_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1476_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1477_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1477_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1477_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1477_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1477_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1478_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1478_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1478_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1478_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1478_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1479_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1479_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1479_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1479_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1479_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1480_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1480_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1480_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1480_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1480_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1481_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1481_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1481_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1481_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1481_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_44_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_44_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_44_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_44_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1482_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1482_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1482_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1482_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1482_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1483_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1483_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1483_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1483_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1483_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1484_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1484_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1484_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1484_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1484_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1485_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1485_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1485_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1485_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1485_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1486_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1486_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1486_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1486_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1486_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1487_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1487_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1487_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1487_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1487_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1488_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1488_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1488_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1488_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1488_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1489_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1489_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1489_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1489_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1489_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_45_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_45_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_45_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_45_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1490_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1490_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1490_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1490_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1490_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1491_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1491_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1491_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1491_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1491_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1492_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1492_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1492_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1492_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1492_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1493_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1493_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1493_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1493_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1493_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1494_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1494_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1494_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1494_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1494_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1495_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1495_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1495_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1495_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1495_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1496_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1496_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1496_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1496_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1496_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1497_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1497_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1497_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1497_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1497_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1498_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1498_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1498_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1498_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1498_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1499_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1499_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1499_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1499_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1499_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1500_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1500_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1500_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1500_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1500_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1501_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1501_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1501_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1501_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1501_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1502_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1502_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1502_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1502_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1502_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1503_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1503_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1503_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1503_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1503_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1504_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1504_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1504_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1504_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1504_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1505_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1505_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1505_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1505_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1505_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1506_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1506_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1506_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1506_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1506_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1507_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1507_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1507_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1507_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1507_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1508_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1508_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1508_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1508_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1508_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1509_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1509_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1509_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1509_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1509_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1510_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1510_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1510_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1510_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1510_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1511_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1511_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1511_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1511_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1511_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1512_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1512_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1512_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1512_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1512_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1513_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1513_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1513_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1513_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1513_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1514_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1514_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1514_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1514_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1514_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1515_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1515_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1515_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1515_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1515_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1516_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1516_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1516_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1516_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1516_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1517_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1517_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1517_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1517_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1517_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1518_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1518_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1518_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1518_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1518_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1519_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1519_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1519_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1519_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1519_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1520_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1520_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1520_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1520_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1520_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1521_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1521_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1521_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1521_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1521_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1522_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1522_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1522_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1522_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1522_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1523_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1523_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1523_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1523_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1523_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1524_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1524_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1524_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1524_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1524_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1525_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1525_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1525_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1525_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1525_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1526_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1526_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1526_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1526_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1526_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1527_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1527_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1527_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1527_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1527_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1528_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1528_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1528_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1528_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1528_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1529_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1529_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1529_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1529_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1529_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1530_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1530_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1530_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1530_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1530_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1531_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1531_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1531_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1531_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1531_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1532_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1532_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1532_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1532_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1532_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1533_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1533_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1533_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1533_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1533_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1534_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1534_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1534_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1534_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1534_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1535_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1535_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1535_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1535_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1535_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1536_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1536_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1536_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1536_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1536_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1537_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1537_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1537_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1537_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1537_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1538_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1538_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1538_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1538_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1538_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1539_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1539_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1539_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1539_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1539_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1540_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1540_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1540_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1540_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1540_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1541_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1541_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1541_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1541_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1541_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1542_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1542_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1542_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1542_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1542_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1543_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1543_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1543_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1543_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1543_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1544_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1544_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1544_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1544_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1544_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1545_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1545_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1545_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1545_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1545_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1546_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1546_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1546_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1546_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1546_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1547_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1547_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1547_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1547_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1547_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1548_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1548_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1548_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1548_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1548_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1549_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1549_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1549_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1549_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1549_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1550_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1550_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1550_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1550_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1550_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1551_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1551_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1551_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1551_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1551_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1552_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1552_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1552_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1552_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1552_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1553_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1553_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1553_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1553_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1553_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1554_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1554_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1554_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1554_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1554_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1555_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1555_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1555_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1555_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1555_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1556_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1556_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1556_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1556_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1556_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1557_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1557_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1557_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1557_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1557_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1558_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1558_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1558_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1558_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1558_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1559_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1559_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1559_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1559_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1559_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1560_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1560_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1560_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1560_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1560_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1561_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1561_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1561_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1561_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1561_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1562_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1562_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1562_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1562_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1562_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1563_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1563_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1563_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1563_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1563_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1564_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1564_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1564_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1564_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1564_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1565_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1565_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1565_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1565_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1565_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1566_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1566_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1566_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1566_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1566_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1567_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1567_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1567_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1567_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1567_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1568_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1568_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1568_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1568_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1568_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1569_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1569_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1569_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1569_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1569_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1570_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1570_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1570_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1570_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1570_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1571_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1571_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1571_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1571_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1571_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1572_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1572_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1572_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1572_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1572_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1573_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1573_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1573_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1573_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1573_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1574_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1574_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1574_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1574_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1574_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1575_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1575_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1575_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1575_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1575_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1576_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1576_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1576_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1576_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1576_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_46_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_46_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_46_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_46_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1577_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1577_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1577_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1577_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1577_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1578_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1578_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1578_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1578_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1578_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1579_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1579_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1579_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1579_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1579_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1580_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1580_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1580_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1580_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1580_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1581_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1581_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1581_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1581_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1581_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1582_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1582_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1582_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1582_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1582_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1583_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1583_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1583_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1583_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1583_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1584_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1584_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1584_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1584_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1584_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1585_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1585_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1585_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1585_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1585_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1586_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1586_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1586_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1586_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1586_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1587_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1587_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1587_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1587_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1587_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1588_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1588_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1588_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1588_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1588_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1589_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1589_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1589_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1589_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1589_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1590_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1590_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1590_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1590_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1590_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1591_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1591_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1591_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1591_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1591_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1592_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1592_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1592_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1592_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1592_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1593_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1593_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1593_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1593_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1593_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1594_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1594_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1594_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1594_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1594_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1595_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1595_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1595_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1595_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1595_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1596_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1596_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1596_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1596_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1596_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1597_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1597_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1597_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1597_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1597_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1598_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1598_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1598_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1598_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1598_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1599_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1599_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1599_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1599_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1599_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1600_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1600_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1600_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1600_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1600_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1601_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1601_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1601_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1601_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1601_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1602_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1602_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1602_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1602_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1602_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1603_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1603_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1603_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1603_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1603_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1604_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1604_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1604_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1604_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1604_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1605_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1605_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1605_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1605_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1605_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1606_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1606_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1606_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1606_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1606_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1607_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1607_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1607_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1607_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1607_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1608_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1608_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1608_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1608_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1608_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1609_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1609_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1609_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1609_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1609_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1610_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1610_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1610_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1610_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1610_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1611_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1611_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1611_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1611_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1611_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1612_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1612_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1612_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1612_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1612_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1613_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1613_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1613_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1613_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1613_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1614_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1614_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1614_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1614_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1614_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1615_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1615_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1615_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1615_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1615_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1616_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1616_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1616_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1616_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1616_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1617_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1617_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1617_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1617_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1617_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1618_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1618_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1618_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1618_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1618_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1619_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1619_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1619_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1619_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1619_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1620_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1620_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1620_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1620_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1620_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1621_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1621_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1621_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1621_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1621_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1622_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1622_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1622_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1622_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1622_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1623_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1623_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1623_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1623_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1623_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1624_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1624_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1624_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1624_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1624_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1625_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1625_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1625_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1625_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1625_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1626_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1626_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1626_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1626_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1626_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1627_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1627_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1627_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1627_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1627_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1628_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1628_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1628_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1628_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1628_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1629_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1629_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1629_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1629_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1629_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1630_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1630_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1630_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1630_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1630_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1631_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1631_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1631_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1631_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1631_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1632_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1632_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1632_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1632_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1632_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1633_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1633_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1633_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1633_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1633_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1634_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1634_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1634_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1634_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1634_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1635_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1635_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1635_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1635_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1635_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1636_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1636_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1636_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1636_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1636_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1637_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1637_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1637_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1637_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1637_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1638_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1638_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1638_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1638_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1638_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1639_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1639_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1639_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1639_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1639_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1640_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1640_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1640_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1640_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1640_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1641_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1641_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1641_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1641_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1641_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1642_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1642_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1642_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1642_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1642_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1643_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1643_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1643_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1643_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1643_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1644_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1644_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1644_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1644_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1644_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1645_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1645_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1645_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1645_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1645_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1646_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1646_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1646_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1646_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1646_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1647_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1647_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1647_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1647_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1647_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1648_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1648_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1648_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1648_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1648_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1649_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1649_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1649_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1649_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1649_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1650_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1650_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1650_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1650_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1650_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1651_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1651_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1651_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1651_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1651_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1652_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1652_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1652_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1652_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1652_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1653_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1653_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1653_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1653_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1653_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1654_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1654_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1654_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1654_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1654_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1655_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1655_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1655_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1655_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1655_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1656_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1656_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1656_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1656_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1656_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1657_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1657_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1657_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1657_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1657_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_47_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_47_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_47_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_47_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1658_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1658_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1658_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1658_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1658_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1659_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1659_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1659_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1659_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1659_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1660_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1660_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1660_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1660_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1660_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1661_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1661_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1661_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1661_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1661_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1662_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1662_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1662_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1662_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1662_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1663_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1663_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1663_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1663_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1663_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1664_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1664_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1664_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1664_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1664_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1665_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1665_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1665_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1665_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1665_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1666_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1666_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1666_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1666_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1666_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1667_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1667_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1667_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1667_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1667_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1668_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1668_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1668_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1668_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1668_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1669_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1669_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1669_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1669_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1669_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_48_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_48_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_48_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_48_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1670_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1670_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1670_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1670_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1670_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1671_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1671_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1671_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1671_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1671_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1672_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1672_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1672_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1672_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1672_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1673_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1673_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1673_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1673_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1673_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1674_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1674_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1674_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1674_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1674_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1675_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1675_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1675_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1675_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1675_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1676_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1676_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1676_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1676_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1676_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1677_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1677_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1677_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1677_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1677_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1678_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1678_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1678_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1678_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1678_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1679_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1679_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1679_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1679_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1679_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1680_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1680_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1680_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1680_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1680_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1681_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1681_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1681_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1681_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1681_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1682_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1682_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1682_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1682_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1682_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1683_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1683_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1683_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1683_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1683_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1684_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1684_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1684_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1684_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1684_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1685_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1685_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1685_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1685_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1685_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1686_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1686_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1686_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1686_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1686_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1687_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1687_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1687_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1687_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1687_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1688_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1688_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1688_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1688_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1688_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1689_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1689_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1689_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1689_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1689_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1690_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1690_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1690_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1690_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1690_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1691_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1691_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1691_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1691_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1691_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1692_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1692_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1692_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1692_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1692_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1693_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1693_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1693_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1693_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1693_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1694_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1694_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1694_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1694_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1694_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1695_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1695_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1695_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1695_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1695_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1696_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1696_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1696_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1696_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1696_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1697_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1697_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1697_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1697_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1697_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1698_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1698_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1698_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1698_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1698_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1699_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1699_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1699_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1699_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1699_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1700_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1700_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1700_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1700_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1700_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1701_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1701_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1701_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1701_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1701_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1702_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1702_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1702_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1702_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1702_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1703_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1703_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1703_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1703_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1703_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1704_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1704_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1704_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1704_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1704_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1705_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1705_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1705_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1705_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1705_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1706_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1706_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1706_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1706_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1706_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1707_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1707_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1707_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1707_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1707_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1708_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1708_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1708_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1708_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1708_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1709_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1709_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1709_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1709_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1709_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1710_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1710_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1710_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1710_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1710_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1711_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1711_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1711_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1711_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1711_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1712_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1712_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1712_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1712_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1712_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1713_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1713_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1713_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1713_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1713_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1714_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1714_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1714_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1714_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1714_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1715_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1715_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1715_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1715_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1715_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1716_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1716_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1716_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1716_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1716_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1717_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1717_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1717_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1717_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1717_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1718_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1718_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1718_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1718_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1718_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1719_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1719_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1719_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1719_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1719_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1720_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1720_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1720_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1720_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1720_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1721_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1721_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1721_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1721_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1721_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1722_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1722_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1722_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1722_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1722_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1723_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1723_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1723_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1723_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1723_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1724_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1724_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1724_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1724_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1724_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1725_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1725_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1725_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1725_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1725_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1726_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1726_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1726_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1726_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1726_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1727_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1727_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1727_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1727_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1727_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1728_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1728_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1728_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1728_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1728_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1729_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1729_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1729_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1729_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1729_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1730_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1730_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1730_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1730_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1730_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1731_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1731_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1731_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1731_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1731_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1732_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1732_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1732_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1732_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1732_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1733_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1733_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1733_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1733_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1733_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1734_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1734_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1734_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1734_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1734_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1735_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1735_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1735_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1735_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1735_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1736_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1736_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1736_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1736_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1736_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1737_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1737_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1737_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1737_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1737_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1738_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1738_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1738_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1738_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1738_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1739_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1739_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1739_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1739_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1739_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1740_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1740_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1740_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1740_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1740_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1741_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1741_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1741_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1741_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1741_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1742_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1742_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1742_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1742_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1742_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1743_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1743_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1743_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1743_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1743_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1744_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1744_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1744_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1744_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1744_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1745_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1745_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1745_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1745_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1745_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1746_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1746_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1746_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1746_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1746_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1747_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1747_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1747_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1747_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1747_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1748_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1748_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1748_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1748_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1748_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1749_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1749_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1749_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1749_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1749_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1750_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1750_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1750_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1750_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1750_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1751_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1751_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1751_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1751_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1751_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1752_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1752_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1752_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1752_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1752_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1753_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1753_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1753_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1753_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1753_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1754_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1754_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1754_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1754_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1754_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1755_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1755_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1755_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1755_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1755_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1756_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1756_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1756_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1756_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1756_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1757_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1757_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1757_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1757_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1757_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1758_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1758_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1758_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1758_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1758_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1759_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1759_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1759_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1759_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1759_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1760_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1760_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1760_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1760_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1760_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1761_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1761_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1761_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1761_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1761_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1762_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1762_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1762_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1762_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1762_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1763_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1763_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1763_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1763_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1763_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1764_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1764_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1764_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1764_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1764_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1765_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1765_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1765_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1765_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1765_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1766_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1766_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1766_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1766_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1766_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1767_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1767_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1767_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1767_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1767_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1768_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1768_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1768_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1768_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1768_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1769_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1769_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1769_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1769_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1769_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1770_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1770_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1770_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1770_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1770_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1771_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1771_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1771_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1771_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1771_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1772_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1772_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1772_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1772_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1772_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1773_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1773_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1773_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1773_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1773_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1774_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1774_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1774_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1774_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1774_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1775_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1775_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1775_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1775_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1775_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1776_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1776_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1776_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1776_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1776_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1777_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1777_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1777_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1777_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1777_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1778_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1778_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1778_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1778_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1778_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1779_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1779_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1779_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1779_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1779_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1780_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1780_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1780_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1780_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1780_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1781_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1781_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1781_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1781_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1781_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1782_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1782_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1782_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1782_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1782_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1783_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1783_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1783_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1783_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1783_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1784_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1784_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1784_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1784_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1784_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1785_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1785_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1785_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1785_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1785_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1786_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1786_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1786_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1786_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1786_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1787_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1787_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1787_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1787_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1787_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1788_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1788_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1788_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1788_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1788_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1789_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1789_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1789_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1789_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1789_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1790_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1790_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1790_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1790_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1790_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1791_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1791_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1791_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1791_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1791_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1792_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1792_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1792_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1792_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1792_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1793_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1793_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1793_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1793_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1793_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1794_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1794_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1794_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1794_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1794_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1795_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1795_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1795_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1795_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1795_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1796_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1796_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1796_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1796_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1796_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1797_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1797_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1797_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1797_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1797_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1798_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1798_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1798_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1798_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1798_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1799_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1799_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1799_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1799_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1799_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1800_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1800_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1800_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1800_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1800_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1801_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1801_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1801_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1801_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1801_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1802_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1802_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1802_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1802_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1802_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1803_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1803_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1803_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1803_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1803_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_49_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_49_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_49_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_49_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1804_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1804_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1804_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1804_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1804_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1805_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1805_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1805_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1805_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1805_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1806_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1806_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1806_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1806_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1806_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1807_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1807_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1807_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1807_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1807_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1808_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1808_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1808_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1808_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1808_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1809_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1809_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1809_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1809_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1809_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1810_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1810_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1810_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1810_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1810_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1811_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1811_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1811_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1811_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1811_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1812_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1812_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1812_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1812_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1812_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1813_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1813_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1813_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1813_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1813_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1814_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1814_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1814_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1814_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1814_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1815_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1815_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1815_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1815_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1815_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1816_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1816_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1816_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1816_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1816_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1817_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1817_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1817_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1817_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1817_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1818_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1818_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1818_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1818_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1818_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1819_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1819_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1819_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1819_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1819_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1820_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1820_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1820_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1820_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1820_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1821_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1821_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1821_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1821_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1821_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1822_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1822_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1822_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1822_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1822_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1823_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1823_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1823_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1823_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1823_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1824_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1824_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1824_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1824_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1824_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1825_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1825_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1825_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1825_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1825_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1826_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1826_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1826_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1826_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1826_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1827_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1827_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1827_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1827_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1827_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1828_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1828_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1828_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1828_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1828_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1829_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1829_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1829_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1829_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1829_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1830_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1830_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1830_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1830_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1830_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1831_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1831_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1831_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1831_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1831_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1832_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1832_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1832_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1832_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1832_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1833_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1833_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1833_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1833_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1833_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1834_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1834_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1834_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1834_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1834_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1835_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1835_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1835_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1835_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1835_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1836_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1836_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1836_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1836_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1836_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1837_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1837_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1837_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1837_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1837_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1838_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1838_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1838_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1838_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1838_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1839_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1839_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1839_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1839_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1839_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1840_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1840_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1840_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1840_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1840_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1841_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1841_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1841_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1841_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1841_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1842_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1842_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1842_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1842_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1842_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1843_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1843_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1843_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1843_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1843_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1844_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1844_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1844_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1844_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1844_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1845_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1845_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1845_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1845_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1845_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1846_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1846_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1846_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1846_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1846_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1847_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1847_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1847_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1847_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1847_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1848_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1848_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1848_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1848_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1848_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1849_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1849_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1849_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1849_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1849_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1850_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1850_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1850_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1850_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1850_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1851_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1851_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1851_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1851_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1851_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1852_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1852_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1852_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1852_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1852_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1853_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1853_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1853_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1853_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1853_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1854_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1854_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1854_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1854_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1854_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1855_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1855_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1855_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1855_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1855_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1856_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1856_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1856_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1856_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1856_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1857_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1857_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1857_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1857_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1857_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1858_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1858_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1858_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1858_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1858_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1859_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1859_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1859_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1859_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1859_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1860_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1860_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1860_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1860_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1860_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1861_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1861_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1861_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1861_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1861_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1862_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1862_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1862_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1862_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1862_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1863_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1863_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1863_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1863_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1863_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1864_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1864_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1864_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1864_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1864_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1865_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1865_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1865_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1865_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1865_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1866_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1866_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1866_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1866_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1866_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1867_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1867_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1867_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1867_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1867_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1868_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1868_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1868_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1868_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1868_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1869_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1869_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1869_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1869_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1869_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1870_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1870_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1870_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1870_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1870_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1871_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1871_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1871_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1871_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1871_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1872_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1872_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1872_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1872_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1872_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1873_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1873_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1873_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1873_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1873_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1874_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1874_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1874_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1874_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1874_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1875_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1875_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1875_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1875_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1875_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1876_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1876_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1876_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1876_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1876_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1877_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1877_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1877_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1877_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1877_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1878_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1878_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1878_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1878_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1878_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1879_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1879_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1879_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1879_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1879_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1880_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1880_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1880_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1880_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1880_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1881_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1881_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1881_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1881_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1881_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1882_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1882_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1882_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1882_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1882_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1883_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1883_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1883_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1883_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1883_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1884_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1884_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1884_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1884_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1884_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1885_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1885_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1885_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1885_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1885_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1886_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1886_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1886_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1886_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1886_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1887_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1887_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1887_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1887_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1887_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1888_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1888_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1888_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1888_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1888_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1889_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1889_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1889_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1889_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1889_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1890_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1890_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1890_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1890_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1890_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1891_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1891_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1891_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1891_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1891_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1892_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1892_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1892_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1892_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1892_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1893_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1893_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1893_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1893_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1893_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1894_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1894_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1894_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1894_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1894_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1895_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1895_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1895_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1895_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1895_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1896_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1896_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1896_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1896_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1896_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1897_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1897_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1897_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1897_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1897_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1898_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1898_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1898_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1898_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1898_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1899_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1899_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1899_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1899_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1899_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1900_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1900_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1900_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1900_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1900_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1901_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1901_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1901_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1901_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1901_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1902_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1902_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1902_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1902_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1902_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1903_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1903_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1903_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1903_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1903_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1904_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1904_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1904_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1904_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1904_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1905_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1905_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1905_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1905_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1905_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1906_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1906_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1906_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1906_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1906_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1907_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1907_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1907_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1907_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1907_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1908_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1908_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1908_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1908_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1908_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1909_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1909_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1909_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1909_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1909_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1910_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1910_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1910_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1910_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1910_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1911_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1911_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1911_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1911_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1911_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1912_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1912_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1912_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1912_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1912_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1913_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1913_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1913_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1913_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1913_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1914_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1914_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1914_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1914_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1914_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1915_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1915_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1915_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1915_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1915_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1916_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1916_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1916_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1916_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1916_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1917_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1917_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1917_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1917_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1917_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1918_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1918_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1918_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1918_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1918_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1919_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1919_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1919_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1919_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1919_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1920_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1920_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1920_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1920_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1920_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1921_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1921_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1921_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1921_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1921_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1922_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1922_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1922_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1922_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1922_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1923_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1923_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1923_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1923_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1923_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1924_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1924_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1924_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1924_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1924_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1925_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1925_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1925_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1925_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1925_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_50_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_50_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_50_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_50_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1926_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1926_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1926_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1926_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1926_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1927_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1927_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1927_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1927_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1927_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1928_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1928_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1928_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1928_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1928_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1929_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1929_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1929_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1929_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1929_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1930_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1930_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1930_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1930_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1930_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1931_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1931_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1931_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1931_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1931_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1932_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1932_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1932_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1932_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1932_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1933_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1933_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1933_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1933_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1933_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1934_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1934_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1934_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1934_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1934_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1935_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1935_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1935_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1935_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1935_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1936_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1936_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1936_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1936_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1936_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1937_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1937_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1937_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1937_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1937_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1938_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1938_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1938_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1938_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1938_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1939_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1939_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1939_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1939_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1939_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1940_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1940_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1940_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1940_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1940_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1941_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1941_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1941_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1941_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1941_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1942_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1942_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1942_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1942_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1942_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1943_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1943_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1943_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1943_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1943_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1944_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1944_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1944_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1944_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1944_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1945_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1945_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1945_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1945_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1945_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1946_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1946_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1946_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1946_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1946_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1947_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1947_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1947_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1947_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1947_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1948_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1948_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1948_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1948_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1948_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1949_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1949_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1949_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1949_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1949_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1950_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1950_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1950_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1950_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1950_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1951_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1951_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1951_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1951_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1951_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1952_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1952_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1952_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1952_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1952_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1953_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1953_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1953_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1953_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1953_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1954_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1954_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1954_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1954_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1954_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1955_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1955_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1955_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1955_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1955_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1956_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1956_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1956_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1956_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1956_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1957_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1957_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1957_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1957_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1957_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1958_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1958_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1958_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1958_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1958_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1959_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1959_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1959_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1959_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1959_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1960_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1960_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1960_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1960_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1960_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1961_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1961_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1961_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1961_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1961_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1962_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1962_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1962_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1962_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1962_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1963_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1963_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1963_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1963_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1963_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1964_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1964_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1964_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1964_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1964_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1965_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1965_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1965_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1965_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1965_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1966_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1966_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1966_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1966_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1966_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1967_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1967_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1967_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1967_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1967_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1968_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1968_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1968_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1968_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1968_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_51_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_51_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_51_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_51_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_1969_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1969_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1969_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1969_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1969_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1970_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1970_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1970_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1970_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1970_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1971_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1971_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1971_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1971_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1971_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1972_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1972_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1972_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1972_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1972_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1973_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1973_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1973_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1973_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1973_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1974_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1974_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1974_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1974_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1974_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1975_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1975_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1975_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1975_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1975_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1976_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1976_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1976_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1976_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1976_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1977_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1977_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1977_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1977_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1977_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1978_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1978_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1978_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1978_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1978_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1979_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1979_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1979_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1979_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1979_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1980_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1980_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1980_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1980_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1980_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1981_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1981_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1981_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1981_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1981_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1982_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1982_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1982_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1982_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1982_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1983_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1983_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1983_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1983_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1983_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1984_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1984_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1984_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1984_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1984_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1985_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1985_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1985_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1985_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1985_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1986_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1986_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1986_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1986_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1986_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1987_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1987_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1987_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1987_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1987_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1988_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1988_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1988_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1988_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1988_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1989_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1989_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1989_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1989_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1989_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1990_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1990_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1990_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1990_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1990_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1991_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1991_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1991_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1991_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1991_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1992_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1992_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1992_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1992_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1992_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1993_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1993_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1993_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1993_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1993_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1994_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1994_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1994_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1994_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1994_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1995_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1995_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1995_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1995_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1995_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1996_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1996_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1996_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1996_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1996_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1997_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1997_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1997_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1997_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1997_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1998_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1998_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1998_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1998_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1998_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_1999_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_1999_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_1999_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_1999_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_1999_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2000_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2000_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2000_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2000_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2000_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2001_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2001_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2001_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2001_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2001_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2002_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2002_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2002_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2002_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2002_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2003_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2003_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2003_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2003_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2003_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2004_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2004_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2004_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2004_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2004_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2005_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2005_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2005_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2005_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2005_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2006_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2006_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2006_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2006_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2006_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2007_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2007_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2007_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2007_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2007_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2008_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2008_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2008_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2008_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2008_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2009_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2009_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2009_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2009_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2009_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2010_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2010_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2010_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2010_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2010_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2011_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2011_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2011_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2011_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2011_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2012_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2012_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2012_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2012_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2012_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2013_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2013_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2013_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2013_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2013_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2014_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2014_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2014_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2014_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2014_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2015_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2015_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2015_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2015_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2015_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2016_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2016_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2016_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2016_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2016_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_52_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_52_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_52_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_52_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2017_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2017_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2017_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2017_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2017_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2018_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2018_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2018_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2018_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2018_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2019_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2019_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2019_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2019_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2019_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2020_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2020_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2020_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2020_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2020_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2021_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2021_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2021_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2021_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2021_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2022_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2022_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2022_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2022_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2022_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2023_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2023_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2023_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2023_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2023_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2024_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2024_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2024_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2024_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2024_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2025_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2025_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2025_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2025_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2025_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2026_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2026_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2026_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2026_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2026_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2027_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2027_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2027_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2027_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2027_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2028_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2028_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2028_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2028_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2028_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2029_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2029_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2029_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2029_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2029_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2030_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2030_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2030_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2030_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2030_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2031_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2031_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2031_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2031_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2031_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2032_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2032_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2032_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2032_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2032_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2033_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2033_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2033_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2033_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2033_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2034_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2034_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2034_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2034_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2034_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2035_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2035_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2035_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2035_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2035_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2036_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2036_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2036_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2036_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2036_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2037_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2037_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2037_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2037_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2037_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2038_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2038_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2038_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2038_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2038_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2039_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2039_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2039_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2039_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2039_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2040_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2040_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2040_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2040_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2040_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2041_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2041_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2041_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2041_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2041_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2042_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2042_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2042_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2042_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2042_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2043_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2043_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2043_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2043_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2043_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2044_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2044_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2044_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2044_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2044_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2045_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2045_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2045_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2045_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2045_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2046_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2046_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2046_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2046_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2046_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2047_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2047_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2047_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2047_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2047_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2048_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2048_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2048_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2048_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2048_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2049_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2049_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2049_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2049_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2049_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2050_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2050_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2050_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2050_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2050_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2051_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2051_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2051_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2051_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2051_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_53_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_53_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_53_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_53_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2052_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2052_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2052_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2052_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2052_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2053_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2053_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2053_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2053_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2053_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2054_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2054_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2054_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2054_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2054_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2055_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2055_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2055_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2055_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2055_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2056_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2056_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2056_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2056_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2056_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2057_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2057_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2057_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2057_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2057_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2058_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2058_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2058_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2058_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2058_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2059_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2059_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2059_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2059_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2059_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2060_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2060_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2060_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2060_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2060_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2061_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2061_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2061_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2061_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2061_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2062_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2062_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2062_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2062_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2062_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2063_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2063_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2063_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2063_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2063_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2064_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2064_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2064_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2064_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2064_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2065_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2065_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2065_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2065_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2065_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2066_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2066_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2066_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2066_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2066_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2067_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2067_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2067_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2067_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2067_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2068_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2068_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2068_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2068_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2068_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2069_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2069_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2069_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2069_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2069_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2070_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2070_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2070_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2070_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2070_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2071_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2071_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2071_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2071_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2071_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2072_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2072_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2072_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2072_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2072_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2073_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2073_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2073_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2073_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2073_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2074_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2074_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2074_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2074_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2074_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2075_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2075_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2075_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2075_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2075_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2076_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2076_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2076_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2076_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2076_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2077_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2077_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2077_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2077_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2077_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2078_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2078_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2078_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2078_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2078_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2079_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2079_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2079_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2079_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2079_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2080_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2080_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2080_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2080_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2080_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2081_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2081_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2081_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2081_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2081_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2082_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2082_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2082_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2082_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2082_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2083_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2083_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2083_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2083_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2083_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2084_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2084_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2084_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2084_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2084_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2085_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2085_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2085_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2085_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2085_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2086_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2086_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2086_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2086_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2086_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2087_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2087_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2087_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2087_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2087_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2088_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2088_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2088_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2088_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2088_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2089_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2089_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2089_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2089_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2089_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_54_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_54_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_54_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_54_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2090_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2090_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2090_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2090_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2090_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2091_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2091_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2091_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2091_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2091_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2092_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2092_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2092_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2092_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2092_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2093_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2093_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2093_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2093_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2093_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2094_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2094_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2094_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2094_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2094_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2095_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2095_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2095_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2095_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2095_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2096_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2096_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2096_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2096_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2096_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2097_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2097_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2097_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2097_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2097_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2098_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2098_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2098_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2098_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2098_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2099_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2099_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2099_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2099_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2099_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2100_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2100_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2100_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2100_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2100_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2101_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2101_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2101_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2101_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2101_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2102_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2102_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2102_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2102_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2102_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2103_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2103_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2103_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2103_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2103_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2104_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2104_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2104_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2104_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2104_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2105_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2105_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2105_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2105_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2105_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2106_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2106_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2106_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2106_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2106_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2107_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2107_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2107_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2107_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2107_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2108_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2108_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2108_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2108_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2108_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2109_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2109_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2109_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2109_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2109_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2110_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2110_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2110_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2110_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2110_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2111_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2111_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2111_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2111_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2111_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2112_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2112_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2112_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2112_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2112_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2113_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2113_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2113_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2113_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2113_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2114_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2114_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2114_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2114_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2114_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2115_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2115_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2115_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2115_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2115_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2116_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2116_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2116_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2116_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2116_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_55_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_55_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_55_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_55_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2117_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2117_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2117_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2117_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2117_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2118_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2118_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2118_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2118_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2118_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2119_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2119_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2119_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2119_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2119_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2120_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2120_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2120_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2120_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2120_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2121_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2121_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2121_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2121_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2121_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2122_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2122_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2122_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2122_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2122_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2123_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2123_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2123_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2123_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2123_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2124_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2124_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2124_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2124_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2124_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2125_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2125_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2125_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2125_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2125_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2126_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2126_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2126_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2126_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2126_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2127_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2127_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2127_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2127_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2127_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2128_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2128_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2128_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2128_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2128_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2129_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2129_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2129_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2129_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2129_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2130_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2130_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2130_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2130_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2130_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2131_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2131_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2131_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2131_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2131_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2132_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2132_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2132_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2132_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2132_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2133_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2133_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2133_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2133_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2133_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_56_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_56_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_56_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_56_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2134_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2134_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2134_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2134_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2134_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2135_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2135_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2135_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2135_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2135_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2136_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2136_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2136_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2136_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2136_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2137_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2137_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2137_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2137_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2137_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2138_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2138_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2138_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2138_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2138_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2139_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2139_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2139_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2139_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2139_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2140_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2140_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2140_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2140_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2140_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2141_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2141_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2141_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2141_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2141_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2142_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2142_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2142_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2142_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2142_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2143_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2143_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2143_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2143_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2143_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2144_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2144_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2144_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2144_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2144_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2145_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2145_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2145_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2145_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2145_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2146_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2146_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2146_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2146_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2146_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2147_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2147_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2147_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2147_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2147_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2148_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2148_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2148_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2148_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2148_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2149_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2149_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2149_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2149_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2149_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2150_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2150_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2150_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2150_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2150_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2151_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2151_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2151_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2151_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2151_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2152_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2152_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2152_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2152_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2152_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2153_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2153_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2153_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2153_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2153_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2154_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2154_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2154_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2154_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2154_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2155_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2155_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2155_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2155_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2155_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2156_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2156_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2156_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2156_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2156_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2157_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2157_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2157_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2157_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2157_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2158_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2158_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2158_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2158_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2158_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2159_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2159_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2159_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2159_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2159_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2160_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2160_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2160_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2160_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2160_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2161_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2161_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2161_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2161_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2161_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2162_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2162_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2162_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2162_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2162_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2163_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2163_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2163_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2163_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2163_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_57_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_57_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_57_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_57_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2164_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2164_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2164_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2164_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2164_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2165_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2165_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2165_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2165_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2165_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2166_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2166_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2166_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2166_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2166_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2167_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2167_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2167_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2167_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2167_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2168_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2168_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2168_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2168_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2168_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2169_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2169_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2169_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2169_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2169_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2170_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2170_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2170_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2170_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2170_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2171_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2171_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2171_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2171_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2171_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2172_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2172_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2172_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2172_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2172_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2173_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2173_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2173_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2173_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2173_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2174_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2174_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2174_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2174_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2174_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2175_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2175_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2175_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2175_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2175_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2176_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2176_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2176_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2176_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2176_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2177_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2177_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2177_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2177_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2177_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2178_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2178_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2178_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2178_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2178_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_58_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_58_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_58_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_58_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2179_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2179_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2179_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2179_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2179_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2180_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2180_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2180_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2180_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2180_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2181_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2181_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2181_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2181_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2181_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_59_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_59_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_59_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_59_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2182_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2182_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2182_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2182_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2182_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2183_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2183_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2183_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2183_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2183_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2184_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2184_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2184_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2184_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2184_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2185_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2185_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2185_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2185_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2185_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2186_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2186_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2186_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2186_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2186_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2187_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2187_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2187_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2187_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2187_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2188_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2188_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2188_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2188_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2188_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2189_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2189_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2189_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2189_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2189_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2190_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2190_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2190_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2190_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2190_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2191_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2191_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2191_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2191_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2191_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2192_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2192_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2192_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2192_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2192_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2193_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2193_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2193_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2193_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2193_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_60_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_60_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_60_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_60_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_61_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_61_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_61_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_61_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2194_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2194_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2194_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2194_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2194_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2195_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2195_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2195_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2195_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2195_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2196_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2196_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2196_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2196_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2196_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2197_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2197_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2197_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2197_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2197_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2198_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2198_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2198_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2198_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2198_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_62_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_62_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_62_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_62_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2199_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2199_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2199_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2199_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2199_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_63_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_63_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_63_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_63_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2200_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2200_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2200_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2200_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2200_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_64_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_64_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_64_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_64_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2201_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2201_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2201_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2201_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2201_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_65_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_65_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_65_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_65_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_66_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_66_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_66_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_66_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_67_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_67_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_67_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_67_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_68_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_68_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_68_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_68_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_69_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_69_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_69_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_69_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2202_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2202_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2202_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2202_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2202_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2203_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2203_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2203_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2203_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2203_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_70_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_70_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_70_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_70_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_71_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_71_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_71_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_71_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2204_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2204_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2204_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2204_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2204_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2205_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2205_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2205_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2205_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2205_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2206_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2206_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2206_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2206_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2206_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2207_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2207_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2207_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2207_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2207_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2208_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2208_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2208_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2208_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2208_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2209_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2209_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2209_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2209_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2209_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2210_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2210_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2210_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2210_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2210_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2211_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2211_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2211_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2211_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2211_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2212_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2212_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2212_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2212_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2212_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2213_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2213_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2213_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2213_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2213_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2214_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2214_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2214_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2214_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2214_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2215_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2215_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2215_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2215_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2215_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2216_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2216_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2216_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2216_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2216_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2217_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2217_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2217_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2217_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2217_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_72_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_72_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_72_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_72_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2218_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2218_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2218_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2218_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2218_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2219_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2219_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2219_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2219_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2219_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2220_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2220_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2220_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2220_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2220_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2221_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2221_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2221_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2221_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2221_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_73_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_73_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_73_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_73_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2222_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2222_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2222_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2222_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2222_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2223_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2223_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2223_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2223_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2223_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2224_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2224_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2224_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2224_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2224_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2225_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2225_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2225_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2225_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2225_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2226_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2226_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2226_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2226_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2226_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2227_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2227_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2227_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2227_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2227_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2228_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2228_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2228_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2228_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2228_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2229_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2229_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2229_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2229_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2229_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2230_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2230_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2230_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2230_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2230_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2231_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2231_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2231_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2231_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2231_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2232_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2232_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2232_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2232_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2232_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2233_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2233_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2233_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2233_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2233_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2234_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2234_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2234_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2234_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2234_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2235_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2235_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2235_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2235_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2235_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2236_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2236_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2236_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2236_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2236_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2237_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2237_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2237_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2237_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2237_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2238_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2238_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2238_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2238_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2238_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2239_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2239_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2239_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2239_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2239_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_74_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_74_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_74_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_74_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2240_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2240_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2240_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2240_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2240_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2241_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2241_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2241_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2241_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2241_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2242_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2242_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2242_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2242_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2242_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2243_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2243_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2243_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2243_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2243_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2244_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2244_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2244_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2244_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2244_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2245_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2245_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2245_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2245_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2245_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2246_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2246_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2246_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2246_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2246_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2247_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2247_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2247_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2247_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2247_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2248_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2248_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2248_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2248_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2248_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2249_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2249_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2249_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2249_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2249_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2250_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2250_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2250_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2250_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2250_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2251_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2251_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2251_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2251_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2251_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2252_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2252_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2252_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2252_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2252_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2253_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2253_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2253_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2253_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2253_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2254_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2254_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2254_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2254_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2254_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2255_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2255_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2255_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2255_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2255_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2256_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2256_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2256_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2256_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2256_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2257_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2257_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2257_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2257_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2257_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2258_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2258_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2258_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2258_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2258_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2259_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2259_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2259_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2259_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2259_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2260_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2260_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2260_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2260_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2260_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2261_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2261_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2261_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2261_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2261_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2262_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2262_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2262_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2262_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2262_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2263_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2263_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2263_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2263_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2263_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2264_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2264_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2264_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2264_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2264_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2265_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2265_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2265_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2265_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2265_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2266_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2266_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2266_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2266_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2266_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2267_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2267_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2267_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2267_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2267_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2268_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2268_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2268_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2268_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2268_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2269_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2269_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2269_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2269_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2269_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2270_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2270_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2270_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2270_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2270_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2271_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2271_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2271_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2271_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2271_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2272_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2272_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2272_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2272_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2272_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2273_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2273_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2273_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2273_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2273_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2274_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2274_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2274_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2274_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2274_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2275_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2275_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2275_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2275_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2275_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2276_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2276_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2276_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2276_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2276_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2277_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2277_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2277_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2277_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2277_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2278_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2278_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2278_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2278_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2278_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2279_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2279_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2279_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2279_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2279_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2280_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2280_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2280_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2280_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2280_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2281_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2281_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2281_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2281_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2281_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2282_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2282_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2282_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2282_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2282_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2283_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2283_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2283_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2283_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2283_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2284_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2284_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2284_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2284_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2284_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2285_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2285_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2285_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2285_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2285_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2286_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2286_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2286_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2286_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2286_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2287_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2287_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2287_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2287_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2287_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2288_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2288_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2288_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2288_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2288_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2289_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2289_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2289_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2289_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2289_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2290_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2290_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2290_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2290_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2290_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2291_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2291_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2291_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2291_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2291_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2292_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2292_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2292_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2292_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2292_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2293_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2293_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2293_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2293_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2293_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2294_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2294_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2294_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2294_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2294_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2295_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2295_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2295_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2295_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2295_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2296_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2296_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2296_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2296_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2296_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2297_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2297_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2297_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2297_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2297_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2298_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2298_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2298_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2298_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2298_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2299_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2299_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2299_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2299_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2299_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2300_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2300_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2300_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2300_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2300_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2301_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2301_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2301_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2301_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2301_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2302_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2302_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2302_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2302_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2302_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2303_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2303_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2303_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2303_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2303_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2304_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2304_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2304_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2304_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2304_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2305_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2305_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2305_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2305_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2305_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2306_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2306_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2306_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2306_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2306_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2307_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2307_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2307_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2307_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2307_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2308_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2308_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2308_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2308_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2308_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2309_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2309_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2309_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2309_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2309_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2310_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2310_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2310_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2310_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2310_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2311_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2311_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2311_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2311_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2311_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2312_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2312_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2312_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2312_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2312_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2313_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2313_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2313_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2313_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2313_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2314_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2314_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2314_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2314_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2314_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2315_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2315_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2315_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2315_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2315_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2316_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2316_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2316_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2316_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2316_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2317_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2317_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2317_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2317_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2317_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2318_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2318_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2318_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2318_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2318_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2319_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2319_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2319_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2319_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2319_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2320_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2320_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2320_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2320_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2320_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2321_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2321_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2321_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2321_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2321_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2322_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2322_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2322_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2322_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2322_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2323_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2323_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2323_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2323_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2323_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2324_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2324_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2324_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2324_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2324_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2325_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2325_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2325_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2325_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2325_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2326_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2326_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2326_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2326_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2326_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2327_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2327_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2327_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2327_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2327_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2328_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2328_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2328_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2328_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2328_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2329_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2329_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2329_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2329_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2329_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2330_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2330_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2330_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2330_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2330_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2331_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2331_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2331_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2331_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2331_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2332_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2332_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2332_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2332_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2332_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2333_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2333_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2333_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2333_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2333_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2334_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2334_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2334_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2334_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2334_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2335_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2335_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2335_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2335_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2335_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2336_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2336_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2336_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2336_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2336_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2337_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2337_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2337_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2337_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2337_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2338_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2338_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2338_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2338_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2338_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_75_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_75_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_75_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_75_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2339_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2339_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2339_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2339_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2339_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2340_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2340_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2340_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2340_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2340_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2341_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2341_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2341_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2341_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2341_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2342_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2342_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2342_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2342_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2342_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2343_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2343_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2343_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2343_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2343_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2344_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2344_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2344_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2344_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2344_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_76_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_76_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_76_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_76_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2345_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2345_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2345_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2345_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2345_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2346_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2346_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2346_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2346_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2346_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2347_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2347_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2347_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2347_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2347_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2348_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2348_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2348_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2348_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2348_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2349_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2349_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2349_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2349_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2349_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2350_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2350_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2350_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2350_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2350_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2351_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2351_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2351_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2351_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2351_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2352_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2352_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2352_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2352_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2352_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2353_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2353_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2353_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2353_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2353_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2354_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2354_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2354_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2354_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2354_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2355_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2355_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2355_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2355_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2355_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2356_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2356_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2356_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2356_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2356_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2357_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2357_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2357_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2357_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2357_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2358_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2358_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2358_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2358_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2358_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2359_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2359_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2359_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2359_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2359_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2360_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2360_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2360_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2360_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2360_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2361_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2361_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2361_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2361_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2361_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2362_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2362_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2362_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2362_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2362_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2363_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2363_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2363_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2363_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2363_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2364_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2364_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2364_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2364_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2364_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2365_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2365_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2365_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2365_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2365_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2366_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2366_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2366_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2366_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2366_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2367_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2367_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2367_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2367_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2367_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2368_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2368_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2368_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2368_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2368_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2369_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2369_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2369_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2369_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2369_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2370_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2370_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2370_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2370_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2370_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2371_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2371_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2371_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2371_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2371_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2372_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2372_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2372_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2372_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2372_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2373_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2373_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2373_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2373_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2373_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2374_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2374_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2374_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2374_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2374_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2375_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2375_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2375_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2375_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2375_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2376_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2376_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2376_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2376_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2376_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2377_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2377_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2377_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2377_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2377_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2378_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2378_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2378_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2378_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2378_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2379_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2379_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2379_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2379_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2379_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2380_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2380_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2380_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2380_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2380_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2381_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2381_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2381_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2381_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2381_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2382_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2382_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2382_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2382_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2382_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2383_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2383_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2383_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2383_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2383_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2384_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2384_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2384_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2384_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2384_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2385_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2385_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2385_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2385_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2385_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_77_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_77_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_77_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_77_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2386_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2386_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2386_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2386_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2386_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2387_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2387_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2387_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2387_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2387_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2388_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2388_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2388_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2388_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2388_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2389_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2389_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2389_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2389_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2389_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2390_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2390_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2390_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2390_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2390_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2391_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2391_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2391_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2391_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2391_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2392_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2392_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2392_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2392_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2392_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2393_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2393_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2393_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2393_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2393_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2394_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2394_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2394_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2394_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2394_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2395_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2395_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2395_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2395_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2395_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2396_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2396_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2396_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2396_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2396_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2397_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2397_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2397_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2397_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2397_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2398_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2398_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2398_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2398_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2398_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2399_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2399_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2399_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2399_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2399_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2400_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2400_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2400_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2400_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2400_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2401_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2401_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2401_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2401_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2401_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2402_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2402_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2402_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2402_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2402_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2403_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2403_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2403_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2403_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2403_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2404_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2404_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2404_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2404_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2404_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2405_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2405_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2405_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2405_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2405_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2406_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2406_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2406_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2406_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2406_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2407_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2407_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2407_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2407_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2407_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2408_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2408_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2408_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2408_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2408_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2409_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2409_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2409_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2409_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2409_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2410_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2410_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2410_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2410_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2410_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2411_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2411_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2411_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2411_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2411_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2412_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2412_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2412_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2412_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2412_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2413_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2413_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2413_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2413_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2413_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2414_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2414_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2414_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2414_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2414_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2415_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2415_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2415_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2415_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2415_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2416_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2416_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2416_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2416_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2416_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2417_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2417_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2417_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2417_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2417_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2418_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2418_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2418_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2418_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2418_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2419_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2419_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2419_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2419_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2419_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2420_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2420_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2420_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2420_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2420_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2421_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2421_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2421_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2421_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2421_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2422_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2422_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2422_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2422_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2422_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2423_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2423_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2423_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2423_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2423_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2424_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2424_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2424_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2424_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2424_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2425_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2425_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2425_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2425_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2425_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2426_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2426_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2426_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2426_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2426_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2427_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2427_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2427_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2427_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2427_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2428_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2428_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2428_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2428_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2428_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2429_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2429_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2429_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2429_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2429_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2430_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2430_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2430_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2430_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2430_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2431_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2431_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2431_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2431_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2431_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2432_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2432_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2432_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2432_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2432_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2433_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2433_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2433_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2433_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2433_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2434_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2434_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2434_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2434_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2434_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2435_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2435_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2435_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2435_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2435_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2436_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2436_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2436_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2436_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2436_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2437_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2437_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2437_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2437_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2437_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2438_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2438_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2438_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2438_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2438_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2439_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2439_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2439_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2439_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2439_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2440_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2440_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2440_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2440_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2440_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2441_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2441_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2441_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2441_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2441_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2442_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2442_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2442_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2442_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2442_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2443_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2443_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2443_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2443_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2443_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2444_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2444_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2444_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2444_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2444_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2445_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2445_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2445_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2445_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2445_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2446_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2446_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2446_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2446_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2446_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2447_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2447_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2447_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2447_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2447_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2448_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2448_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2448_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2448_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2448_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2449_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2449_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2449_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2449_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2449_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2450_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2450_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2450_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2450_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2450_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2451_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2451_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2451_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2451_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2451_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2452_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2452_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2452_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2452_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2452_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2453_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2453_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2453_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2453_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2453_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2454_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2454_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2454_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2454_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2454_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2455_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2455_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2455_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2455_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2455_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2456_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2456_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2456_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2456_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2456_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2457_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2457_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2457_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2457_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2457_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2458_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2458_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2458_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2458_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2458_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2459_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2459_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2459_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2459_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2459_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2460_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2460_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2460_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2460_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2460_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2461_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2461_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2461_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2461_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2461_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2462_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2462_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2462_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2462_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2462_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2463_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2463_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2463_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2463_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2463_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2464_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2464_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2464_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2464_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2464_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2465_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2465_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2465_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2465_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2465_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2466_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2466_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2466_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2466_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2466_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2467_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2467_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2467_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2467_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2467_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2468_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2468_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2468_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2468_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2468_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2469_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2469_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2469_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2469_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2469_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2470_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2470_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2470_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2470_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2470_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2471_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2471_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2471_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2471_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2471_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2472_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2472_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2472_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2472_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2472_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2473_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2473_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2473_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2473_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2473_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2474_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2474_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2474_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2474_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2474_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2475_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2475_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2475_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2475_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2475_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2476_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2476_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2476_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2476_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2476_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2477_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2477_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2477_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2477_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2477_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2478_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2478_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2478_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2478_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2478_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2479_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2479_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2479_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2479_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2479_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2480_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2480_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2480_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2480_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2480_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2481_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2481_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2481_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2481_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2481_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2482_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2482_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2482_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2482_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2482_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2483_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2483_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2483_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2483_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2483_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2484_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2484_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2484_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2484_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2484_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2485_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2485_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2485_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2485_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2485_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2486_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2486_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2486_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2486_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2486_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2487_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2487_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2487_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2487_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2487_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2488_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2488_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2488_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2488_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2488_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2489_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2489_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2489_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2489_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2489_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2490_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2490_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2490_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2490_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2490_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2491_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2491_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2491_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2491_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2491_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2492_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2492_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2492_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2492_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2492_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2493_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2493_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2493_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2493_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2493_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2494_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2494_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2494_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2494_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2494_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2495_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2495_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2495_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2495_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2495_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2496_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2496_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2496_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2496_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2496_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2497_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2497_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2497_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2497_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2497_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2498_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2498_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2498_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2498_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2498_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2499_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2499_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2499_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2499_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2499_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2500_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2500_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2500_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2500_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2500_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2501_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2501_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2501_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2501_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2501_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2502_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2502_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2502_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2502_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2502_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2503_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2503_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2503_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2503_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2503_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2504_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2504_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2504_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2504_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2504_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2505_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2505_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2505_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2505_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2505_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_78_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_78_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_78_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_78_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2506_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2506_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2506_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2506_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2506_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2507_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2507_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2507_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2507_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2507_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2508_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2508_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2508_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2508_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2508_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2509_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2509_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2509_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2509_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2509_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2510_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2510_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2510_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2510_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2510_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2511_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2511_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2511_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2511_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2511_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2512_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2512_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2512_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2512_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2512_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2513_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2513_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2513_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2513_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2513_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2514_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2514_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2514_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2514_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2514_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2515_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2515_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2515_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2515_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2515_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2516_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2516_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2516_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2516_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2516_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2517_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2517_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2517_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2517_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2517_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2518_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2518_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2518_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2518_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2518_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2519_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2519_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2519_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2519_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2519_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2520_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2520_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2520_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2520_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2520_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2521_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2521_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2521_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2521_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2521_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2522_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2522_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2522_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2522_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2522_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2523_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2523_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2523_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2523_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2523_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2524_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2524_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2524_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2524_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2524_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2525_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2525_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2525_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2525_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2525_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2526_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2526_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2526_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2526_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2526_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2527_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2527_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2527_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2527_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2527_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2528_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2528_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2528_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2528_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2528_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2529_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2529_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2529_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2529_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2529_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2530_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2530_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2530_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2530_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2530_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2531_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2531_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2531_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2531_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2531_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2532_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2532_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2532_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2532_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2532_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2533_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2533_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2533_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2533_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2533_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2534_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2534_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2534_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2534_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2534_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2535_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2535_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2535_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2535_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2535_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2536_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2536_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2536_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2536_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2536_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2537_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2537_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2537_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2537_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2537_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2538_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2538_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2538_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2538_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2538_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2539_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2539_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2539_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2539_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2539_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2540_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2540_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2540_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2540_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2540_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2541_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2541_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2541_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2541_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2541_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2542_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2542_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2542_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2542_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2542_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2543_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2543_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2543_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2543_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2543_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2544_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2544_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2544_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2544_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2544_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2545_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2545_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2545_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2545_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2545_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2546_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2546_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2546_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2546_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2546_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2547_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2547_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2547_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2547_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2547_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2548_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2548_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2548_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2548_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2548_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2549_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2549_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2549_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2549_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2549_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_79_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_79_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_79_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_79_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2550_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2550_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2550_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2550_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2550_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2551_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2551_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2551_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2551_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2551_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2552_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2552_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2552_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2552_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2552_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2553_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2553_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2553_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2553_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2553_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2554_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2554_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2554_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2554_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2554_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2555_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2555_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2555_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2555_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2555_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2556_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2556_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2556_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2556_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2556_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2557_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2557_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2557_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2557_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2557_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2558_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2558_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2558_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2558_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2558_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2559_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2559_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2559_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2559_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2559_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2560_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2560_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2560_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2560_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2560_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2561_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2561_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2561_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2561_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2561_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2562_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2562_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2562_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2562_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2562_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2563_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2563_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2563_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2563_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2563_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2564_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2564_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2564_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2564_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2564_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2565_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2565_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2565_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2565_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2565_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2566_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2566_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2566_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2566_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2566_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2567_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2567_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2567_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2567_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2567_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2568_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2568_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2568_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2568_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2568_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2569_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2569_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2569_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2569_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2569_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2570_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2570_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2570_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2570_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2570_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2571_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2571_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2571_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2571_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2571_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2572_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2572_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2572_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2572_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2572_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2573_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2573_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2573_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2573_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2573_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2574_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2574_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2574_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2574_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2574_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2575_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2575_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2575_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2575_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2575_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2576_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2576_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2576_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2576_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2576_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2577_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2577_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2577_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2577_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2577_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2578_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2578_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2578_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2578_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2578_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2579_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2579_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2579_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2579_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2579_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2580_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2580_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2580_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2580_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2580_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2581_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2581_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2581_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2581_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2581_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2582_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2582_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2582_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2582_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2582_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2583_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2583_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2583_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2583_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2583_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2584_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2584_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2584_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2584_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2584_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2585_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2585_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2585_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2585_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2585_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2586_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2586_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2586_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2586_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2586_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2587_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2587_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2587_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2587_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2587_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2588_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2588_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2588_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2588_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2588_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2589_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2589_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2589_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2589_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2589_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2590_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2590_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2590_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2590_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2590_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2591_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2591_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2591_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2591_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2591_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2592_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2592_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2592_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2592_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2592_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2593_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2593_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2593_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2593_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2593_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2594_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2594_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2594_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2594_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2594_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2595_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2595_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2595_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2595_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2595_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2596_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2596_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2596_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2596_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2596_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2597_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2597_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2597_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2597_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2597_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2598_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2598_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2598_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2598_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2598_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2599_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2599_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2599_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2599_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2599_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2600_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2600_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2600_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2600_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2600_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2601_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2601_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2601_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2601_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2601_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2602_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2602_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2602_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2602_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2602_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2603_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2603_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2603_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2603_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2603_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_80_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_80_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_80_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_80_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2604_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2604_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2604_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2604_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2604_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2605_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2605_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2605_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2605_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2605_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2606_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2606_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2606_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2606_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2606_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2607_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2607_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2607_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2607_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2607_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2608_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2608_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2608_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2608_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2608_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2609_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2609_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2609_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2609_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2609_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2610_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2610_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2610_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2610_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2610_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2611_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2611_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2611_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2611_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2611_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2612_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2612_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2612_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2612_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2612_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2613_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2613_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2613_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2613_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2613_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2614_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2614_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2614_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2614_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2614_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2615_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2615_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2615_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2615_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2615_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2616_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2616_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2616_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2616_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2616_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2617_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2617_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2617_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2617_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2617_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2618_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2618_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2618_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2618_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2618_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2619_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2619_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2619_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2619_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2619_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2620_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2620_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2620_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2620_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2620_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2621_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2621_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2621_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2621_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2621_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2622_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2622_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2622_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2622_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2622_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2623_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2623_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2623_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2623_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2623_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2624_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2624_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2624_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2624_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2624_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2625_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2625_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2625_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2625_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2625_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2626_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2626_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2626_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2626_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2626_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2627_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2627_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2627_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2627_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2627_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2628_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2628_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2628_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2628_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2628_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2629_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2629_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2629_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2629_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2629_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2630_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2630_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2630_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2630_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2630_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2631_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2631_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2631_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2631_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2631_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2632_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2632_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2632_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2632_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2632_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2633_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2633_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2633_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2633_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2633_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2634_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2634_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2634_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2634_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2634_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2635_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2635_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2635_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2635_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2635_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2636_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2636_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2636_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2636_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2636_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2637_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2637_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2637_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2637_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2637_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2638_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2638_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2638_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2638_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2638_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2639_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2639_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2639_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2639_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2639_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2640_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2640_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2640_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2640_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2640_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2641_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2641_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2641_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2641_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2641_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2642_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2642_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2642_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2642_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2642_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2643_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2643_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2643_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2643_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2643_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2644_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2644_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2644_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2644_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2644_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_81_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_81_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_81_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_81_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2645_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2645_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2645_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2645_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2645_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2646_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2646_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2646_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2646_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2646_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2647_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2647_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2647_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2647_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2647_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2648_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2648_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2648_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2648_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2648_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2649_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2649_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2649_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2649_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2649_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2650_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2650_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2650_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2650_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2650_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2651_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2651_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2651_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2651_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2651_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2652_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2652_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2652_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2652_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2652_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2653_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2653_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2653_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2653_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2653_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2654_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2654_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2654_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2654_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2654_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2655_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2655_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2655_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2655_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2655_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2656_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2656_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2656_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2656_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2656_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2657_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2657_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2657_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2657_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2657_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2658_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2658_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2658_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2658_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2658_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2659_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2659_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2659_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2659_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2659_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2660_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2660_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2660_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2660_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2660_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2661_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2661_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2661_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2661_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2661_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2662_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2662_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2662_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2662_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2662_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2663_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2663_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2663_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2663_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2663_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2664_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2664_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2664_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2664_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2664_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2665_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2665_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2665_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2665_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2665_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2666_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2666_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2666_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2666_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2666_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2667_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2667_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2667_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2667_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2667_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2668_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2668_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2668_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2668_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2668_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2669_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2669_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2669_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2669_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2669_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2670_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2670_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2670_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2670_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2670_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2671_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2671_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2671_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2671_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2671_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2672_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2672_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2672_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2672_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2672_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2673_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2673_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2673_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2673_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2673_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2674_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2674_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2674_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2674_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2674_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2675_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2675_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2675_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2675_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2675_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2676_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2676_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2676_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2676_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2676_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2677_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2677_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2677_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2677_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2677_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2678_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2678_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2678_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2678_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2678_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2679_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2679_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2679_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2679_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2679_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2680_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2680_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2680_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2680_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2680_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2681_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2681_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2681_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2681_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2681_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2682_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2682_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2682_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2682_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2682_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2683_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2683_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2683_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2683_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2683_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2684_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2684_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2684_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2684_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2684_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2685_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2685_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2685_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2685_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2685_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2686_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2686_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2686_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2686_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2686_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2687_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2687_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2687_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2687_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2687_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2688_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2688_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2688_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2688_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2688_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2689_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2689_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2689_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2689_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2689_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2690_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2690_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2690_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2690_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2690_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2691_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2691_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2691_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2691_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2691_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_82_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_82_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_82_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_82_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2692_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2692_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2692_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2692_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2692_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2693_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2693_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2693_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2693_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2693_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2694_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2694_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2694_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2694_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2694_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2695_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2695_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2695_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2695_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2695_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2696_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2696_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2696_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2696_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2696_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_83_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_83_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_83_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_83_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2697_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2697_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2697_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2697_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2697_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2698_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2698_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2698_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2698_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2698_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2699_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2699_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2699_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2699_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2699_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2700_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2700_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2700_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2700_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2700_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2701_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2701_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2701_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2701_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2701_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2702_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2702_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2702_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2702_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2702_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2703_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2703_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2703_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2703_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2703_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2704_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2704_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2704_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2704_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2704_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2705_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2705_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2705_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2705_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2705_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2706_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2706_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2706_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2706_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2706_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2707_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2707_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2707_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2707_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2707_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2708_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2708_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2708_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2708_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2708_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2709_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2709_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2709_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2709_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2709_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2710_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2710_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2710_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2710_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2710_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2711_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2711_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2711_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2711_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2711_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2712_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2712_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2712_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2712_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2712_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2713_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2713_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2713_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2713_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2713_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2714_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2714_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2714_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2714_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2714_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2715_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2715_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2715_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2715_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2715_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2716_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2716_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2716_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2716_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2716_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2717_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2717_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2717_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2717_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2717_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2718_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2718_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2718_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2718_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2718_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2719_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2719_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2719_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2719_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2719_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2720_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2720_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2720_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2720_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2720_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2721_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2721_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2721_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2721_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2721_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2722_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2722_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2722_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2722_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2722_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2723_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2723_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2723_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2723_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2723_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2724_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2724_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2724_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2724_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2724_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_84_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_84_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_84_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_84_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2725_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2725_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2725_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2725_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2725_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2726_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2726_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2726_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2726_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2726_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2727_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2727_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2727_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2727_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2727_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2728_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2728_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2728_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2728_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2728_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2729_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2729_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2729_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2729_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2729_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2730_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2730_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2730_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2730_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2730_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2731_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2731_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2731_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2731_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2731_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2732_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2732_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2732_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2732_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2732_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2733_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2733_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2733_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2733_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2733_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2734_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2734_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2734_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2734_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2734_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2735_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2735_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2735_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2735_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2735_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2736_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2736_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2736_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2736_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2736_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2737_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2737_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2737_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2737_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2737_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2738_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2738_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2738_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2738_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2738_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2739_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2739_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2739_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2739_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2739_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2740_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2740_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2740_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2740_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2740_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2741_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2741_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2741_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2741_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2741_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2742_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2742_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2742_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2742_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2742_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2743_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2743_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2743_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2743_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2743_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2744_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2744_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2744_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2744_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2744_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2745_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2745_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2745_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2745_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2745_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2746_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2746_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2746_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2746_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2746_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2747_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2747_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2747_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2747_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2747_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2748_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2748_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2748_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2748_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2748_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2749_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2749_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2749_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2749_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2749_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2750_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2750_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2750_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2750_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2750_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_85_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_85_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_85_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_85_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2751_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2751_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2751_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2751_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2751_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2752_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2752_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2752_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2752_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2752_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2753_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2753_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2753_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2753_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2753_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2754_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2754_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2754_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2754_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2754_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2755_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2755_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2755_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2755_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2755_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2756_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2756_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2756_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2756_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2756_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2757_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2757_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2757_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2757_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2757_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2758_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2758_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2758_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2758_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2758_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2759_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2759_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2759_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2759_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2759_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2760_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2760_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2760_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2760_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2760_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2761_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2761_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2761_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2761_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2761_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2762_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2762_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2762_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2762_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2762_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2763_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2763_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2763_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2763_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2763_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2764_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2764_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2764_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2764_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2764_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2765_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2765_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2765_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2765_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2765_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2766_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2766_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2766_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2766_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2766_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2767_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2767_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2767_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2767_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2767_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2768_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2768_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2768_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2768_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2768_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2769_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2769_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2769_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2769_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2769_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_86_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_86_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_86_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_86_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2770_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2770_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2770_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2770_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2770_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2771_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2771_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2771_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2771_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2771_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2772_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2772_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2772_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2772_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2772_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2773_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2773_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2773_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2773_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2773_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2774_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2774_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2774_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2774_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2774_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2775_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2775_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2775_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2775_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2775_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2776_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2776_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2776_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2776_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2776_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2777_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2777_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2777_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2777_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2777_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2778_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2778_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2778_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2778_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2778_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_87_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_87_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_87_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_87_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_88_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_88_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_88_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_88_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2779_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2779_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2779_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2779_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2779_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_89_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_89_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_89_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_89_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2780_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2780_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2780_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2780_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2780_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2781_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2781_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2781_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2781_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2781_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2782_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2782_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2782_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2782_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2782_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2783_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2783_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2783_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2783_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2783_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_90_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_90_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_90_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_90_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_91_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_91_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_91_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_91_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_92_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_92_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_92_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_92_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_93_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_93_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_93_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_93_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_94_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_94_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_94_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_94_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_95_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_95_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_95_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_95_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2784_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2784_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2784_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2784_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2784_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_96_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_96_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_96_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_96_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2785_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2785_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2785_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2785_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2785_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2786_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2786_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2786_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2786_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2786_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2787_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2787_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2787_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2787_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2787_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2788_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2788_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2788_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2788_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2788_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2789_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2789_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2789_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2789_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2789_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2790_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2790_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2790_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2790_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2790_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2791_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2791_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2791_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2791_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2791_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2792_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2792_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2792_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2792_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2792_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2793_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2793_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2793_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2793_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2793_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2794_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2794_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2794_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2794_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2794_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2795_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2795_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2795_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2795_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2795_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2796_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2796_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2796_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2796_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2796_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2797_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2797_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2797_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2797_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2797_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2798_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2798_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2798_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2798_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2798_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2799_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2799_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2799_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2799_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2799_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2800_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2800_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2800_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2800_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2800_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2801_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2801_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2801_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2801_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2801_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2802_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2802_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2802_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2802_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2802_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2803_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2803_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2803_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2803_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2803_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2804_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2804_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2804_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2804_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2804_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2805_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2805_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2805_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2805_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2805_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2806_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2806_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2806_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2806_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2806_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2807_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2807_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2807_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2807_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2807_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2808_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2808_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2808_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2808_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2808_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2809_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2809_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2809_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2809_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2809_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2810_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2810_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2810_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2810_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2810_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2811_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2811_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2811_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2811_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2811_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2812_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2812_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2812_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2812_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2812_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2813_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2813_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2813_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2813_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2813_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2814_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2814_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2814_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2814_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2814_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2815_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2815_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2815_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2815_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2815_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2816_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2816_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2816_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2816_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2816_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2817_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2817_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2817_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2817_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2817_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2818_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2818_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2818_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2818_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2818_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2819_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2819_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2819_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2819_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2819_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2820_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2820_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2820_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2820_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2820_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2821_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2821_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2821_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2821_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2821_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_97_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_97_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_97_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_97_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2822_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2822_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2822_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2822_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2822_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2823_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2823_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2823_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2823_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2823_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2824_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2824_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2824_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2824_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2824_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2825_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2825_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2825_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2825_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2825_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2826_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2826_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2826_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2826_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2826_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2827_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2827_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2827_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2827_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2827_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2828_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2828_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2828_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2828_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2828_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2829_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2829_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2829_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2829_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2829_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2830_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2830_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2830_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2830_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2830_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2831_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2831_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2831_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2831_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2831_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2832_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2832_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2832_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2832_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2832_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2833_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2833_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2833_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2833_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2833_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2834_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2834_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2834_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2834_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2834_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2835_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2835_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2835_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2835_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2835_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2836_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2836_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2836_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2836_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2836_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2837_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2837_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2837_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2837_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2837_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2838_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2838_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2838_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2838_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2838_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2839_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2839_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2839_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2839_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2839_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_98_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_98_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_98_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_98_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2840_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2840_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2840_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2840_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2840_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2841_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2841_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2841_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2841_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2841_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2842_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2842_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2842_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2842_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2842_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_99_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_99_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_99_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_99_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2843_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2843_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2843_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2843_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2843_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2844_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2844_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2844_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2844_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2844_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2845_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2845_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2845_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2845_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2845_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_100_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_100_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_100_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_100_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2846_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2846_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2846_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2846_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2846_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2847_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2847_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2847_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2847_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2847_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2848_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2848_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2848_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2848_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2848_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2849_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2849_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2849_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2849_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2849_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2850_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2850_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2850_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2850_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2850_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2851_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2851_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2851_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2851_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2851_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2852_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2852_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2852_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2852_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2852_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2853_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2853_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2853_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2853_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2853_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2854_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2854_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2854_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2854_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2854_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2855_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2855_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2855_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2855_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2855_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2856_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2856_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2856_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2856_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2856_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2857_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2857_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2857_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2857_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2857_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2858_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2858_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2858_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2858_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2858_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2859_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2859_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2859_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2859_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2859_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2860_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2860_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2860_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2860_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2860_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2861_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2861_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2861_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2861_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2861_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2862_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2862_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2862_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2862_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2862_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2863_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2863_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2863_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2863_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2863_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2864_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2864_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2864_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2864_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2864_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2865_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2865_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2865_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2865_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2865_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2866_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2866_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2866_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2866_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2866_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2867_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2867_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2867_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2867_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2867_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2868_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2868_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2868_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2868_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2868_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2869_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2869_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2869_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2869_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2869_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2870_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2870_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2870_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2870_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2870_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2871_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2871_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2871_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2871_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2871_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2872_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2872_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2872_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2872_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2872_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2873_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2873_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2873_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2873_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2873_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2874_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2874_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2874_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2874_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2874_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2875_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2875_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2875_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2875_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2875_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2876_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2876_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2876_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2876_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2876_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2877_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2877_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2877_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2877_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2877_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2878_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2878_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2878_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2878_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2878_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_101_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_101_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_101_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_101_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2879_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2879_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2879_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2879_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2879_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2880_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2880_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2880_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2880_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2880_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2881_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2881_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2881_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2881_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2881_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2882_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2882_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2882_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2882_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2882_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2883_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2883_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2883_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2883_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2883_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2884_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2884_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2884_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2884_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2884_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2885_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2885_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2885_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2885_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2885_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2886_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2886_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2886_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2886_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2886_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2887_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2887_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2887_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2887_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2887_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2888_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2888_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2888_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2888_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2888_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2889_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2889_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2889_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2889_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2889_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2890_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2890_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2890_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2890_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2890_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2891_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2891_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2891_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2891_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2891_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2892_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2892_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2892_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2892_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2892_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2893_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2893_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2893_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2893_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2893_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2894_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2894_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2894_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2894_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2894_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2895_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2895_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2895_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2895_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2895_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2896_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2896_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2896_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2896_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2896_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2897_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2897_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2897_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2897_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2897_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2898_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2898_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2898_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2898_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2898_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2899_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2899_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2899_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2899_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2899_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2900_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2900_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2900_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2900_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2900_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2901_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2901_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2901_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2901_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2901_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2902_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2902_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2902_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2902_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2902_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2903_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2903_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2903_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2903_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2903_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2904_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2904_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2904_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2904_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2904_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2905_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2905_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2905_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2905_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2905_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2906_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2906_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2906_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2906_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2906_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2907_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2907_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2907_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2907_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2907_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2908_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2908_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2908_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2908_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2908_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2909_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2909_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2909_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2909_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2909_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2910_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2910_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2910_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2910_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2910_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2911_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2911_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2911_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2911_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2911_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2912_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2912_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2912_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2912_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2912_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2913_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2913_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2913_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2913_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2913_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2914_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2914_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2914_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2914_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2914_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2915_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2915_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2915_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2915_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2915_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2916_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2916_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2916_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2916_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2916_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2917_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2917_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2917_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2917_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2917_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2918_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2918_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2918_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2918_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2918_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2919_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2919_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2919_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2919_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2919_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2920_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2920_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2920_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2920_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2920_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2921_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2921_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2921_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2921_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2921_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2922_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2922_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2922_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2922_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2922_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2923_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2923_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2923_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2923_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2923_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2924_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2924_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2924_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2924_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2924_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2925_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2925_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2925_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2925_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2925_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2926_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2926_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2926_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2926_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2926_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2927_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2927_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2927_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2927_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2927_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2928_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2928_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2928_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2928_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2928_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2929_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2929_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2929_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2929_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2929_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2930_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2930_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2930_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2930_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2930_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2931_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2931_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2931_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2931_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2931_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2932_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2932_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2932_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2932_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2932_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_102_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_102_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_102_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_102_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2933_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2933_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2933_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2933_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2933_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2934_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2934_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2934_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2934_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2934_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2935_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2935_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2935_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2935_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2935_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2936_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2936_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2936_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2936_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2936_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2937_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2937_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2937_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2937_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2937_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2938_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2938_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2938_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2938_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2938_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2939_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2939_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2939_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2939_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2939_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2940_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2940_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2940_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2940_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2940_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2941_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2941_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2941_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2941_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2941_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2942_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2942_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2942_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2942_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2942_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2943_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2943_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2943_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2943_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2943_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2944_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2944_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2944_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2944_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2944_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2945_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2945_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2945_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2945_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2945_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2946_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2946_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2946_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2946_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2946_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2947_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2947_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2947_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2947_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2947_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2948_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2948_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2948_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2948_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2948_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2949_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2949_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2949_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2949_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2949_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2950_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2950_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2950_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2950_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2950_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2951_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2951_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2951_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2951_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2951_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2952_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2952_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2952_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2952_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2952_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2953_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2953_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2953_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2953_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2953_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2954_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2954_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2954_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2954_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2954_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2955_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2955_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2955_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2955_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2955_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2956_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2956_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2956_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2956_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2956_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2957_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2957_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2957_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2957_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2957_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2958_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2958_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2958_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2958_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2958_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2959_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2959_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2959_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2959_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2959_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2960_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2960_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2960_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2960_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2960_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2961_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2961_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2961_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2961_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2961_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2962_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2962_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2962_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2962_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2962_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2963_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2963_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2963_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2963_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2963_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2964_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2964_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2964_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2964_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2964_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2965_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2965_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2965_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2965_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2965_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2966_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2966_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2966_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2966_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2966_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2967_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2967_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2967_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2967_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2967_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2968_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2968_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2968_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2968_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2968_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2969_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2969_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2969_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2969_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2969_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2970_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2970_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2970_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2970_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2970_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2971_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2971_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2971_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2971_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2971_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2972_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2972_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2972_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2972_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2972_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2973_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2973_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2973_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2973_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2973_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2974_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2974_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2974_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2974_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2974_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2975_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2975_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2975_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2975_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2975_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2976_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2976_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2976_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2976_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2976_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2977_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2977_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2977_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2977_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2977_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2978_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2978_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2978_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2978_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2978_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2979_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2979_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2979_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2979_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2979_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2980_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2980_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2980_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2980_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2980_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2981_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2981_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2981_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2981_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2981_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2982_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2982_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2982_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2982_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2982_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2983_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2983_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2983_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2983_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2983_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2984_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2984_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2984_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2984_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2984_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2985_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2985_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2985_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2985_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2985_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2986_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2986_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2986_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2986_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2986_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_103_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_103_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_103_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_103_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_2987_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2987_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2987_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2987_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2987_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2988_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2988_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2988_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2988_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2988_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2989_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2989_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2989_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2989_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2989_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2990_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2990_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2990_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2990_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2990_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2991_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2991_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2991_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2991_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2991_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2992_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2992_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2992_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2992_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2992_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2993_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2993_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2993_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2993_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2993_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2994_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2994_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2994_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2994_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2994_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2995_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2995_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2995_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2995_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2995_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2996_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2996_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2996_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2996_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2996_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2997_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2997_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2997_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2997_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2997_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2998_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2998_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2998_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2998_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2998_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_2999_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_2999_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_2999_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_2999_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_2999_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3000_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3000_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3000_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3000_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3000_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3001_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3001_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3001_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3001_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3001_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3002_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3002_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3002_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3002_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3002_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3003_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3003_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3003_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3003_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3003_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3004_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3004_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3004_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3004_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3004_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3005_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3005_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3005_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3005_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3005_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3006_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3006_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3006_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3006_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3006_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3007_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3007_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3007_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3007_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3007_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3008_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3008_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3008_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3008_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3008_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3009_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3009_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3009_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3009_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3009_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3010_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3010_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3010_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3010_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3010_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3011_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3011_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3011_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3011_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3011_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3012_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3012_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3012_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3012_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3012_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3013_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3013_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3013_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3013_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3013_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3014_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3014_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3014_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3014_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3014_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3015_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3015_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3015_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3015_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3015_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3016_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3016_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3016_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3016_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3016_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3017_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3017_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3017_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3017_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3017_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3018_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3018_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3018_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3018_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3018_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3019_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3019_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3019_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3019_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3019_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3020_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3020_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3020_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3020_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3020_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3021_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3021_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3021_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3021_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3021_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3022_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3022_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3022_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3022_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3022_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3023_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3023_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3023_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3023_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3023_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3024_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3024_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3024_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3024_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3024_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3025_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3025_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3025_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3025_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3025_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3026_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3026_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3026_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3026_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3026_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_104_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_104_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_104_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_104_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3027_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3027_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3027_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3027_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3027_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3028_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3028_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3028_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3028_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3028_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3029_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3029_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3029_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3029_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3029_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3030_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3030_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3030_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3030_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3030_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3031_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3031_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3031_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3031_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3031_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_105_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_105_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_105_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_105_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3032_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3032_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3032_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3032_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3032_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3033_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3033_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3033_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3033_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3033_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3034_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3034_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3034_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3034_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3034_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3035_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3035_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3035_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3035_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3035_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3036_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3036_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3036_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3036_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3036_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3037_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3037_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3037_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3037_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3037_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3038_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3038_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3038_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3038_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3038_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3039_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3039_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3039_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3039_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3039_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3040_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3040_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3040_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3040_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3040_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3041_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3041_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3041_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3041_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3041_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3042_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3042_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3042_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3042_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3042_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3043_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3043_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3043_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3043_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3043_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3044_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3044_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3044_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3044_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3044_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3045_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3045_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3045_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3045_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3045_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3046_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3046_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3046_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3046_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3046_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3047_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3047_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3047_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3047_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3047_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3048_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3048_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3048_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3048_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3048_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3049_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3049_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3049_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3049_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3049_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3050_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3050_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3050_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3050_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3050_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3051_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3051_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3051_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3051_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3051_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3052_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3052_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3052_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3052_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3052_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3053_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3053_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3053_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3053_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3053_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3054_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3054_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3054_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3054_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3054_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3055_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3055_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3055_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3055_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3055_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3056_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3056_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3056_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3056_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3056_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3057_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3057_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3057_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3057_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3057_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3058_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3058_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3058_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3058_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3058_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3059_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3059_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3059_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3059_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3059_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3060_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3060_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3060_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3060_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3060_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3061_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3061_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3061_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3061_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3061_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3062_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3062_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3062_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3062_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3062_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3063_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3063_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3063_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3063_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3063_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3064_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3064_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3064_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3064_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3064_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3065_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3065_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3065_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3065_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3065_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3066_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3066_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3066_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3066_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3066_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3067_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3067_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3067_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3067_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3067_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3068_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3068_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3068_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3068_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3068_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3069_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3069_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3069_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3069_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3069_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3070_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3070_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3070_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3070_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3070_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3071_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3071_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3071_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3071_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3071_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3072_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3072_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3072_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3072_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3072_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3073_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3073_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3073_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3073_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3073_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3074_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3074_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3074_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3074_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3074_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3075_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3075_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3075_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3075_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3075_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3076_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3076_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3076_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3076_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3076_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_106_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_106_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_106_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_106_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3077_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3077_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3077_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3077_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3077_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3078_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3078_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3078_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3078_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3078_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3079_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3079_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3079_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3079_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3079_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3080_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3080_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3080_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3080_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3080_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3081_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3081_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3081_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3081_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3081_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3082_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3082_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3082_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3082_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3082_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3083_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3083_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3083_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3083_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3083_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3084_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3084_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3084_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3084_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3084_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3085_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3085_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3085_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3085_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3085_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3086_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3086_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3086_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3086_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3086_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3087_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3087_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3087_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3087_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3087_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3088_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3088_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3088_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3088_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3088_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3089_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3089_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3089_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3089_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3089_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3090_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3090_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3090_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3090_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3090_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3091_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3091_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3091_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3091_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3091_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3092_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3092_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3092_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3092_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3092_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3093_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3093_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3093_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3093_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3093_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3094_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3094_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3094_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3094_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3094_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3095_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3095_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3095_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3095_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3095_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3096_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3096_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3096_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3096_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3096_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3097_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3097_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3097_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3097_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3097_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3098_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3098_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3098_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3098_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3098_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3099_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3099_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3099_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3099_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3099_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3100_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3100_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3100_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3100_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3100_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3101_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3101_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3101_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3101_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3101_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3102_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3102_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3102_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3102_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3102_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3103_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3103_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3103_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3103_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3103_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3104_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3104_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3104_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3104_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3104_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3105_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3105_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3105_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3105_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3105_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3106_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3106_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3106_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3106_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3106_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3107_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3107_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3107_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3107_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3107_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3108_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3108_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3108_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3108_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3108_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3109_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3109_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3109_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3109_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3109_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3110_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3110_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3110_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3110_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3110_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3111_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3111_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3111_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3111_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3111_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3112_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3112_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3112_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3112_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3112_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3113_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3113_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3113_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3113_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3113_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3114_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3114_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3114_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3114_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3114_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3115_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3115_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3115_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3115_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3115_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3116_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3116_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3116_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3116_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3116_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3117_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3117_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3117_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3117_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3117_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3118_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3118_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3118_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3118_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3118_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_107_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_107_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_107_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_107_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3119_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3119_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3119_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3119_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3119_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3120_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3120_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3120_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3120_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3120_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3121_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3121_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3121_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3121_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3121_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3122_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3122_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3122_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3122_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3122_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3123_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3123_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3123_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3123_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3123_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3124_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3124_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3124_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3124_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3124_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3125_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3125_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3125_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3125_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3125_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3126_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3126_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3126_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3126_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3126_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3127_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3127_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3127_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3127_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3127_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3128_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3128_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3128_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3128_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3128_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3129_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3129_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3129_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3129_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3129_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3130_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3130_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3130_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3130_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3130_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3131_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3131_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3131_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3131_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3131_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3132_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3132_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3132_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3132_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3132_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3133_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3133_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3133_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3133_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3133_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3134_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3134_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3134_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3134_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3134_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3135_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3135_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3135_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3135_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3135_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3136_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3136_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3136_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3136_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3136_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3137_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3137_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3137_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3137_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3137_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3138_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3138_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3138_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3138_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3138_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3139_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3139_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3139_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3139_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3139_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3140_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3140_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3140_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3140_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3140_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3141_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3141_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3141_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3141_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3141_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3142_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3142_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3142_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3142_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3142_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3143_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3143_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3143_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3143_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3143_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3144_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3144_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3144_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3144_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3144_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3145_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3145_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3145_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3145_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3145_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3146_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3146_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3146_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3146_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3146_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3147_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3147_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3147_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3147_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3147_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3148_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3148_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3148_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3148_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3148_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3149_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3149_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3149_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3149_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3149_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3150_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3150_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3150_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3150_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3150_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3151_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3151_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3151_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3151_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3151_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3152_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3152_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3152_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3152_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3152_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3153_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3153_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3153_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3153_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3153_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3154_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3154_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3154_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3154_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3154_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3155_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3155_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3155_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3155_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3155_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3156_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3156_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3156_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3156_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3156_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3157_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3157_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3157_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3157_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3157_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3158_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3158_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3158_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3158_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3158_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3159_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3159_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3159_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3159_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3159_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3160_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3160_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3160_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3160_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3160_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3161_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3161_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3161_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3161_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3161_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3162_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3162_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3162_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3162_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3162_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3163_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3163_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3163_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3163_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3163_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3164_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3164_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3164_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3164_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3164_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3165_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3165_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3165_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3165_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3165_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3166_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3166_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3166_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3166_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3166_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3167_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3167_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3167_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3167_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3167_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_108_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_108_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_108_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_108_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3168_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3168_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3168_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3168_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3168_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3169_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3169_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3169_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3169_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3169_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_109_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_109_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_109_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_109_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3170_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3170_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3170_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3170_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3170_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3171_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3171_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3171_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3171_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3171_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3172_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3172_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3172_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3172_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3172_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_110_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_110_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_110_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_110_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_111_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_111_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_111_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_111_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3173_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3173_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3173_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3173_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3173_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3174_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3174_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3174_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3174_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3174_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3175_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3175_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3175_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3175_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3175_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_112_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_112_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_112_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_112_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_113_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_113_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_113_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_113_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_114_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_114_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_114_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_114_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_115_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_115_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_115_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_115_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3176_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3176_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3176_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3176_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3176_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_116_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_116_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_116_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_116_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_117_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_117_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_117_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_117_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3177_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3177_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3177_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3177_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3177_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_118_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_118_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_118_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_118_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_119_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_119_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_119_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_119_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3178_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3178_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3178_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3178_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3178_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3179_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3179_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3179_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3179_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3179_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3180_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3180_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3180_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3180_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3180_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3181_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3181_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3181_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3181_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3181_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3182_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3182_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3182_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3182_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3182_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3183_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3183_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3183_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3183_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3183_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3184_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3184_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3184_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3184_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3184_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3185_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3185_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3185_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3185_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3185_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3186_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3186_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3186_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3186_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3186_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3187_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3187_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3187_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3187_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3187_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3188_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3188_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3188_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3188_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3188_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_120_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_120_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_120_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_120_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3189_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3189_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3189_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3189_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3189_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_121_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_121_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_121_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_121_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3190_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3190_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3190_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3190_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3190_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3191_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3191_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3191_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3191_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3191_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3192_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3192_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3192_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3192_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3192_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3193_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3193_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3193_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3193_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3193_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3194_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3194_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3194_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3194_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3194_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3195_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3195_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3195_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3195_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3195_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3196_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3196_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3196_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3196_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3196_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3197_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3197_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3197_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3197_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3197_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3198_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3198_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3198_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3198_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3198_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3199_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3199_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3199_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3199_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3199_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3200_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3200_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3200_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3200_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3200_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3201_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3201_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3201_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3201_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3201_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3202_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3202_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3202_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3202_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3202_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3203_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3203_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3203_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3203_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3203_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3204_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3204_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3204_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3204_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3204_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3205_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3205_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3205_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3205_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3205_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3206_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3206_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3206_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3206_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3206_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3207_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3207_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3207_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3207_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3207_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3208_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3208_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3208_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3208_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3208_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3209_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3209_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3209_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3209_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3209_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3210_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3210_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3210_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3210_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3210_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3211_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3211_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3211_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3211_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3211_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3212_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3212_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3212_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3212_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3212_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3213_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3213_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3213_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3213_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3213_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3214_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3214_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3214_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3214_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3214_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_122_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_122_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_122_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_122_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3215_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3215_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3215_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3215_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3215_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3216_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3216_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3216_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3216_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3216_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_123_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_123_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_123_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_123_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3217_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3217_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3217_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3217_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3217_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3218_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3218_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3218_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3218_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3218_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_124_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_124_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_124_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_124_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3219_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3219_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3219_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3219_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3219_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3220_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3220_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3220_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3220_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3220_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3221_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3221_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3221_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3221_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3221_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3222_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3222_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3222_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3222_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3222_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3223_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3223_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3223_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3223_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3223_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3224_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3224_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3224_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3224_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3224_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3225_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3225_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3225_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3225_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3225_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_125_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_125_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_125_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_125_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3226_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3226_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3226_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3226_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3226_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3227_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3227_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3227_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3227_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3227_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_126_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_126_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_126_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_126_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3228_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3228_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3228_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3228_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3228_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3229_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3229_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3229_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3229_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3229_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3230_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3230_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3230_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3230_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3230_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3231_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3231_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3231_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3231_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3231_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3232_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3232_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3232_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3232_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3232_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3233_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3233_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3233_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3233_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3233_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3234_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3234_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3234_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3234_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3234_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3235_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3235_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3235_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3235_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3235_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3236_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3236_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3236_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3236_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3236_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3237_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3237_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3237_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3237_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3237_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3238_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3238_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3238_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3238_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3238_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3239_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3239_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3239_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3239_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3239_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3240_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3240_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3240_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3240_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3240_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3241_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3241_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3241_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3241_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3241_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3242_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3242_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3242_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3242_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3242_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3243_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3243_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3243_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3243_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3243_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3244_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3244_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3244_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3244_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3244_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3245_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3245_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3245_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3245_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3245_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3246_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3246_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3246_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3246_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3246_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3247_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3247_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3247_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3247_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3247_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3248_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3248_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3248_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3248_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3248_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3249_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3249_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3249_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3249_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3249_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3250_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3250_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3250_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3250_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3250_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3251_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3251_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3251_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3251_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3251_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3252_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3252_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3252_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3252_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3252_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3253_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3253_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3253_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3253_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3253_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3254_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3254_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3254_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3254_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3254_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3255_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3255_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3255_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3255_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3255_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3256_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3256_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3256_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3256_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3256_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3257_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3257_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3257_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3257_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3257_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3258_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3258_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3258_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3258_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3258_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3259_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3259_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3259_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3259_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3259_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3260_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3260_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3260_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3260_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3260_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3261_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3261_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3261_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3261_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3261_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_127_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_127_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_127_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_127_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3262_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3262_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3262_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3262_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3262_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3263_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3263_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3263_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3263_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3263_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3264_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3264_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3264_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3264_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3264_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_128_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_128_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_128_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_128_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3265_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3265_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3265_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3265_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3265_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3266_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3266_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3266_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3266_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3266_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3267_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3267_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3267_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3267_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3267_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_129_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_129_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_129_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_129_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3268_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3268_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3268_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3268_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3268_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3269_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3269_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3269_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3269_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3269_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3270_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3270_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3270_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3270_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3270_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3271_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3271_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3271_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3271_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3271_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3272_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3272_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3272_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3272_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3272_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3273_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3273_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3273_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3273_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3273_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3274_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3274_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3274_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3274_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3274_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3275_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3275_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3275_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3275_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3275_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3276_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3276_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3276_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3276_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3276_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3277_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3277_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3277_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3277_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3277_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3278_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3278_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3278_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3278_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3278_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3279_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3279_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3279_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3279_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3279_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3280_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3280_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3280_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3280_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3280_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3281_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3281_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3281_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3281_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3281_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3282_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3282_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3282_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3282_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3282_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3283_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3283_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3283_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3283_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3283_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3284_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3284_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3284_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3284_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3284_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3285_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3285_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3285_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3285_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3285_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3286_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3286_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3286_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3286_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3286_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3287_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3287_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3287_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3287_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3287_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3288_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3288_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3288_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3288_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3288_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3289_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3289_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3289_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3289_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3289_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3290_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3290_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3290_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3290_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3290_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3291_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3291_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3291_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3291_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3291_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3292_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3292_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3292_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3292_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3292_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3293_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3293_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3293_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3293_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3293_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3294_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3294_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3294_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3294_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3294_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3295_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3295_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3295_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3295_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3295_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3296_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3296_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3296_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3296_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3296_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3297_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3297_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3297_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3297_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3297_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3298_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3298_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3298_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3298_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3298_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3299_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3299_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3299_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3299_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3299_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3300_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3300_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3300_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3300_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3300_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3301_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3301_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3301_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3301_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3301_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3302_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3302_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3302_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3302_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3302_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3303_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3303_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3303_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3303_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3303_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3304_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3304_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3304_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3304_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3304_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3305_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3305_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3305_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3305_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3305_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3306_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3306_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3306_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3306_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3306_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3307_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3307_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3307_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3307_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3307_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_130_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_130_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_130_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_130_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3308_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3308_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3308_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3308_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3308_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3309_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3309_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3309_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3309_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3309_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3310_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3310_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3310_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3310_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3310_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3311_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3311_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3311_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3311_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3311_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3312_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3312_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3312_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3312_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3312_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3313_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3313_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3313_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3313_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3313_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3314_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3314_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3314_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3314_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3314_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3315_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3315_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3315_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3315_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3315_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3316_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3316_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3316_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3316_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3316_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3317_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3317_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3317_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3317_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3317_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3318_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3318_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3318_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3318_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3318_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3319_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3319_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3319_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3319_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3319_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3320_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3320_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3320_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3320_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3320_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3321_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3321_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3321_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3321_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3321_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3322_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3322_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3322_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3322_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3322_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3323_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3323_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3323_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3323_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3323_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3324_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3324_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3324_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3324_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3324_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3325_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3325_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3325_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3325_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3325_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3326_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3326_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3326_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3326_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3326_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3327_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3327_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3327_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3327_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3327_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3328_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3328_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3328_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3328_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3328_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3329_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3329_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3329_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3329_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3329_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3330_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3330_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3330_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3330_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3330_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3331_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3331_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3331_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3331_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3331_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3332_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3332_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3332_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3332_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3332_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3333_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3333_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3333_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3333_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3333_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3334_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3334_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3334_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3334_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3334_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3335_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3335_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3335_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3335_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3335_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3336_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3336_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3336_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3336_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3336_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3337_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3337_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3337_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3337_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3337_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3338_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3338_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3338_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3338_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3338_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3339_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3339_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3339_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3339_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3339_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3340_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3340_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3340_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3340_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3340_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3341_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3341_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3341_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3341_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3341_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3342_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3342_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3342_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3342_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3342_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3343_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3343_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3343_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3343_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3343_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3344_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3344_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3344_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3344_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3344_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3345_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3345_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3345_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3345_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3345_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3346_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3346_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3346_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3346_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3346_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3347_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3347_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3347_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3347_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3347_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3348_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3348_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3348_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3348_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3348_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_131_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_131_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_131_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_131_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3349_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3349_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3349_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3349_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3349_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3350_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3350_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3350_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3350_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3350_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3351_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3351_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3351_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3351_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3351_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3352_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3352_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3352_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3352_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3352_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3353_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3353_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3353_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3353_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3353_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3354_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3354_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3354_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3354_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3354_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3355_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3355_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3355_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3355_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3355_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3356_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3356_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3356_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3356_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3356_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3357_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3357_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3357_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3357_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3357_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3358_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3358_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3358_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3358_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3358_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3359_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3359_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3359_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3359_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3359_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3360_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3360_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3360_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3360_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3360_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3361_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3361_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3361_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3361_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3361_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3362_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3362_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3362_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3362_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3362_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3363_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3363_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3363_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3363_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3363_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3364_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3364_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3364_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3364_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3364_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3365_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3365_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3365_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3365_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3365_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3366_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3366_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3366_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3366_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3366_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3367_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3367_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3367_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3367_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3367_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3368_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3368_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3368_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3368_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3368_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3369_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3369_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3369_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3369_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3369_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3370_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3370_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3370_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3370_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3370_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3371_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3371_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3371_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3371_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3371_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3372_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3372_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3372_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3372_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3372_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3373_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3373_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3373_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3373_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3373_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3374_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3374_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3374_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3374_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3374_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3375_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3375_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3375_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3375_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3375_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3376_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3376_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3376_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3376_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3376_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3377_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3377_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3377_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3377_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3377_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3378_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3378_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3378_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3378_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3378_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3379_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3379_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3379_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3379_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3379_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3380_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3380_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3380_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3380_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3380_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3381_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3381_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3381_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3381_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3381_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3382_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3382_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3382_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3382_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3382_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3383_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3383_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3383_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3383_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3383_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3384_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3384_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3384_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3384_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3384_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3385_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3385_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3385_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3385_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3385_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3386_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3386_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3386_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3386_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3386_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3387_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3387_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3387_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3387_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3387_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3388_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3388_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3388_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3388_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3388_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_132_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_132_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_132_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_132_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3389_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3389_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3389_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3389_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3389_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3390_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3390_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3390_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3390_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3390_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3391_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3391_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3391_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3391_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3391_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3392_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3392_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3392_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3392_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3392_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3393_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3393_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3393_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3393_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3393_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3394_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3394_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3394_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3394_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3394_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3395_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3395_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3395_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3395_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3395_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3396_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3396_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3396_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3396_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3396_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3397_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3397_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3397_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3397_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3397_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3398_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3398_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3398_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3398_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3398_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3399_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3399_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3399_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3399_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3399_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3400_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3400_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3400_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3400_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3400_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3401_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3401_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3401_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3401_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3401_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3402_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3402_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3402_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3402_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3402_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_133_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_133_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_133_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_133_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3403_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3403_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3403_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3403_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3403_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3404_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3404_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3404_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3404_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3404_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3405_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3405_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3405_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3405_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3405_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3406_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3406_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3406_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3406_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3406_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3407_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3407_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3407_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3407_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3407_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3408_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3408_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3408_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3408_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3408_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3409_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3409_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3409_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3409_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3409_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3410_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3410_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3410_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3410_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3410_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3411_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3411_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3411_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3411_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3411_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3412_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3412_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3412_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3412_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3412_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3413_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3413_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3413_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3413_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3413_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3414_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3414_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3414_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3414_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3414_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3415_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3415_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3415_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3415_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3415_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3416_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3416_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3416_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3416_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3416_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3417_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3417_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3417_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3417_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3417_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3418_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3418_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3418_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3418_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3418_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3419_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3419_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3419_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3419_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3419_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3420_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3420_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3420_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3420_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3420_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3421_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3421_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3421_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3421_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3421_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3422_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3422_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3422_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3422_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3422_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3423_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3423_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3423_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3423_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3423_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_134_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_134_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_134_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_134_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3424_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3424_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3424_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3424_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3424_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_135_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_135_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_135_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_135_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3425_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3425_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3425_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3425_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3425_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_136_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_136_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_136_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_136_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3426_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3426_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3426_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3426_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3426_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3427_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3427_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3427_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3427_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3427_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3428_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3428_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3428_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3428_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3428_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3429_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3429_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3429_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3429_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3429_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3430_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3430_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3430_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3430_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3430_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3431_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3431_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3431_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3431_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3431_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3432_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3432_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3432_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3432_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3432_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3433_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3433_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3433_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3433_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3433_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3434_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3434_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3434_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3434_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3434_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_137_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_137_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_137_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_137_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_138_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_138_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_138_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_138_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_139_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_139_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_139_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_139_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_140_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_140_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_140_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_140_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_141_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_141_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_141_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_141_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_142_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_142_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_142_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_142_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_143_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_143_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_143_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_143_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_144_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_144_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_144_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_144_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_145_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_145_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_145_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_145_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_146_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_146_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_146_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_146_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_147_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_147_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_147_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_147_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_148_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_148_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_148_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_148_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_149_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_149_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_149_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_149_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3435_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3435_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3435_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3435_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3435_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_150_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_150_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_150_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_150_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3436_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3436_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3436_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3436_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3436_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3437_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3437_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3437_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3437_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3437_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3438_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3438_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3438_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3438_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3438_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3439_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3439_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3439_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3439_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3439_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3440_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3440_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3440_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3440_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3440_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3441_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3441_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3441_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3441_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3441_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3442_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3442_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3442_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3442_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3442_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3443_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3443_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3443_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3443_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3443_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3444_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3444_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3444_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3444_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3444_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3445_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3445_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3445_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3445_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3445_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3446_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3446_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3446_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3446_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3446_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3447_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3447_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3447_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3447_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3447_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3448_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3448_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3448_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3448_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3448_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3449_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3449_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3449_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3449_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3449_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_151_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_151_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_151_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_151_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_152_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_152_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_152_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_152_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3450_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3450_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3450_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3450_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3450_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3451_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3451_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3451_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3451_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3451_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3452_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3452_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3452_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3452_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3452_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3453_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3453_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3453_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3453_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3453_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3454_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3454_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3454_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3454_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3454_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_153_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_153_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_153_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_153_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3455_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3455_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3455_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3455_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3455_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3456_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3456_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3456_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3456_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3456_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3457_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3457_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3457_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3457_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3457_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3458_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3458_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3458_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3458_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3458_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3459_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3459_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3459_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3459_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3459_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_154_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_154_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_154_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_154_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3460_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3460_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3460_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3460_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3460_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3461_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3461_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3461_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3461_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3461_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3462_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3462_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3462_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3462_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3462_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3463_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3463_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3463_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3463_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3463_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3464_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3464_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3464_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3464_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3464_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3465_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3465_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3465_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3465_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3465_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3466_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3466_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3466_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3466_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3466_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_155_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_155_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_155_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_155_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_156_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_156_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_156_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_156_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_157_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_157_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_157_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_157_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3467_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3467_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3467_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3467_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3467_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3468_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3468_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3468_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3468_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3468_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3469_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3469_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3469_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3469_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3469_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3470_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3470_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3470_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3470_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3470_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3471_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3471_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3471_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3471_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3471_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3472_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3472_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3472_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3472_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3472_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3473_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3473_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3473_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3473_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3473_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3474_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3474_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3474_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3474_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3474_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3475_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3475_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3475_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3475_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3475_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3476_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3476_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3476_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3476_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3476_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3477_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3477_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3477_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3477_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3477_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3478_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3478_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3478_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3478_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3478_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3479_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3479_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3479_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3479_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3479_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3480_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3480_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3480_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3480_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3480_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3481_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3481_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3481_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3481_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3481_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3482_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3482_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3482_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3482_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3482_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3483_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3483_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3483_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3483_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3483_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3484_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3484_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3484_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3484_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3484_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_158_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_158_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_158_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_158_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3485_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3485_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3485_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3485_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3485_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3486_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3486_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3486_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3486_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3486_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3487_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3487_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3487_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3487_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3487_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3488_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3488_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3488_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3488_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3488_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3489_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3489_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3489_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3489_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3489_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3490_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3490_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3490_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3490_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3490_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_159_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_159_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_159_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_159_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3491_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3491_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3491_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3491_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3491_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3492_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3492_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3492_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3492_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3492_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3493_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3493_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3493_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3493_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3493_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3494_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3494_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3494_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3494_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3494_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_160_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_160_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_160_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_160_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3495_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3495_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3495_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3495_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3495_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3496_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3496_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3496_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3496_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3496_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_161_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_161_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_161_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_161_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3497_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3497_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3497_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3497_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3497_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3498_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3498_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3498_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3498_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3498_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3499_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3499_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3499_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3499_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3499_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3500_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3500_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3500_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3500_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3500_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3501_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3501_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3501_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3501_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3501_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3502_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3502_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3502_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3502_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3502_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3503_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3503_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3503_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3503_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3503_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3504_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3504_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3504_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3504_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3504_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_162_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_162_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_162_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_162_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3505_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3505_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3505_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3505_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3505_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3506_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3506_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3506_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3506_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3506_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_163_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_163_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_163_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_163_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3507_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3507_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3507_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3507_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3507_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_164_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_164_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_164_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_164_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_165_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_165_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_165_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_165_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_166_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_166_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_166_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_166_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3508_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3508_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3508_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3508_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3508_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3509_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3509_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3509_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3509_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3509_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3510_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3510_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3510_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3510_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3510_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3511_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3511_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3511_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3511_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3511_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3512_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3512_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3512_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3512_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3512_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3513_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3513_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3513_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3513_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3513_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3514_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3514_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3514_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3514_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3514_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3515_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3515_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3515_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3515_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3515_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3516_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3516_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3516_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3516_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3516_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3517_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3517_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3517_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3517_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3517_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3518_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3518_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3518_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3518_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3518_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3519_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3519_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3519_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3519_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3519_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3520_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3520_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3520_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3520_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3520_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3521_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3521_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3521_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3521_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3521_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3522_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3522_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3522_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3522_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3522_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3523_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3523_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3523_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3523_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3523_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3524_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3524_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3524_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3524_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3524_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3525_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3525_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3525_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3525_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3525_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3526_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3526_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3526_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3526_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3526_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3527_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3527_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3527_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3527_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3527_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3528_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3528_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3528_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3528_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3528_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3529_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3529_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3529_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3529_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3529_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3530_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3530_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3530_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3530_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3530_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3531_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3531_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3531_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3531_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3531_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3532_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3532_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3532_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3532_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3532_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3533_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3533_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3533_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3533_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3533_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3534_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3534_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3534_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3534_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3534_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_167_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_167_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_167_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_167_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3535_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3535_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3535_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3535_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3535_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3536_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3536_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3536_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3536_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3536_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3537_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3537_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3537_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3537_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3537_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3538_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3538_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3538_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3538_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3538_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3539_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3539_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3539_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3539_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3539_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3540_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3540_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3540_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3540_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3540_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3541_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3541_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3541_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3541_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3541_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3542_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3542_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3542_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3542_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3542_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3543_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3543_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3543_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3543_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3543_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3544_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3544_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3544_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3544_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3544_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3545_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3545_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3545_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3545_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3545_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3546_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3546_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3546_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3546_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3546_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3547_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3547_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3547_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3547_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3547_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3548_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3548_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3548_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3548_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3548_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3549_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3549_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3549_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3549_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3549_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3550_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3550_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3550_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3550_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3550_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3551_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3551_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3551_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3551_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3551_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3552_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3552_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3552_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3552_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3552_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3553_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3553_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3553_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3553_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3553_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3554_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3554_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3554_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3554_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3554_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3555_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3555_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3555_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3555_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3555_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3556_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3556_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3556_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3556_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3556_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3557_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3557_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3557_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3557_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3557_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3558_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3558_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3558_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3558_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3558_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3559_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3559_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3559_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3559_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3559_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3560_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3560_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3560_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3560_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3560_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3561_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3561_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3561_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3561_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3561_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3562_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3562_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3562_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3562_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3562_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3563_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3563_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3563_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3563_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3563_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3564_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3564_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3564_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3564_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3564_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3565_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3565_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3565_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3565_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3565_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3566_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3566_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3566_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3566_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3566_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_168_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_168_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_168_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_168_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3567_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3567_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3567_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3567_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3567_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3568_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3568_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3568_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3568_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3568_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3569_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3569_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3569_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3569_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3569_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3570_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3570_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3570_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3570_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3570_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3571_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3571_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3571_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3571_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3571_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3572_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3572_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3572_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3572_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3572_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3573_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3573_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3573_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3573_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3573_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3574_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3574_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3574_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3574_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3574_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3575_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3575_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3575_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3575_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3575_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3576_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3576_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3576_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3576_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3576_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_169_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_169_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_169_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_169_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3577_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3577_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3577_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3577_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3577_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3578_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3578_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3578_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3578_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3578_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_170_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_170_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_170_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_170_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3579_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3579_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3579_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3579_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3579_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3580_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3580_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3580_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3580_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3580_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3581_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3581_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3581_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3581_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3581_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3582_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3582_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3582_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3582_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3582_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3583_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3583_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3583_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3583_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3583_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3584_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3584_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3584_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3584_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3584_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3585_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3585_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3585_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3585_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3585_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3586_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3586_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3586_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3586_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3586_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3587_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3587_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3587_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3587_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3587_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3588_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3588_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3588_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3588_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3588_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3589_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3589_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3589_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3589_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3589_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3590_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3590_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3590_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3590_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3590_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3591_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3591_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3591_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3591_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3591_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3592_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3592_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3592_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3592_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3592_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_171_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_171_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_171_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_171_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3593_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3593_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3593_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3593_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3593_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3594_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3594_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3594_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3594_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3594_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_172_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_172_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_172_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_172_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3595_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3595_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3595_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3595_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3595_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3596_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3596_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3596_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3596_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3596_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3597_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3597_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3597_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3597_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3597_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3598_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3598_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3598_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3598_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3598_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_173_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_173_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_173_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_173_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3599_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3599_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3599_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3599_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3599_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_174_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_174_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_174_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_174_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_175_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_175_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_175_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_175_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3600_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3600_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3600_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3600_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3600_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_176_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_176_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_176_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_176_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_177_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_177_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_177_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_177_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_178_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_178_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_178_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_178_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3601_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3601_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3601_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3601_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3601_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3602_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3602_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3602_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3602_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3602_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3603_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3603_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3603_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3603_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3603_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3604_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3604_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3604_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3604_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3604_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_179_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_179_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_179_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_179_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3605_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3605_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3605_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3605_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3605_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3606_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3606_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3606_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3606_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3606_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3607_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3607_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3607_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3607_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3607_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_180_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_180_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_180_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_180_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3608_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3608_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3608_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3608_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3608_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3609_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3609_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3609_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3609_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3609_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3610_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3610_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3610_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3610_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3610_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3611_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3611_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3611_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3611_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3611_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3612_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3612_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3612_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3612_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3612_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_181_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_181_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_181_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_181_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3613_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3613_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3613_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3613_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3613_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3614_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3614_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3614_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3614_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3614_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3615_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3615_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3615_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3615_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3615_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3616_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3616_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3616_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3616_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3616_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3617_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3617_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3617_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3617_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3617_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3618_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3618_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3618_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3618_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3618_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_182_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_182_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_182_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_182_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_183_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_183_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_183_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_183_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3619_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3619_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3619_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3619_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3619_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3620_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3620_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3620_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3620_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3620_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3621_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3621_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3621_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3621_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3621_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3622_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3622_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3622_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3622_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3622_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_184_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_184_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_184_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_184_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_185_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_185_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_185_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_185_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_186_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_186_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_186_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_186_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3623_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3623_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3623_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3623_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3623_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3624_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3624_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3624_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3624_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3624_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_187_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_187_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_187_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_187_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3625_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3625_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3625_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3625_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3625_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3626_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3626_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3626_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3626_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3626_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_188_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_188_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_188_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_188_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_189_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_189_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_189_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_189_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3627_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3627_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3627_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3627_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3627_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3628_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3628_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3628_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3628_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3628_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3629_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3629_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3629_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3629_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3629_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3630_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3630_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3630_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3630_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3630_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3631_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3631_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3631_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3631_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3631_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_190_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_190_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_190_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_190_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3632_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3632_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3632_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3632_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3632_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3633_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3633_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3633_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3633_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3633_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3634_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3634_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3634_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3634_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3634_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3635_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3635_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3635_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3635_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3635_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3636_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3636_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3636_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3636_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3636_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3637_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3637_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3637_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3637_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3637_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3638_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3638_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3638_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3638_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3638_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3639_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3639_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3639_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3639_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3639_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3640_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3640_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3640_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3640_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3640_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3641_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3641_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3641_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3641_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3641_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_191_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_191_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_191_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_191_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3642_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3642_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3642_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3642_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3642_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3643_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3643_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3643_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3643_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3643_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3644_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3644_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3644_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3644_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3644_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3645_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3645_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3645_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3645_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3645_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3646_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3646_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3646_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3646_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3646_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3647_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3647_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3647_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3647_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3647_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3648_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3648_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3648_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3648_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3648_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3649_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3649_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3649_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3649_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3649_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3650_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3650_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3650_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3650_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3650_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3651_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3651_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3651_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3651_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3651_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_192_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_192_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_192_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_192_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_193_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_193_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_193_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_193_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_194_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_194_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_194_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_194_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3652_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3652_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3652_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3652_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3652_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3653_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3653_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3653_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3653_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3653_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3654_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3654_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3654_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3654_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3654_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3655_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3655_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3655_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3655_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3655_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3656_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3656_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3656_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3656_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3656_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3657_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3657_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3657_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3657_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3657_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3658_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3658_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3658_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3658_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3658_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3659_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3659_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3659_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3659_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3659_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3660_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3660_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3660_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3660_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3660_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_195_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_195_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_195_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_195_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3661_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3661_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3661_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3661_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3661_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3662_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3662_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3662_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3662_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3662_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3663_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3663_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3663_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3663_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3663_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3664_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3664_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3664_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3664_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3664_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3665_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3665_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3665_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3665_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3665_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3666_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3666_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3666_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3666_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3666_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3667_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3667_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3667_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3667_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3667_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3668_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3668_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3668_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3668_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3668_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3669_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3669_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3669_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3669_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3669_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3670_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3670_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3670_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3670_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3670_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3671_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3671_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3671_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3671_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3671_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3672_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3672_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3672_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3672_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3672_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3673_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3673_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3673_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3673_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3673_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3674_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3674_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3674_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3674_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3674_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3675_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3675_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3675_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3675_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3675_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3676_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3676_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3676_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3676_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3676_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3677_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3677_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3677_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3677_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3677_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3678_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3678_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3678_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3678_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3678_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_196_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_196_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_196_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_196_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3679_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3679_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3679_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3679_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3679_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3680_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3680_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3680_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3680_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3680_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3681_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3681_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3681_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3681_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3681_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3682_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3682_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3682_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3682_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3682_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_197_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_197_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_197_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_197_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3683_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3683_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3683_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3683_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3683_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3684_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3684_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3684_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3684_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3684_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3685_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3685_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3685_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3685_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3685_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3686_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3686_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3686_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3686_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3686_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3687_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3687_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3687_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3687_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3687_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3688_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3688_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3688_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3688_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3688_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3689_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3689_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3689_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3689_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3689_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3690_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3690_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3690_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3690_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3690_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3691_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3691_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3691_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3691_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3691_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3692_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3692_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3692_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3692_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3692_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3693_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3693_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3693_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3693_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3693_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3694_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3694_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3694_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3694_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3694_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3695_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3695_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3695_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3695_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3695_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3696_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3696_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3696_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3696_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3696_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3697_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3697_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3697_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3697_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3697_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3698_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3698_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3698_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3698_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3698_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3699_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3699_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3699_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3699_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3699_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3700_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3700_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3700_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3700_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3700_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3701_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3701_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3701_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3701_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3701_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3702_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3702_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3702_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3702_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3702_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_198_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_198_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_198_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_198_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3703_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3703_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3703_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3703_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3703_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3704_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3704_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3704_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3704_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3704_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3705_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3705_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3705_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3705_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3705_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3706_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3706_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3706_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3706_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3706_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_199_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_199_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_199_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_199_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_200_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_200_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_200_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_200_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3707_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3707_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3707_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3707_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3707_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3708_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3708_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3708_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3708_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3708_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3709_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3709_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3709_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3709_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3709_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_201_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_201_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_201_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_201_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3710_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3710_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3710_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3710_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3710_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_202_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_202_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_202_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_202_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_203_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_203_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_203_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_203_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3711_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3711_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3711_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3711_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3711_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_204_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_204_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_204_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_204_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_205_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_205_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_205_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_205_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3712_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3712_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3712_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3712_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3712_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_206_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_206_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_206_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_206_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_207_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_207_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_207_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_207_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_208_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_208_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_208_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_208_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3713_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3713_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3713_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3713_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3713_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_209_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_209_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_209_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_209_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3714_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3714_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3714_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3714_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3714_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_210_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_210_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_210_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_210_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3715_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3715_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3715_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3715_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3715_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3716_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3716_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3716_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3716_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3716_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3717_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3717_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3717_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3717_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3717_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3718_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3718_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3718_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3718_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3718_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3719_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3719_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3719_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3719_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3719_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3720_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3720_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3720_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3720_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3720_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_211_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_211_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_211_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_211_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_212_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_212_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_212_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_212_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_213_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_213_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_213_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_213_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3721_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3721_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3721_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3721_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3721_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3722_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3722_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3722_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3722_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3722_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3723_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3723_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3723_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3723_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3723_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_214_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_214_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_214_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_214_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_215_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_215_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_215_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_215_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3724_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3724_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3724_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3724_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3724_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3725_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3725_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3725_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3725_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3725_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3726_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3726_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3726_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3726_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3726_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3727_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3727_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3727_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3727_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3727_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_216_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_216_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_216_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_216_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_217_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_217_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_217_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_217_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3728_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3728_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3728_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3728_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3728_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3729_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3729_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3729_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3729_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3729_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3730_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3730_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3730_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3730_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3730_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3731_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3731_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3731_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3731_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3731_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3732_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3732_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3732_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3732_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3732_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3733_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3733_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3733_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3733_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3733_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3734_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3734_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3734_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3734_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3734_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3735_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3735_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3735_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3735_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3735_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3736_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3736_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3736_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3736_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3736_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3737_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3737_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3737_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3737_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3737_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3738_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3738_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3738_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3738_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3738_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3739_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3739_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3739_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3739_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3739_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3740_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3740_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3740_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3740_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3740_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3741_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3741_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3741_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3741_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3741_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3742_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3742_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3742_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3742_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3742_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3743_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3743_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3743_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3743_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3743_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_218_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_218_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_218_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_218_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_219_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_219_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_219_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_219_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_220_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_220_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_220_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_220_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3744_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3744_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3744_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3744_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3744_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_221_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_221_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_221_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_221_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3745_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3745_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3745_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3745_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3745_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3746_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3746_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3746_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3746_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3746_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3747_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3747_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3747_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3747_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3747_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3748_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3748_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3748_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3748_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3748_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3749_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3749_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3749_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3749_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3749_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3750_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3750_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3750_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3750_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3750_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3751_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3751_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3751_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3751_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3751_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3752_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3752_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3752_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3752_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3752_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3753_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3753_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3753_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3753_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3753_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3754_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3754_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3754_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3754_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3754_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3755_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3755_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3755_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3755_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3755_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3756_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3756_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3756_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3756_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3756_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3757_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3757_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3757_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3757_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3757_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3758_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3758_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3758_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3758_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3758_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3759_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3759_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3759_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3759_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3759_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3760_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3760_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3760_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3760_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3760_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3761_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3761_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3761_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3761_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3761_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3762_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3762_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3762_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3762_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3762_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3763_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3763_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3763_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3763_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3763_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3764_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3764_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3764_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3764_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3764_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3765_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3765_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3765_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3765_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3765_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3766_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3766_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3766_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3766_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3766_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3767_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3767_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3767_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3767_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3767_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3768_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3768_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3768_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3768_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3768_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_222_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_222_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_222_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_222_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3769_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3769_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3769_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3769_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3769_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3770_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3770_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3770_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3770_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3770_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3771_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3771_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3771_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3771_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3771_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3772_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3772_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3772_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3772_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3772_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_223_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_223_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_223_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_223_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3773_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3773_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3773_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3773_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3773_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_224_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_224_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_224_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_224_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3774_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3774_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3774_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3774_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3774_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_225_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_225_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_225_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_225_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3775_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3775_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3775_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3775_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3775_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3776_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3776_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3776_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3776_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3776_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_226_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_226_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_226_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_226_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3777_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3777_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3777_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3777_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3777_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3778_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3778_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3778_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3778_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3778_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3779_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3779_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3779_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3779_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3779_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3780_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3780_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3780_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3780_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3780_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3781_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3781_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3781_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3781_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3781_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_227_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_227_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_227_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_227_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3782_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3782_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3782_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3782_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3782_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_228_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_228_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_228_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_228_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_229_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_229_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_229_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_229_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3783_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3783_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3783_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3783_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3783_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3784_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3784_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3784_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3784_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3784_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3785_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3785_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3785_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3785_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3785_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3786_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3786_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3786_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3786_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3786_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_230_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_230_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_230_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_230_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3787_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3787_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3787_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3787_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3787_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_231_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_231_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_231_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_231_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3788_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3788_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3788_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3788_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3788_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3789_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3789_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3789_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3789_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3789_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3790_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3790_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3790_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3790_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3790_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_232_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_232_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_232_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_232_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3791_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3791_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3791_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3791_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3791_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3792_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3792_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3792_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3792_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3792_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3793_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3793_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3793_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3793_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3793_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_233_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_233_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_233_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_233_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3794_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3794_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3794_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3794_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3794_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_234_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_234_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_234_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_234_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3795_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3795_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3795_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3795_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3795_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3796_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3796_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3796_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3796_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3796_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_235_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_235_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_235_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_235_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3797_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3797_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3797_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3797_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3797_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3798_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3798_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3798_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3798_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3798_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3799_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3799_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3799_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3799_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3799_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3800_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3800_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3800_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3800_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3800_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3801_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3801_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3801_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3801_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3801_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3802_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3802_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3802_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3802_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3802_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3803_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3803_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3803_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3803_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3803_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3804_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3804_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3804_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3804_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3804_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3805_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3805_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3805_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3805_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3805_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3806_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3806_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3806_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3806_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3806_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3807_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3807_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3807_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3807_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3807_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3808_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3808_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3808_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3808_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3808_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3809_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3809_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3809_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3809_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3809_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3810_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3810_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3810_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3810_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3810_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3811_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3811_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3811_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3811_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3811_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_236_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_236_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_236_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_236_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_237_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_237_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_237_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_237_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_238_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_238_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_238_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_238_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3812_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3812_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3812_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3812_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3812_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3813_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3813_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3813_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3813_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3813_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3814_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3814_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3814_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3814_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3814_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3815_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3815_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3815_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3815_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3815_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_239_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_239_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_239_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_239_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3816_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3816_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3816_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3816_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3816_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3817_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3817_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3817_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3817_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3817_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3818_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3818_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3818_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3818_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3818_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3819_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3819_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3819_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3819_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3819_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3820_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3820_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3820_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3820_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3820_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3821_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3821_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3821_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3821_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3821_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3822_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3822_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3822_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3822_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3822_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_240_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_240_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_240_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_240_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3823_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3823_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3823_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3823_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3823_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3824_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3824_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3824_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3824_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3824_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_241_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_241_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_241_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_241_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3825_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3825_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3825_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3825_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3825_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3826_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3826_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3826_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3826_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3826_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3827_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3827_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3827_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3827_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3827_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_242_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_242_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_242_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_242_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3828_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3828_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3828_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3828_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3828_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3829_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3829_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3829_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3829_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3829_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_243_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_243_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_243_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_243_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3830_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3830_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3830_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3830_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3830_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_244_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_244_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_244_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_244_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3831_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3831_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3831_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3831_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3831_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_245_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_245_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_245_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_245_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_246_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_246_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_246_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_246_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_247_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_247_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_247_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_247_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3832_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3832_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3832_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3832_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3832_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3833_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3833_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3833_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3833_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3833_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_248_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_248_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_248_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_248_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3834_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3834_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3834_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3834_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3834_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3835_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3835_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3835_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3835_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3835_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3836_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3836_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3836_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3836_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3836_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3837_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3837_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3837_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3837_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3837_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3838_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3838_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3838_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3838_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3838_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_249_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_249_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_249_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_249_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3839_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3839_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3839_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3839_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3839_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3840_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3840_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3840_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3840_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3840_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3841_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3841_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3841_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3841_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3841_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_250_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_250_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_250_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_250_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3842_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3842_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3842_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3842_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3842_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3843_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3843_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3843_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3843_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3843_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3844_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3844_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3844_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3844_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3844_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_251_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_251_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_251_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_251_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_252_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_252_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_252_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_252_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3845_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3845_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3845_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3845_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3845_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_253_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_253_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_253_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_253_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3846_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3846_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3846_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3846_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3846_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3847_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3847_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3847_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3847_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3847_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_254_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_254_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_254_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_254_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3848_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3848_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3848_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3848_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3848_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3849_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3849_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3849_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3849_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3849_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_255_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_255_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_255_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_255_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_256_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_256_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_256_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_256_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3850_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3850_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3850_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3850_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3850_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3851_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3851_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3851_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3851_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3851_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3852_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3852_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3852_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3852_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3852_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_257_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_257_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_257_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_257_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_258_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_258_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_258_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_258_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_259_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_259_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_259_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_259_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_260_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_260_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_260_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_260_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_261_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_261_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_261_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_261_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3853_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3853_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3853_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3853_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3853_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3854_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3854_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3854_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3854_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3854_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3855_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3855_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3855_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3855_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3855_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3856_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3856_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3856_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3856_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3856_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3857_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3857_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3857_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3857_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3857_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3858_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3858_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3858_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3858_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3858_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3859_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3859_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3859_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3859_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3859_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3860_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3860_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3860_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3860_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3860_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3861_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3861_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3861_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3861_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3861_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3862_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3862_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3862_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3862_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3862_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_262_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_262_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_262_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_262_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3863_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3863_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3863_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3863_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3863_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3864_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3864_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3864_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3864_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3864_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3865_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3865_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3865_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3865_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3865_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_263_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_263_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_263_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_263_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3866_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3866_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3866_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3866_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3866_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3867_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3867_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3867_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3867_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3867_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3868_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3868_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3868_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3868_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3868_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_264_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_264_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_264_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_264_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_265_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_265_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_265_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_265_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_266_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_266_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_266_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_266_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3869_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3869_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3869_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3869_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3869_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3870_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3870_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3870_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3870_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3870_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3871_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3871_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3871_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3871_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3871_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_267_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_267_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_267_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_267_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3872_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3872_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3872_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3872_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3872_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3873_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3873_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3873_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3873_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3873_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_268_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_268_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_268_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_268_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_269_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_269_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_269_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_269_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3874_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3874_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3874_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3874_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3874_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3875_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3875_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3875_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3875_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3875_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3876_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3876_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3876_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3876_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3876_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_270_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_270_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_270_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_270_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3877_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3877_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3877_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3877_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3877_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_271_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_271_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_271_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_271_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3878_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3878_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3878_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3878_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3878_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3879_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3879_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3879_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3879_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3879_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_272_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_272_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_272_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_272_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3880_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3880_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3880_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3880_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3880_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3881_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3881_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3881_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3881_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3881_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3882_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3882_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3882_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3882_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3882_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_273_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_273_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_273_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_273_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3883_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3883_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3883_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3883_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3883_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3884_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3884_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3884_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3884_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3884_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3885_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3885_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3885_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3885_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3885_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3886_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3886_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3886_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3886_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3886_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3887_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3887_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3887_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3887_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3887_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3888_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3888_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3888_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3888_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3888_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_274_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_274_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_274_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_274_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_275_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_275_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_275_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_275_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3889_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3889_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3889_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3889_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3889_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3890_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3890_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3890_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3890_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3890_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3891_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3891_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3891_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3891_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3891_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_276_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_276_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_276_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_276_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3892_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3892_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3892_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3892_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3892_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_277_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_277_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_277_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_277_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_278_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_278_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_278_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_278_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_279_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_279_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_279_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_279_io_co; // @[wallace.scala 57:25]
  wire  HalfAdder_280_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_280_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_280_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_280_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3893_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3893_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3893_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3893_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3893_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3894_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3894_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3894_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3894_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3894_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_281_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_281_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_281_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_281_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3895_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3895_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3895_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3895_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3895_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3896_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3896_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3896_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3896_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3896_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_282_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_282_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_282_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_282_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3897_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3897_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3897_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3897_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3897_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3898_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3898_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3898_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3898_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3898_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_283_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_283_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_283_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_283_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3899_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3899_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3899_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3899_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3899_io_co; // @[wallace.scala 67:25]
  wire  HalfAdder_284_io_a; // @[wallace.scala 57:25]
  wire  HalfAdder_284_io_b; // @[wallace.scala 57:25]
  wire  HalfAdder_284_io_s; // @[wallace.scala 57:25]
  wire  HalfAdder_284_io_co; // @[wallace.scala 57:25]
  wire  FullAdder_3900_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3900_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3900_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3900_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3900_io_co; // @[wallace.scala 67:25]
  wire  FullAdder_3901_io_a; // @[wallace.scala 67:25]
  wire  FullAdder_3901_io_b; // @[wallace.scala 67:25]
  wire  FullAdder_3901_io_ci; // @[wallace.scala 67:25]
  wire  FullAdder_3901_io_s; // @[wallace.scala 67:25]
  wire  FullAdder_3901_io_co; // @[wallace.scala 67:25]
  wire  res0_0 = io_pp_0[0]; // @[wallace.scala 34:43]
  wire  res0_1 = io_pp_0[1]; // @[wallace.scala 34:43]
  wire  res1_1 = io_pp_1[0]; // @[wallace.scala 34:43]
  wire  res0_126 = HalfAdder_283_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_125 = HalfAdder_281_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_124 = FullAdder_3886_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_123 = HalfAdder_265_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_122 = FullAdder_3834_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_121 = HalfAdder_229_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_120 = HalfAdder_205_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_119 = FullAdder_3601_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_118 = HalfAdder_149_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_117 = FullAdder_3435_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [9:0] _T_4104 = {res0_126,res0_125,res0_124,res0_123,res0_122,res0_121,res0_120,res0_119,res0_118,res0_117}; // @[Cat.scala 29:58]
  wire  res0_116 = FullAdder_3602_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_115 = FullAdder_3835_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_114 = FullAdder_3783_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_113 = FullAdder_3712_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_112 = FullAdder_3836_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_111 = FullAdder_3784_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_110 = HalfAdder_206_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_109 = FullAdder_3785_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_108 = HalfAdder_207_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [18:0] _T_4113 = {_T_4104,res0_116,res0_115,res0_114,res0_113,res0_112,res0_111,res0_110,res0_109,res0_108}; // @[Cat.scala 29:58]
  wire  res0_107 = FullAdder_3786_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_106 = HalfAdder_230_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_105 = FullAdder_3887_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_104 = HalfAdder_266_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_103 = FullAdder_3837_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_102 = FullAdder_3787_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_101 = FullAdder_3838_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_100 = HalfAdder_249_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_99 = FullAdder_3839_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [27:0] _T_4122 = {_T_4113,res0_107,res0_106,res0_105,res0_104,res0_103,res0_102,res0_101,res0_100,res0_99}; // @[Cat.scala 29:58]
  wire  res0_98 = FullAdder_3788_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_97 = FullAdder_3869_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_96 = FullAdder_3840_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_95 = FullAdder_3870_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_94 = FullAdder_3841_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_93 = HalfAdder_250_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_92 = FullAdder_3842_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_91 = FullAdder_3871_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_90 = FullAdder_3895_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [36:0] _T_4131 = {_T_4122,res0_98,res0_97,res0_96,res0_95,res0_94,res0_93,res0_92,res0_91,res0_90}; // @[Cat.scala 29:58]
  wire  res0_89 = FullAdder_3888_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_88 = HalfAdder_267_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_87 = FullAdder_3872_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_86 = HalfAdder_274_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_85 = FullAdder_3896_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_84 = HalfAdder_275_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_83 = HalfAdder_269_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_82 = FullAdder_3874_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_81 = FullAdder_3846_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [45:0] _T_4140 = {_T_4131,res0_89,res0_88,res0_87,res0_86,res0_85,res0_84,res0_83,res0_82,res0_81}; // @[Cat.scala 29:58]
  wire  res0_80 = FullAdder_3847_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_79 = HalfAdder_254_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_78 = FullAdder_3889_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_77 = FullAdder_3875_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_76 = FullAdder_3848_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_75 = FullAdder_3849_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_74 = HalfAdder_255_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_73 = HalfAdder_256_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_72 = FullAdder_3890_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [54:0] _T_4149 = {_T_4140,res0_80,res0_79,res0_78,res0_77,res0_76,res0_75,res0_74,res0_73,res0_72}; // @[Cat.scala 29:58]
  wire  res0_71 = FullAdder_3901_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_70 = FullAdder_3899_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_69 = HalfAdder_284_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_68 = FullAdder_3892_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_67 = HalfAdder_277_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_66 = HalfAdder_278_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_65 = FullAdder_3878_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_64 = FullAdder_3900_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_63 = FullAdder_3897_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [63:0] _T_4158 = {_T_4149,res0_71,res0_70,res0_69,res0_68,res0_67,res0_66,res0_65,res0_64,res0_63}; // @[Cat.scala 29:58]
  wire  res0_62 = HalfAdder_279_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_61 = FullAdder_3880_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_60 = FullAdder_3853_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_59 = FullAdder_3818_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_58 = FullAdder_3854_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_57 = FullAdder_3881_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_56 = FullAdder_3855_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_55 = FullAdder_3856_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_54 = FullAdder_3821_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [72:0] _T_4167 = {_T_4158,res0_62,res0_61,res0_60,res0_59,res0_58,res0_57,res0_56,res0_55,res0_54}; // @[Cat.scala 29:58]
  wire  res0_53 = FullAdder_3857_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_52 = FullAdder_3858_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_51 = FullAdder_3882_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_50 = FullAdder_3859_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_49 = FullAdder_3824_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_48 = FullAdder_3860_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_47 = HalfAdder_241_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_46 = FullAdder_3825_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_45 = FullAdder_3826_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [81:0] _T_4176 = {_T_4167,res0_53,res0_52,res0_51,res0_50,res0_49,res0_48,res0_47,res0_46,res0_45}; // @[Cat.scala 29:58]
  wire  res0_44 = FullAdder_3861_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_43 = FullAdder_3827_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_42 = FullAdder_3862_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_41 = HalfAdder_262_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_40 = FullAdder_3863_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_39 = FullAdder_3828_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_38 = FullAdder_3829_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_37 = FullAdder_3864_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_36 = HalfAdder_273_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [90:0] _T_4185 = {_T_4176,res0_44,res0_43,res0_42,res0_41,res0_40,res0_39,res0_38,res0_37,res0_36}; // @[Cat.scala 29:58]
  wire  res0_35 = FullAdder_3865_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_34 = FullAdder_3830_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_33 = HalfAdder_244_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_32 = FullAdder_3774_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_31 = FullAdder_3831_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_30 = HalfAdder_263_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_29 = HalfAdder_280_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_28 = FullAdder_3883_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_27 = FullAdder_3866_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [99:0] _T_4194 = {_T_4185,res0_35,res0_34,res0_33,res0_32,res0_31,res0_30,res0_29,res0_28,res0_27}; // @[Cat.scala 29:58]
  wire  res0_26 = HalfAdder_246_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_25 = FullAdder_3777_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_24 = FullAdder_3898_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_23 = FullAdder_3893_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_22 = FullAdder_3884_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_21 = FullAdder_3867_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_20 = HalfAdder_247_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_19 = FullAdder_3778_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_18 = FullAdder_3707_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [108:0] _T_4203 = {_T_4194,res0_26,res0_25,res0_24,res0_23,res0_22,res0_21,res0_20,res0_19,res0_18}; // @[Cat.scala 29:58]
  wire  res0_17 = FullAdder_3708_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_16 = FullAdder_3894_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_15 = FullAdder_3885_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_14 = FullAdder_3868_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_13 = FullAdder_3832_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_12 = FullAdder_3779_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_11 = FullAdder_3780_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_10 = HalfAdder_201_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_9 = FullAdder_3599_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [117:0] _T_4212 = {_T_4203,res0_17,res0_16,res0_15,res0_14,res0_13,res0_12,res0_11,res0_10,res0_9}; // @[Cat.scala 29:58]
  wire  res0_8 = FullAdder_3833_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_7 = FullAdder_3781_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_6 = FullAdder_3710_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_5 = HalfAdder_174_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_4 = HalfAdder_143_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_3 = HalfAdder_91_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire  res0_2 = HalfAdder_65_io_s; // @[wallace.scala 78:49 wallace.scala 83:13]
  wire [126:0] _T_4221 = {_T_4212,res0_8,res0_7,res0_6,res0_5,res0_4,res0_3,res0_2,res0_1,res0_0}; // @[Cat.scala 29:58]
  wire  res1_118 = FullAdder_3435_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_117 = FullAdder_3602_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_116 = FullAdder_3835_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_113 = FullAdder_3836_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_110 = FullAdder_3785_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [16:0] _T_4237 = {8'h0,res1_118,res1_117,res1_116,1'h0,1'h0,res1_113,1'h0,1'h0,res1_110}; // @[Cat.scala 29:58]
  wire  res1_108 = FullAdder_3786_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_107 = HalfAdder_230_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_106 = FullAdder_3887_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_102 = FullAdder_3838_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_101 = HalfAdder_249_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [25:0] _T_4246 = {_T_4237,1'h0,res1_108,res1_107,res1_106,1'h0,1'h0,1'h0,res1_102,res1_101}; // @[Cat.scala 29:58]
  wire  res1_100 = FullAdder_3839_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_98 = FullAdder_3869_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_96 = FullAdder_3870_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_94 = HalfAdder_250_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_93 = FullAdder_3842_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_92 = FullAdder_3871_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [34:0] _T_4255 = {_T_4246,res1_100,1'h0,res1_98,1'h0,res1_96,1'h0,res1_94,res1_93,res1_92}; // @[Cat.scala 29:58]
  wire  res1_91 = FullAdder_3895_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_88 = FullAdder_3872_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_87 = HalfAdder_274_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_86 = FullAdder_3896_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_83 = FullAdder_3874_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [43:0] _T_4264 = {_T_4255,res1_91,1'h0,1'h0,res1_88,res1_87,res1_86,1'h0,1'h0,res1_83}; // @[Cat.scala 29:58]
  wire  res1_81 = FullAdder_3847_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_80 = HalfAdder_254_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_79 = FullAdder_3889_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_76 = FullAdder_3849_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_75 = HalfAdder_255_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_74 = HalfAdder_256_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [52:0] _T_4273 = {_T_4264,1'h0,res1_81,res1_80,res1_79,1'h0,1'h0,res1_76,res1_75,res1_74}; // @[Cat.scala 29:58]
  wire  res1_73 = FullAdder_3890_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_72 = FullAdder_3901_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_70 = HalfAdder_284_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_68 = HalfAdder_277_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_67 = HalfAdder_278_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_65 = FullAdder_3900_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [61:0] _T_4282 = {_T_4273,res1_73,res1_72,1'h0,res1_70,1'h0,res1_68,res1_67,1'h0,res1_65}; // @[Cat.scala 29:58]
  wire  res1_59 = FullAdder_3854_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_58 = FullAdder_3881_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_56 = FullAdder_3856_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [70:0] _T_4291 = {_T_4282,1'h0,1'h0,1'h0,1'h0,1'h0,res1_59,res1_58,1'h0,res1_56}; // @[Cat.scala 29:58]
  wire  res1_54 = FullAdder_3857_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_53 = FullAdder_3858_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_52 = FullAdder_3882_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_49 = FullAdder_3860_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_47 = FullAdder_3825_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [79:0] _T_4300 = {_T_4291,1'h0,res1_54,res1_53,res1_52,1'h0,1'h0,res1_49,1'h0,res1_47}; // @[Cat.scala 29:58]
  wire  res1_46 = FullAdder_3826_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_45 = FullAdder_3861_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_43 = FullAdder_3862_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_42 = HalfAdder_262_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_41 = FullAdder_3863_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_39 = FullAdder_3829_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_38 = FullAdder_3864_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [88:0] _T_4309 = {_T_4300,res1_46,res1_45,1'h0,res1_43,res1_42,res1_41,1'h0,res1_39,res1_38}; // @[Cat.scala 29:58]
  wire  res1_37 = HalfAdder_273_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_34 = HalfAdder_244_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_32 = FullAdder_3831_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_31 = HalfAdder_263_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_30 = HalfAdder_280_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [97:0] _T_4318 = {_T_4309,res1_37,1'h0,1'h0,res1_34,1'h0,res1_32,res1_31,res1_30,1'h0}; // @[Cat.scala 29:58]
  wire  res1_25 = FullAdder_3898_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [106:0] _T_4327 = {_T_4318,1'h0,1'h0,1'h0,res1_25,1'h0,1'h0,1'h0,1'h0,1'h0}; // @[Cat.scala 29:58]
  wire  res1_18 = FullAdder_3708_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_17 = FullAdder_3894_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire  res1_12 = FullAdder_3780_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [115:0] _T_4336 = {_T_4327,1'h0,res1_18,res1_17,1'h0,1'h0,1'h0,1'h0,res1_12,1'h0}; // @[Cat.scala 29:58]
  wire  res1_9 = FullAdder_3833_io_co; // @[wallace.scala 79:49 wallace.scala 87:15]
  wire [124:0] _T_4345 = {_T_4336,1'h0,res1_9,1'h0,1'h0,1'h0,1'h0,1'h0,1'h0,1'h0}; // @[Cat.scala 29:58]
  wire [126:0] _T_4347 = {_T_4345,res1_1,1'h0}; // @[Cat.scala 29:58]
  HalfAdder HalfAdder ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_io_a),
    .io_b(HalfAdder_io_b),
    .io_s(HalfAdder_io_s),
    .io_co(HalfAdder_io_co)
  );
  FullAdder FullAdder ( // @[wallace.scala 67:25]
    .io_a(FullAdder_io_a),
    .io_b(FullAdder_io_b),
    .io_ci(FullAdder_io_ci),
    .io_s(FullAdder_io_s),
    .io_co(FullAdder_io_co)
  );
  FullAdder FullAdder_1 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1_io_a),
    .io_b(FullAdder_1_io_b),
    .io_ci(FullAdder_1_io_ci),
    .io_s(FullAdder_1_io_s),
    .io_co(FullAdder_1_io_co)
  );
  FullAdder FullAdder_2 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2_io_a),
    .io_b(FullAdder_2_io_b),
    .io_ci(FullAdder_2_io_ci),
    .io_s(FullAdder_2_io_s),
    .io_co(FullAdder_2_io_co)
  );
  HalfAdder HalfAdder_1 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_1_io_a),
    .io_b(HalfAdder_1_io_b),
    .io_s(HalfAdder_1_io_s),
    .io_co(HalfAdder_1_io_co)
  );
  FullAdder FullAdder_3 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3_io_a),
    .io_b(FullAdder_3_io_b),
    .io_ci(FullAdder_3_io_ci),
    .io_s(FullAdder_3_io_s),
    .io_co(FullAdder_3_io_co)
  );
  FullAdder FullAdder_4 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_4_io_a),
    .io_b(FullAdder_4_io_b),
    .io_ci(FullAdder_4_io_ci),
    .io_s(FullAdder_4_io_s),
    .io_co(FullAdder_4_io_co)
  );
  FullAdder FullAdder_5 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_5_io_a),
    .io_b(FullAdder_5_io_b),
    .io_ci(FullAdder_5_io_ci),
    .io_s(FullAdder_5_io_s),
    .io_co(FullAdder_5_io_co)
  );
  FullAdder FullAdder_6 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_6_io_a),
    .io_b(FullAdder_6_io_b),
    .io_ci(FullAdder_6_io_ci),
    .io_s(FullAdder_6_io_s),
    .io_co(FullAdder_6_io_co)
  );
  FullAdder FullAdder_7 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_7_io_a),
    .io_b(FullAdder_7_io_b),
    .io_ci(FullAdder_7_io_ci),
    .io_s(FullAdder_7_io_s),
    .io_co(FullAdder_7_io_co)
  );
  FullAdder FullAdder_8 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_8_io_a),
    .io_b(FullAdder_8_io_b),
    .io_ci(FullAdder_8_io_ci),
    .io_s(FullAdder_8_io_s),
    .io_co(FullAdder_8_io_co)
  );
  HalfAdder HalfAdder_2 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_2_io_a),
    .io_b(HalfAdder_2_io_b),
    .io_s(HalfAdder_2_io_s),
    .io_co(HalfAdder_2_io_co)
  );
  FullAdder FullAdder_9 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_9_io_a),
    .io_b(FullAdder_9_io_b),
    .io_ci(FullAdder_9_io_ci),
    .io_s(FullAdder_9_io_s),
    .io_co(FullAdder_9_io_co)
  );
  FullAdder FullAdder_10 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_10_io_a),
    .io_b(FullAdder_10_io_b),
    .io_ci(FullAdder_10_io_ci),
    .io_s(FullAdder_10_io_s),
    .io_co(FullAdder_10_io_co)
  );
  FullAdder FullAdder_11 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_11_io_a),
    .io_b(FullAdder_11_io_b),
    .io_ci(FullAdder_11_io_ci),
    .io_s(FullAdder_11_io_s),
    .io_co(FullAdder_11_io_co)
  );
  FullAdder FullAdder_12 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_12_io_a),
    .io_b(FullAdder_12_io_b),
    .io_ci(FullAdder_12_io_ci),
    .io_s(FullAdder_12_io_s),
    .io_co(FullAdder_12_io_co)
  );
  FullAdder FullAdder_13 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_13_io_a),
    .io_b(FullAdder_13_io_b),
    .io_ci(FullAdder_13_io_ci),
    .io_s(FullAdder_13_io_s),
    .io_co(FullAdder_13_io_co)
  );
  FullAdder FullAdder_14 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_14_io_a),
    .io_b(FullAdder_14_io_b),
    .io_ci(FullAdder_14_io_ci),
    .io_s(FullAdder_14_io_s),
    .io_co(FullAdder_14_io_co)
  );
  FullAdder FullAdder_15 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_15_io_a),
    .io_b(FullAdder_15_io_b),
    .io_ci(FullAdder_15_io_ci),
    .io_s(FullAdder_15_io_s),
    .io_co(FullAdder_15_io_co)
  );
  FullAdder FullAdder_16 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_16_io_a),
    .io_b(FullAdder_16_io_b),
    .io_ci(FullAdder_16_io_ci),
    .io_s(FullAdder_16_io_s),
    .io_co(FullAdder_16_io_co)
  );
  FullAdder FullAdder_17 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_17_io_a),
    .io_b(FullAdder_17_io_b),
    .io_ci(FullAdder_17_io_ci),
    .io_s(FullAdder_17_io_s),
    .io_co(FullAdder_17_io_co)
  );
  HalfAdder HalfAdder_3 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_3_io_a),
    .io_b(HalfAdder_3_io_b),
    .io_s(HalfAdder_3_io_s),
    .io_co(HalfAdder_3_io_co)
  );
  FullAdder FullAdder_18 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_18_io_a),
    .io_b(FullAdder_18_io_b),
    .io_ci(FullAdder_18_io_ci),
    .io_s(FullAdder_18_io_s),
    .io_co(FullAdder_18_io_co)
  );
  FullAdder FullAdder_19 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_19_io_a),
    .io_b(FullAdder_19_io_b),
    .io_ci(FullAdder_19_io_ci),
    .io_s(FullAdder_19_io_s),
    .io_co(FullAdder_19_io_co)
  );
  FullAdder FullAdder_20 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_20_io_a),
    .io_b(FullAdder_20_io_b),
    .io_ci(FullAdder_20_io_ci),
    .io_s(FullAdder_20_io_s),
    .io_co(FullAdder_20_io_co)
  );
  FullAdder FullAdder_21 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_21_io_a),
    .io_b(FullAdder_21_io_b),
    .io_ci(FullAdder_21_io_ci),
    .io_s(FullAdder_21_io_s),
    .io_co(FullAdder_21_io_co)
  );
  FullAdder FullAdder_22 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_22_io_a),
    .io_b(FullAdder_22_io_b),
    .io_ci(FullAdder_22_io_ci),
    .io_s(FullAdder_22_io_s),
    .io_co(FullAdder_22_io_co)
  );
  FullAdder FullAdder_23 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_23_io_a),
    .io_b(FullAdder_23_io_b),
    .io_ci(FullAdder_23_io_ci),
    .io_s(FullAdder_23_io_s),
    .io_co(FullAdder_23_io_co)
  );
  FullAdder FullAdder_24 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_24_io_a),
    .io_b(FullAdder_24_io_b),
    .io_ci(FullAdder_24_io_ci),
    .io_s(FullAdder_24_io_s),
    .io_co(FullAdder_24_io_co)
  );
  FullAdder FullAdder_25 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_25_io_a),
    .io_b(FullAdder_25_io_b),
    .io_ci(FullAdder_25_io_ci),
    .io_s(FullAdder_25_io_s),
    .io_co(FullAdder_25_io_co)
  );
  FullAdder FullAdder_26 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_26_io_a),
    .io_b(FullAdder_26_io_b),
    .io_ci(FullAdder_26_io_ci),
    .io_s(FullAdder_26_io_s),
    .io_co(FullAdder_26_io_co)
  );
  FullAdder FullAdder_27 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_27_io_a),
    .io_b(FullAdder_27_io_b),
    .io_ci(FullAdder_27_io_ci),
    .io_s(FullAdder_27_io_s),
    .io_co(FullAdder_27_io_co)
  );
  FullAdder FullAdder_28 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_28_io_a),
    .io_b(FullAdder_28_io_b),
    .io_ci(FullAdder_28_io_ci),
    .io_s(FullAdder_28_io_s),
    .io_co(FullAdder_28_io_co)
  );
  FullAdder FullAdder_29 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_29_io_a),
    .io_b(FullAdder_29_io_b),
    .io_ci(FullAdder_29_io_ci),
    .io_s(FullAdder_29_io_s),
    .io_co(FullAdder_29_io_co)
  );
  FullAdder FullAdder_30 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_30_io_a),
    .io_b(FullAdder_30_io_b),
    .io_ci(FullAdder_30_io_ci),
    .io_s(FullAdder_30_io_s),
    .io_co(FullAdder_30_io_co)
  );
  FullAdder FullAdder_31 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_31_io_a),
    .io_b(FullAdder_31_io_b),
    .io_ci(FullAdder_31_io_ci),
    .io_s(FullAdder_31_io_s),
    .io_co(FullAdder_31_io_co)
  );
  FullAdder FullAdder_32 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_32_io_a),
    .io_b(FullAdder_32_io_b),
    .io_ci(FullAdder_32_io_ci),
    .io_s(FullAdder_32_io_s),
    .io_co(FullAdder_32_io_co)
  );
  FullAdder FullAdder_33 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_33_io_a),
    .io_b(FullAdder_33_io_b),
    .io_ci(FullAdder_33_io_ci),
    .io_s(FullAdder_33_io_s),
    .io_co(FullAdder_33_io_co)
  );
  FullAdder FullAdder_34 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_34_io_a),
    .io_b(FullAdder_34_io_b),
    .io_ci(FullAdder_34_io_ci),
    .io_s(FullAdder_34_io_s),
    .io_co(FullAdder_34_io_co)
  );
  FullAdder FullAdder_35 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_35_io_a),
    .io_b(FullAdder_35_io_b),
    .io_ci(FullAdder_35_io_ci),
    .io_s(FullAdder_35_io_s),
    .io_co(FullAdder_35_io_co)
  );
  FullAdder FullAdder_36 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_36_io_a),
    .io_b(FullAdder_36_io_b),
    .io_ci(FullAdder_36_io_ci),
    .io_s(FullAdder_36_io_s),
    .io_co(FullAdder_36_io_co)
  );
  FullAdder FullAdder_37 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_37_io_a),
    .io_b(FullAdder_37_io_b),
    .io_ci(FullAdder_37_io_ci),
    .io_s(FullAdder_37_io_s),
    .io_co(FullAdder_37_io_co)
  );
  FullAdder FullAdder_38 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_38_io_a),
    .io_b(FullAdder_38_io_b),
    .io_ci(FullAdder_38_io_ci),
    .io_s(FullAdder_38_io_s),
    .io_co(FullAdder_38_io_co)
  );
  FullAdder FullAdder_39 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_39_io_a),
    .io_b(FullAdder_39_io_b),
    .io_ci(FullAdder_39_io_ci),
    .io_s(FullAdder_39_io_s),
    .io_co(FullAdder_39_io_co)
  );
  FullAdder FullAdder_40 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_40_io_a),
    .io_b(FullAdder_40_io_b),
    .io_ci(FullAdder_40_io_ci),
    .io_s(FullAdder_40_io_s),
    .io_co(FullAdder_40_io_co)
  );
  FullAdder FullAdder_41 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_41_io_a),
    .io_b(FullAdder_41_io_b),
    .io_ci(FullAdder_41_io_ci),
    .io_s(FullAdder_41_io_s),
    .io_co(FullAdder_41_io_co)
  );
  FullAdder FullAdder_42 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_42_io_a),
    .io_b(FullAdder_42_io_b),
    .io_ci(FullAdder_42_io_ci),
    .io_s(FullAdder_42_io_s),
    .io_co(FullAdder_42_io_co)
  );
  FullAdder FullAdder_43 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_43_io_a),
    .io_b(FullAdder_43_io_b),
    .io_ci(FullAdder_43_io_ci),
    .io_s(FullAdder_43_io_s),
    .io_co(FullAdder_43_io_co)
  );
  FullAdder FullAdder_44 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_44_io_a),
    .io_b(FullAdder_44_io_b),
    .io_ci(FullAdder_44_io_ci),
    .io_s(FullAdder_44_io_s),
    .io_co(FullAdder_44_io_co)
  );
  HalfAdder HalfAdder_4 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_4_io_a),
    .io_b(HalfAdder_4_io_b),
    .io_s(HalfAdder_4_io_s),
    .io_co(HalfAdder_4_io_co)
  );
  FullAdder FullAdder_45 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_45_io_a),
    .io_b(FullAdder_45_io_b),
    .io_ci(FullAdder_45_io_ci),
    .io_s(FullAdder_45_io_s),
    .io_co(FullAdder_45_io_co)
  );
  FullAdder FullAdder_46 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_46_io_a),
    .io_b(FullAdder_46_io_b),
    .io_ci(FullAdder_46_io_ci),
    .io_s(FullAdder_46_io_s),
    .io_co(FullAdder_46_io_co)
  );
  FullAdder FullAdder_47 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_47_io_a),
    .io_b(FullAdder_47_io_b),
    .io_ci(FullAdder_47_io_ci),
    .io_s(FullAdder_47_io_s),
    .io_co(FullAdder_47_io_co)
  );
  FullAdder FullAdder_48 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_48_io_a),
    .io_b(FullAdder_48_io_b),
    .io_ci(FullAdder_48_io_ci),
    .io_s(FullAdder_48_io_s),
    .io_co(FullAdder_48_io_co)
  );
  FullAdder FullAdder_49 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_49_io_a),
    .io_b(FullAdder_49_io_b),
    .io_ci(FullAdder_49_io_ci),
    .io_s(FullAdder_49_io_s),
    .io_co(FullAdder_49_io_co)
  );
  FullAdder FullAdder_50 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_50_io_a),
    .io_b(FullAdder_50_io_b),
    .io_ci(FullAdder_50_io_ci),
    .io_s(FullAdder_50_io_s),
    .io_co(FullAdder_50_io_co)
  );
  FullAdder FullAdder_51 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_51_io_a),
    .io_b(FullAdder_51_io_b),
    .io_ci(FullAdder_51_io_ci),
    .io_s(FullAdder_51_io_s),
    .io_co(FullAdder_51_io_co)
  );
  FullAdder FullAdder_52 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_52_io_a),
    .io_b(FullAdder_52_io_b),
    .io_ci(FullAdder_52_io_ci),
    .io_s(FullAdder_52_io_s),
    .io_co(FullAdder_52_io_co)
  );
  FullAdder FullAdder_53 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_53_io_a),
    .io_b(FullAdder_53_io_b),
    .io_ci(FullAdder_53_io_ci),
    .io_s(FullAdder_53_io_s),
    .io_co(FullAdder_53_io_co)
  );
  FullAdder FullAdder_54 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_54_io_a),
    .io_b(FullAdder_54_io_b),
    .io_ci(FullAdder_54_io_ci),
    .io_s(FullAdder_54_io_s),
    .io_co(FullAdder_54_io_co)
  );
  FullAdder FullAdder_55 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_55_io_a),
    .io_b(FullAdder_55_io_b),
    .io_ci(FullAdder_55_io_ci),
    .io_s(FullAdder_55_io_s),
    .io_co(FullAdder_55_io_co)
  );
  FullAdder FullAdder_56 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_56_io_a),
    .io_b(FullAdder_56_io_b),
    .io_ci(FullAdder_56_io_ci),
    .io_s(FullAdder_56_io_s),
    .io_co(FullAdder_56_io_co)
  );
  FullAdder FullAdder_57 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_57_io_a),
    .io_b(FullAdder_57_io_b),
    .io_ci(FullAdder_57_io_ci),
    .io_s(FullAdder_57_io_s),
    .io_co(FullAdder_57_io_co)
  );
  FullAdder FullAdder_58 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_58_io_a),
    .io_b(FullAdder_58_io_b),
    .io_ci(FullAdder_58_io_ci),
    .io_s(FullAdder_58_io_s),
    .io_co(FullAdder_58_io_co)
  );
  FullAdder FullAdder_59 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_59_io_a),
    .io_b(FullAdder_59_io_b),
    .io_ci(FullAdder_59_io_ci),
    .io_s(FullAdder_59_io_s),
    .io_co(FullAdder_59_io_co)
  );
  FullAdder FullAdder_60 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_60_io_a),
    .io_b(FullAdder_60_io_b),
    .io_ci(FullAdder_60_io_ci),
    .io_s(FullAdder_60_io_s),
    .io_co(FullAdder_60_io_co)
  );
  FullAdder FullAdder_61 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_61_io_a),
    .io_b(FullAdder_61_io_b),
    .io_ci(FullAdder_61_io_ci),
    .io_s(FullAdder_61_io_s),
    .io_co(FullAdder_61_io_co)
  );
  FullAdder FullAdder_62 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_62_io_a),
    .io_b(FullAdder_62_io_b),
    .io_ci(FullAdder_62_io_ci),
    .io_s(FullAdder_62_io_s),
    .io_co(FullAdder_62_io_co)
  );
  HalfAdder HalfAdder_5 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_5_io_a),
    .io_b(HalfAdder_5_io_b),
    .io_s(HalfAdder_5_io_s),
    .io_co(HalfAdder_5_io_co)
  );
  FullAdder FullAdder_63 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_63_io_a),
    .io_b(FullAdder_63_io_b),
    .io_ci(FullAdder_63_io_ci),
    .io_s(FullAdder_63_io_s),
    .io_co(FullAdder_63_io_co)
  );
  FullAdder FullAdder_64 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_64_io_a),
    .io_b(FullAdder_64_io_b),
    .io_ci(FullAdder_64_io_ci),
    .io_s(FullAdder_64_io_s),
    .io_co(FullAdder_64_io_co)
  );
  FullAdder FullAdder_65 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_65_io_a),
    .io_b(FullAdder_65_io_b),
    .io_ci(FullAdder_65_io_ci),
    .io_s(FullAdder_65_io_s),
    .io_co(FullAdder_65_io_co)
  );
  FullAdder FullAdder_66 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_66_io_a),
    .io_b(FullAdder_66_io_b),
    .io_ci(FullAdder_66_io_ci),
    .io_s(FullAdder_66_io_s),
    .io_co(FullAdder_66_io_co)
  );
  FullAdder FullAdder_67 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_67_io_a),
    .io_b(FullAdder_67_io_b),
    .io_ci(FullAdder_67_io_ci),
    .io_s(FullAdder_67_io_s),
    .io_co(FullAdder_67_io_co)
  );
  FullAdder FullAdder_68 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_68_io_a),
    .io_b(FullAdder_68_io_b),
    .io_ci(FullAdder_68_io_ci),
    .io_s(FullAdder_68_io_s),
    .io_co(FullAdder_68_io_co)
  );
  FullAdder FullAdder_69 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_69_io_a),
    .io_b(FullAdder_69_io_b),
    .io_ci(FullAdder_69_io_ci),
    .io_s(FullAdder_69_io_s),
    .io_co(FullAdder_69_io_co)
  );
  FullAdder FullAdder_70 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_70_io_a),
    .io_b(FullAdder_70_io_b),
    .io_ci(FullAdder_70_io_ci),
    .io_s(FullAdder_70_io_s),
    .io_co(FullAdder_70_io_co)
  );
  FullAdder FullAdder_71 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_71_io_a),
    .io_b(FullAdder_71_io_b),
    .io_ci(FullAdder_71_io_ci),
    .io_s(FullAdder_71_io_s),
    .io_co(FullAdder_71_io_co)
  );
  FullAdder FullAdder_72 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_72_io_a),
    .io_b(FullAdder_72_io_b),
    .io_ci(FullAdder_72_io_ci),
    .io_s(FullAdder_72_io_s),
    .io_co(FullAdder_72_io_co)
  );
  FullAdder FullAdder_73 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_73_io_a),
    .io_b(FullAdder_73_io_b),
    .io_ci(FullAdder_73_io_ci),
    .io_s(FullAdder_73_io_s),
    .io_co(FullAdder_73_io_co)
  );
  FullAdder FullAdder_74 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_74_io_a),
    .io_b(FullAdder_74_io_b),
    .io_ci(FullAdder_74_io_ci),
    .io_s(FullAdder_74_io_s),
    .io_co(FullAdder_74_io_co)
  );
  FullAdder FullAdder_75 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_75_io_a),
    .io_b(FullAdder_75_io_b),
    .io_ci(FullAdder_75_io_ci),
    .io_s(FullAdder_75_io_s),
    .io_co(FullAdder_75_io_co)
  );
  FullAdder FullAdder_76 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_76_io_a),
    .io_b(FullAdder_76_io_b),
    .io_ci(FullAdder_76_io_ci),
    .io_s(FullAdder_76_io_s),
    .io_co(FullAdder_76_io_co)
  );
  FullAdder FullAdder_77 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_77_io_a),
    .io_b(FullAdder_77_io_b),
    .io_ci(FullAdder_77_io_ci),
    .io_s(FullAdder_77_io_s),
    .io_co(FullAdder_77_io_co)
  );
  FullAdder FullAdder_78 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_78_io_a),
    .io_b(FullAdder_78_io_b),
    .io_ci(FullAdder_78_io_ci),
    .io_s(FullAdder_78_io_s),
    .io_co(FullAdder_78_io_co)
  );
  FullAdder FullAdder_79 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_79_io_a),
    .io_b(FullAdder_79_io_b),
    .io_ci(FullAdder_79_io_ci),
    .io_s(FullAdder_79_io_s),
    .io_co(FullAdder_79_io_co)
  );
  FullAdder FullAdder_80 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_80_io_a),
    .io_b(FullAdder_80_io_b),
    .io_ci(FullAdder_80_io_ci),
    .io_s(FullAdder_80_io_s),
    .io_co(FullAdder_80_io_co)
  );
  FullAdder FullAdder_81 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_81_io_a),
    .io_b(FullAdder_81_io_b),
    .io_ci(FullAdder_81_io_ci),
    .io_s(FullAdder_81_io_s),
    .io_co(FullAdder_81_io_co)
  );
  FullAdder FullAdder_82 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_82_io_a),
    .io_b(FullAdder_82_io_b),
    .io_ci(FullAdder_82_io_ci),
    .io_s(FullAdder_82_io_s),
    .io_co(FullAdder_82_io_co)
  );
  FullAdder FullAdder_83 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_83_io_a),
    .io_b(FullAdder_83_io_b),
    .io_ci(FullAdder_83_io_ci),
    .io_s(FullAdder_83_io_s),
    .io_co(FullAdder_83_io_co)
  );
  HalfAdder HalfAdder_6 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_6_io_a),
    .io_b(HalfAdder_6_io_b),
    .io_s(HalfAdder_6_io_s),
    .io_co(HalfAdder_6_io_co)
  );
  FullAdder FullAdder_84 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_84_io_a),
    .io_b(FullAdder_84_io_b),
    .io_ci(FullAdder_84_io_ci),
    .io_s(FullAdder_84_io_s),
    .io_co(FullAdder_84_io_co)
  );
  FullAdder FullAdder_85 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_85_io_a),
    .io_b(FullAdder_85_io_b),
    .io_ci(FullAdder_85_io_ci),
    .io_s(FullAdder_85_io_s),
    .io_co(FullAdder_85_io_co)
  );
  FullAdder FullAdder_86 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_86_io_a),
    .io_b(FullAdder_86_io_b),
    .io_ci(FullAdder_86_io_ci),
    .io_s(FullAdder_86_io_s),
    .io_co(FullAdder_86_io_co)
  );
  FullAdder FullAdder_87 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_87_io_a),
    .io_b(FullAdder_87_io_b),
    .io_ci(FullAdder_87_io_ci),
    .io_s(FullAdder_87_io_s),
    .io_co(FullAdder_87_io_co)
  );
  FullAdder FullAdder_88 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_88_io_a),
    .io_b(FullAdder_88_io_b),
    .io_ci(FullAdder_88_io_ci),
    .io_s(FullAdder_88_io_s),
    .io_co(FullAdder_88_io_co)
  );
  FullAdder FullAdder_89 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_89_io_a),
    .io_b(FullAdder_89_io_b),
    .io_ci(FullAdder_89_io_ci),
    .io_s(FullAdder_89_io_s),
    .io_co(FullAdder_89_io_co)
  );
  FullAdder FullAdder_90 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_90_io_a),
    .io_b(FullAdder_90_io_b),
    .io_ci(FullAdder_90_io_ci),
    .io_s(FullAdder_90_io_s),
    .io_co(FullAdder_90_io_co)
  );
  FullAdder FullAdder_91 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_91_io_a),
    .io_b(FullAdder_91_io_b),
    .io_ci(FullAdder_91_io_ci),
    .io_s(FullAdder_91_io_s),
    .io_co(FullAdder_91_io_co)
  );
  FullAdder FullAdder_92 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_92_io_a),
    .io_b(FullAdder_92_io_b),
    .io_ci(FullAdder_92_io_ci),
    .io_s(FullAdder_92_io_s),
    .io_co(FullAdder_92_io_co)
  );
  FullAdder FullAdder_93 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_93_io_a),
    .io_b(FullAdder_93_io_b),
    .io_ci(FullAdder_93_io_ci),
    .io_s(FullAdder_93_io_s),
    .io_co(FullAdder_93_io_co)
  );
  FullAdder FullAdder_94 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_94_io_a),
    .io_b(FullAdder_94_io_b),
    .io_ci(FullAdder_94_io_ci),
    .io_s(FullAdder_94_io_s),
    .io_co(FullAdder_94_io_co)
  );
  FullAdder FullAdder_95 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_95_io_a),
    .io_b(FullAdder_95_io_b),
    .io_ci(FullAdder_95_io_ci),
    .io_s(FullAdder_95_io_s),
    .io_co(FullAdder_95_io_co)
  );
  FullAdder FullAdder_96 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_96_io_a),
    .io_b(FullAdder_96_io_b),
    .io_ci(FullAdder_96_io_ci),
    .io_s(FullAdder_96_io_s),
    .io_co(FullAdder_96_io_co)
  );
  FullAdder FullAdder_97 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_97_io_a),
    .io_b(FullAdder_97_io_b),
    .io_ci(FullAdder_97_io_ci),
    .io_s(FullAdder_97_io_s),
    .io_co(FullAdder_97_io_co)
  );
  FullAdder FullAdder_98 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_98_io_a),
    .io_b(FullAdder_98_io_b),
    .io_ci(FullAdder_98_io_ci),
    .io_s(FullAdder_98_io_s),
    .io_co(FullAdder_98_io_co)
  );
  FullAdder FullAdder_99 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_99_io_a),
    .io_b(FullAdder_99_io_b),
    .io_ci(FullAdder_99_io_ci),
    .io_s(FullAdder_99_io_s),
    .io_co(FullAdder_99_io_co)
  );
  FullAdder FullAdder_100 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_100_io_a),
    .io_b(FullAdder_100_io_b),
    .io_ci(FullAdder_100_io_ci),
    .io_s(FullAdder_100_io_s),
    .io_co(FullAdder_100_io_co)
  );
  FullAdder FullAdder_101 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_101_io_a),
    .io_b(FullAdder_101_io_b),
    .io_ci(FullAdder_101_io_ci),
    .io_s(FullAdder_101_io_s),
    .io_co(FullAdder_101_io_co)
  );
  FullAdder FullAdder_102 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_102_io_a),
    .io_b(FullAdder_102_io_b),
    .io_ci(FullAdder_102_io_ci),
    .io_s(FullAdder_102_io_s),
    .io_co(FullAdder_102_io_co)
  );
  FullAdder FullAdder_103 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_103_io_a),
    .io_b(FullAdder_103_io_b),
    .io_ci(FullAdder_103_io_ci),
    .io_s(FullAdder_103_io_s),
    .io_co(FullAdder_103_io_co)
  );
  FullAdder FullAdder_104 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_104_io_a),
    .io_b(FullAdder_104_io_b),
    .io_ci(FullAdder_104_io_ci),
    .io_s(FullAdder_104_io_s),
    .io_co(FullAdder_104_io_co)
  );
  FullAdder FullAdder_105 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_105_io_a),
    .io_b(FullAdder_105_io_b),
    .io_ci(FullAdder_105_io_ci),
    .io_s(FullAdder_105_io_s),
    .io_co(FullAdder_105_io_co)
  );
  FullAdder FullAdder_106 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_106_io_a),
    .io_b(FullAdder_106_io_b),
    .io_ci(FullAdder_106_io_ci),
    .io_s(FullAdder_106_io_s),
    .io_co(FullAdder_106_io_co)
  );
  FullAdder FullAdder_107 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_107_io_a),
    .io_b(FullAdder_107_io_b),
    .io_ci(FullAdder_107_io_ci),
    .io_s(FullAdder_107_io_s),
    .io_co(FullAdder_107_io_co)
  );
  FullAdder FullAdder_108 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_108_io_a),
    .io_b(FullAdder_108_io_b),
    .io_ci(FullAdder_108_io_ci),
    .io_s(FullAdder_108_io_s),
    .io_co(FullAdder_108_io_co)
  );
  FullAdder FullAdder_109 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_109_io_a),
    .io_b(FullAdder_109_io_b),
    .io_ci(FullAdder_109_io_ci),
    .io_s(FullAdder_109_io_s),
    .io_co(FullAdder_109_io_co)
  );
  FullAdder FullAdder_110 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_110_io_a),
    .io_b(FullAdder_110_io_b),
    .io_ci(FullAdder_110_io_ci),
    .io_s(FullAdder_110_io_s),
    .io_co(FullAdder_110_io_co)
  );
  FullAdder FullAdder_111 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_111_io_a),
    .io_b(FullAdder_111_io_b),
    .io_ci(FullAdder_111_io_ci),
    .io_s(FullAdder_111_io_s),
    .io_co(FullAdder_111_io_co)
  );
  FullAdder FullAdder_112 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_112_io_a),
    .io_b(FullAdder_112_io_b),
    .io_ci(FullAdder_112_io_ci),
    .io_s(FullAdder_112_io_s),
    .io_co(FullAdder_112_io_co)
  );
  FullAdder FullAdder_113 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_113_io_a),
    .io_b(FullAdder_113_io_b),
    .io_ci(FullAdder_113_io_ci),
    .io_s(FullAdder_113_io_s),
    .io_co(FullAdder_113_io_co)
  );
  FullAdder FullAdder_114 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_114_io_a),
    .io_b(FullAdder_114_io_b),
    .io_ci(FullAdder_114_io_ci),
    .io_s(FullAdder_114_io_s),
    .io_co(FullAdder_114_io_co)
  );
  FullAdder FullAdder_115 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_115_io_a),
    .io_b(FullAdder_115_io_b),
    .io_ci(FullAdder_115_io_ci),
    .io_s(FullAdder_115_io_s),
    .io_co(FullAdder_115_io_co)
  );
  FullAdder FullAdder_116 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_116_io_a),
    .io_b(FullAdder_116_io_b),
    .io_ci(FullAdder_116_io_ci),
    .io_s(FullAdder_116_io_s),
    .io_co(FullAdder_116_io_co)
  );
  FullAdder FullAdder_117 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_117_io_a),
    .io_b(FullAdder_117_io_b),
    .io_ci(FullAdder_117_io_ci),
    .io_s(FullAdder_117_io_s),
    .io_co(FullAdder_117_io_co)
  );
  FullAdder FullAdder_118 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_118_io_a),
    .io_b(FullAdder_118_io_b),
    .io_ci(FullAdder_118_io_ci),
    .io_s(FullAdder_118_io_s),
    .io_co(FullAdder_118_io_co)
  );
  FullAdder FullAdder_119 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_119_io_a),
    .io_b(FullAdder_119_io_b),
    .io_ci(FullAdder_119_io_ci),
    .io_s(FullAdder_119_io_s),
    .io_co(FullAdder_119_io_co)
  );
  FullAdder FullAdder_120 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_120_io_a),
    .io_b(FullAdder_120_io_b),
    .io_ci(FullAdder_120_io_ci),
    .io_s(FullAdder_120_io_s),
    .io_co(FullAdder_120_io_co)
  );
  FullAdder FullAdder_121 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_121_io_a),
    .io_b(FullAdder_121_io_b),
    .io_ci(FullAdder_121_io_ci),
    .io_s(FullAdder_121_io_s),
    .io_co(FullAdder_121_io_co)
  );
  FullAdder FullAdder_122 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_122_io_a),
    .io_b(FullAdder_122_io_b),
    .io_ci(FullAdder_122_io_ci),
    .io_s(FullAdder_122_io_s),
    .io_co(FullAdder_122_io_co)
  );
  FullAdder FullAdder_123 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_123_io_a),
    .io_b(FullAdder_123_io_b),
    .io_ci(FullAdder_123_io_ci),
    .io_s(FullAdder_123_io_s),
    .io_co(FullAdder_123_io_co)
  );
  FullAdder FullAdder_124 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_124_io_a),
    .io_b(FullAdder_124_io_b),
    .io_ci(FullAdder_124_io_ci),
    .io_s(FullAdder_124_io_s),
    .io_co(FullAdder_124_io_co)
  );
  FullAdder FullAdder_125 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_125_io_a),
    .io_b(FullAdder_125_io_b),
    .io_ci(FullAdder_125_io_ci),
    .io_s(FullAdder_125_io_s),
    .io_co(FullAdder_125_io_co)
  );
  FullAdder FullAdder_126 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_126_io_a),
    .io_b(FullAdder_126_io_b),
    .io_ci(FullAdder_126_io_ci),
    .io_s(FullAdder_126_io_s),
    .io_co(FullAdder_126_io_co)
  );
  FullAdder FullAdder_127 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_127_io_a),
    .io_b(FullAdder_127_io_b),
    .io_ci(FullAdder_127_io_ci),
    .io_s(FullAdder_127_io_s),
    .io_co(FullAdder_127_io_co)
  );
  FullAdder FullAdder_128 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_128_io_a),
    .io_b(FullAdder_128_io_b),
    .io_ci(FullAdder_128_io_ci),
    .io_s(FullAdder_128_io_s),
    .io_co(FullAdder_128_io_co)
  );
  FullAdder FullAdder_129 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_129_io_a),
    .io_b(FullAdder_129_io_b),
    .io_ci(FullAdder_129_io_ci),
    .io_s(FullAdder_129_io_s),
    .io_co(FullAdder_129_io_co)
  );
  FullAdder FullAdder_130 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_130_io_a),
    .io_b(FullAdder_130_io_b),
    .io_ci(FullAdder_130_io_ci),
    .io_s(FullAdder_130_io_s),
    .io_co(FullAdder_130_io_co)
  );
  FullAdder FullAdder_131 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_131_io_a),
    .io_b(FullAdder_131_io_b),
    .io_ci(FullAdder_131_io_ci),
    .io_s(FullAdder_131_io_s),
    .io_co(FullAdder_131_io_co)
  );
  FullAdder FullAdder_132 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_132_io_a),
    .io_b(FullAdder_132_io_b),
    .io_ci(FullAdder_132_io_ci),
    .io_s(FullAdder_132_io_s),
    .io_co(FullAdder_132_io_co)
  );
  FullAdder FullAdder_133 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_133_io_a),
    .io_b(FullAdder_133_io_b),
    .io_ci(FullAdder_133_io_ci),
    .io_s(FullAdder_133_io_s),
    .io_co(FullAdder_133_io_co)
  );
  FullAdder FullAdder_134 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_134_io_a),
    .io_b(FullAdder_134_io_b),
    .io_ci(FullAdder_134_io_ci),
    .io_s(FullAdder_134_io_s),
    .io_co(FullAdder_134_io_co)
  );
  FullAdder FullAdder_135 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_135_io_a),
    .io_b(FullAdder_135_io_b),
    .io_ci(FullAdder_135_io_ci),
    .io_s(FullAdder_135_io_s),
    .io_co(FullAdder_135_io_co)
  );
  FullAdder FullAdder_136 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_136_io_a),
    .io_b(FullAdder_136_io_b),
    .io_ci(FullAdder_136_io_ci),
    .io_s(FullAdder_136_io_s),
    .io_co(FullAdder_136_io_co)
  );
  FullAdder FullAdder_137 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_137_io_a),
    .io_b(FullAdder_137_io_b),
    .io_ci(FullAdder_137_io_ci),
    .io_s(FullAdder_137_io_s),
    .io_co(FullAdder_137_io_co)
  );
  FullAdder FullAdder_138 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_138_io_a),
    .io_b(FullAdder_138_io_b),
    .io_ci(FullAdder_138_io_ci),
    .io_s(FullAdder_138_io_s),
    .io_co(FullAdder_138_io_co)
  );
  FullAdder FullAdder_139 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_139_io_a),
    .io_b(FullAdder_139_io_b),
    .io_ci(FullAdder_139_io_ci),
    .io_s(FullAdder_139_io_s),
    .io_co(FullAdder_139_io_co)
  );
  FullAdder FullAdder_140 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_140_io_a),
    .io_b(FullAdder_140_io_b),
    .io_ci(FullAdder_140_io_ci),
    .io_s(FullAdder_140_io_s),
    .io_co(FullAdder_140_io_co)
  );
  FullAdder FullAdder_141 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_141_io_a),
    .io_b(FullAdder_141_io_b),
    .io_ci(FullAdder_141_io_ci),
    .io_s(FullAdder_141_io_s),
    .io_co(FullAdder_141_io_co)
  );
  FullAdder FullAdder_142 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_142_io_a),
    .io_b(FullAdder_142_io_b),
    .io_ci(FullAdder_142_io_ci),
    .io_s(FullAdder_142_io_s),
    .io_co(FullAdder_142_io_co)
  );
  FullAdder FullAdder_143 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_143_io_a),
    .io_b(FullAdder_143_io_b),
    .io_ci(FullAdder_143_io_ci),
    .io_s(FullAdder_143_io_s),
    .io_co(FullAdder_143_io_co)
  );
  FullAdder FullAdder_144 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_144_io_a),
    .io_b(FullAdder_144_io_b),
    .io_ci(FullAdder_144_io_ci),
    .io_s(FullAdder_144_io_s),
    .io_co(FullAdder_144_io_co)
  );
  FullAdder FullAdder_145 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_145_io_a),
    .io_b(FullAdder_145_io_b),
    .io_ci(FullAdder_145_io_ci),
    .io_s(FullAdder_145_io_s),
    .io_co(FullAdder_145_io_co)
  );
  FullAdder FullAdder_146 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_146_io_a),
    .io_b(FullAdder_146_io_b),
    .io_ci(FullAdder_146_io_ci),
    .io_s(FullAdder_146_io_s),
    .io_co(FullAdder_146_io_co)
  );
  FullAdder FullAdder_147 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_147_io_a),
    .io_b(FullAdder_147_io_b),
    .io_ci(FullAdder_147_io_ci),
    .io_s(FullAdder_147_io_s),
    .io_co(FullAdder_147_io_co)
  );
  FullAdder FullAdder_148 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_148_io_a),
    .io_b(FullAdder_148_io_b),
    .io_ci(FullAdder_148_io_ci),
    .io_s(FullAdder_148_io_s),
    .io_co(FullAdder_148_io_co)
  );
  FullAdder FullAdder_149 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_149_io_a),
    .io_b(FullAdder_149_io_b),
    .io_ci(FullAdder_149_io_ci),
    .io_s(FullAdder_149_io_s),
    .io_co(FullAdder_149_io_co)
  );
  FullAdder FullAdder_150 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_150_io_a),
    .io_b(FullAdder_150_io_b),
    .io_ci(FullAdder_150_io_ci),
    .io_s(FullAdder_150_io_s),
    .io_co(FullAdder_150_io_co)
  );
  FullAdder FullAdder_151 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_151_io_a),
    .io_b(FullAdder_151_io_b),
    .io_ci(FullAdder_151_io_ci),
    .io_s(FullAdder_151_io_s),
    .io_co(FullAdder_151_io_co)
  );
  FullAdder FullAdder_152 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_152_io_a),
    .io_b(FullAdder_152_io_b),
    .io_ci(FullAdder_152_io_ci),
    .io_s(FullAdder_152_io_s),
    .io_co(FullAdder_152_io_co)
  );
  FullAdder FullAdder_153 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_153_io_a),
    .io_b(FullAdder_153_io_b),
    .io_ci(FullAdder_153_io_ci),
    .io_s(FullAdder_153_io_s),
    .io_co(FullAdder_153_io_co)
  );
  FullAdder FullAdder_154 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_154_io_a),
    .io_b(FullAdder_154_io_b),
    .io_ci(FullAdder_154_io_ci),
    .io_s(FullAdder_154_io_s),
    .io_co(FullAdder_154_io_co)
  );
  FullAdder FullAdder_155 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_155_io_a),
    .io_b(FullAdder_155_io_b),
    .io_ci(FullAdder_155_io_ci),
    .io_s(FullAdder_155_io_s),
    .io_co(FullAdder_155_io_co)
  );
  FullAdder FullAdder_156 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_156_io_a),
    .io_b(FullAdder_156_io_b),
    .io_ci(FullAdder_156_io_ci),
    .io_s(FullAdder_156_io_s),
    .io_co(FullAdder_156_io_co)
  );
  FullAdder FullAdder_157 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_157_io_a),
    .io_b(FullAdder_157_io_b),
    .io_ci(FullAdder_157_io_ci),
    .io_s(FullAdder_157_io_s),
    .io_co(FullAdder_157_io_co)
  );
  FullAdder FullAdder_158 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_158_io_a),
    .io_b(FullAdder_158_io_b),
    .io_ci(FullAdder_158_io_ci),
    .io_s(FullAdder_158_io_s),
    .io_co(FullAdder_158_io_co)
  );
  FullAdder FullAdder_159 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_159_io_a),
    .io_b(FullAdder_159_io_b),
    .io_ci(FullAdder_159_io_ci),
    .io_s(FullAdder_159_io_s),
    .io_co(FullAdder_159_io_co)
  );
  FullAdder FullAdder_160 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_160_io_a),
    .io_b(FullAdder_160_io_b),
    .io_ci(FullAdder_160_io_ci),
    .io_s(FullAdder_160_io_s),
    .io_co(FullAdder_160_io_co)
  );
  FullAdder FullAdder_161 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_161_io_a),
    .io_b(FullAdder_161_io_b),
    .io_ci(FullAdder_161_io_ci),
    .io_s(FullAdder_161_io_s),
    .io_co(FullAdder_161_io_co)
  );
  FullAdder FullAdder_162 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_162_io_a),
    .io_b(FullAdder_162_io_b),
    .io_ci(FullAdder_162_io_ci),
    .io_s(FullAdder_162_io_s),
    .io_co(FullAdder_162_io_co)
  );
  FullAdder FullAdder_163 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_163_io_a),
    .io_b(FullAdder_163_io_b),
    .io_ci(FullAdder_163_io_ci),
    .io_s(FullAdder_163_io_s),
    .io_co(FullAdder_163_io_co)
  );
  FullAdder FullAdder_164 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_164_io_a),
    .io_b(FullAdder_164_io_b),
    .io_ci(FullAdder_164_io_ci),
    .io_s(FullAdder_164_io_s),
    .io_co(FullAdder_164_io_co)
  );
  HalfAdder HalfAdder_7 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_7_io_a),
    .io_b(HalfAdder_7_io_b),
    .io_s(HalfAdder_7_io_s),
    .io_co(HalfAdder_7_io_co)
  );
  FullAdder FullAdder_165 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_165_io_a),
    .io_b(FullAdder_165_io_b),
    .io_ci(FullAdder_165_io_ci),
    .io_s(FullAdder_165_io_s),
    .io_co(FullAdder_165_io_co)
  );
  FullAdder FullAdder_166 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_166_io_a),
    .io_b(FullAdder_166_io_b),
    .io_ci(FullAdder_166_io_ci),
    .io_s(FullAdder_166_io_s),
    .io_co(FullAdder_166_io_co)
  );
  FullAdder FullAdder_167 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_167_io_a),
    .io_b(FullAdder_167_io_b),
    .io_ci(FullAdder_167_io_ci),
    .io_s(FullAdder_167_io_s),
    .io_co(FullAdder_167_io_co)
  );
  FullAdder FullAdder_168 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_168_io_a),
    .io_b(FullAdder_168_io_b),
    .io_ci(FullAdder_168_io_ci),
    .io_s(FullAdder_168_io_s),
    .io_co(FullAdder_168_io_co)
  );
  FullAdder FullAdder_169 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_169_io_a),
    .io_b(FullAdder_169_io_b),
    .io_ci(FullAdder_169_io_ci),
    .io_s(FullAdder_169_io_s),
    .io_co(FullAdder_169_io_co)
  );
  FullAdder FullAdder_170 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_170_io_a),
    .io_b(FullAdder_170_io_b),
    .io_ci(FullAdder_170_io_ci),
    .io_s(FullAdder_170_io_s),
    .io_co(FullAdder_170_io_co)
  );
  FullAdder FullAdder_171 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_171_io_a),
    .io_b(FullAdder_171_io_b),
    .io_ci(FullAdder_171_io_ci),
    .io_s(FullAdder_171_io_s),
    .io_co(FullAdder_171_io_co)
  );
  FullAdder FullAdder_172 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_172_io_a),
    .io_b(FullAdder_172_io_b),
    .io_ci(FullAdder_172_io_ci),
    .io_s(FullAdder_172_io_s),
    .io_co(FullAdder_172_io_co)
  );
  FullAdder FullAdder_173 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_173_io_a),
    .io_b(FullAdder_173_io_b),
    .io_ci(FullAdder_173_io_ci),
    .io_s(FullAdder_173_io_s),
    .io_co(FullAdder_173_io_co)
  );
  FullAdder FullAdder_174 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_174_io_a),
    .io_b(FullAdder_174_io_b),
    .io_ci(FullAdder_174_io_ci),
    .io_s(FullAdder_174_io_s),
    .io_co(FullAdder_174_io_co)
  );
  FullAdder FullAdder_175 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_175_io_a),
    .io_b(FullAdder_175_io_b),
    .io_ci(FullAdder_175_io_ci),
    .io_s(FullAdder_175_io_s),
    .io_co(FullAdder_175_io_co)
  );
  FullAdder FullAdder_176 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_176_io_a),
    .io_b(FullAdder_176_io_b),
    .io_ci(FullAdder_176_io_ci),
    .io_s(FullAdder_176_io_s),
    .io_co(FullAdder_176_io_co)
  );
  FullAdder FullAdder_177 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_177_io_a),
    .io_b(FullAdder_177_io_b),
    .io_ci(FullAdder_177_io_ci),
    .io_s(FullAdder_177_io_s),
    .io_co(FullAdder_177_io_co)
  );
  FullAdder FullAdder_178 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_178_io_a),
    .io_b(FullAdder_178_io_b),
    .io_ci(FullAdder_178_io_ci),
    .io_s(FullAdder_178_io_s),
    .io_co(FullAdder_178_io_co)
  );
  FullAdder FullAdder_179 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_179_io_a),
    .io_b(FullAdder_179_io_b),
    .io_ci(FullAdder_179_io_ci),
    .io_s(FullAdder_179_io_s),
    .io_co(FullAdder_179_io_co)
  );
  FullAdder FullAdder_180 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_180_io_a),
    .io_b(FullAdder_180_io_b),
    .io_ci(FullAdder_180_io_ci),
    .io_s(FullAdder_180_io_s),
    .io_co(FullAdder_180_io_co)
  );
  FullAdder FullAdder_181 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_181_io_a),
    .io_b(FullAdder_181_io_b),
    .io_ci(FullAdder_181_io_ci),
    .io_s(FullAdder_181_io_s),
    .io_co(FullAdder_181_io_co)
  );
  FullAdder FullAdder_182 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_182_io_a),
    .io_b(FullAdder_182_io_b),
    .io_ci(FullAdder_182_io_ci),
    .io_s(FullAdder_182_io_s),
    .io_co(FullAdder_182_io_co)
  );
  FullAdder FullAdder_183 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_183_io_a),
    .io_b(FullAdder_183_io_b),
    .io_ci(FullAdder_183_io_ci),
    .io_s(FullAdder_183_io_s),
    .io_co(FullAdder_183_io_co)
  );
  FullAdder FullAdder_184 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_184_io_a),
    .io_b(FullAdder_184_io_b),
    .io_ci(FullAdder_184_io_ci),
    .io_s(FullAdder_184_io_s),
    .io_co(FullAdder_184_io_co)
  );
  FullAdder FullAdder_185 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_185_io_a),
    .io_b(FullAdder_185_io_b),
    .io_ci(FullAdder_185_io_ci),
    .io_s(FullAdder_185_io_s),
    .io_co(FullAdder_185_io_co)
  );
  FullAdder FullAdder_186 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_186_io_a),
    .io_b(FullAdder_186_io_b),
    .io_ci(FullAdder_186_io_ci),
    .io_s(FullAdder_186_io_s),
    .io_co(FullAdder_186_io_co)
  );
  FullAdder FullAdder_187 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_187_io_a),
    .io_b(FullAdder_187_io_b),
    .io_ci(FullAdder_187_io_ci),
    .io_s(FullAdder_187_io_s),
    .io_co(FullAdder_187_io_co)
  );
  FullAdder FullAdder_188 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_188_io_a),
    .io_b(FullAdder_188_io_b),
    .io_ci(FullAdder_188_io_ci),
    .io_s(FullAdder_188_io_s),
    .io_co(FullAdder_188_io_co)
  );
  FullAdder FullAdder_189 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_189_io_a),
    .io_b(FullAdder_189_io_b),
    .io_ci(FullAdder_189_io_ci),
    .io_s(FullAdder_189_io_s),
    .io_co(FullAdder_189_io_co)
  );
  FullAdder FullAdder_190 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_190_io_a),
    .io_b(FullAdder_190_io_b),
    .io_ci(FullAdder_190_io_ci),
    .io_s(FullAdder_190_io_s),
    .io_co(FullAdder_190_io_co)
  );
  FullAdder FullAdder_191 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_191_io_a),
    .io_b(FullAdder_191_io_b),
    .io_ci(FullAdder_191_io_ci),
    .io_s(FullAdder_191_io_s),
    .io_co(FullAdder_191_io_co)
  );
  FullAdder FullAdder_192 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_192_io_a),
    .io_b(FullAdder_192_io_b),
    .io_ci(FullAdder_192_io_ci),
    .io_s(FullAdder_192_io_s),
    .io_co(FullAdder_192_io_co)
  );
  FullAdder FullAdder_193 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_193_io_a),
    .io_b(FullAdder_193_io_b),
    .io_ci(FullAdder_193_io_ci),
    .io_s(FullAdder_193_io_s),
    .io_co(FullAdder_193_io_co)
  );
  FullAdder FullAdder_194 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_194_io_a),
    .io_b(FullAdder_194_io_b),
    .io_ci(FullAdder_194_io_ci),
    .io_s(FullAdder_194_io_s),
    .io_co(FullAdder_194_io_co)
  );
  FullAdder FullAdder_195 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_195_io_a),
    .io_b(FullAdder_195_io_b),
    .io_ci(FullAdder_195_io_ci),
    .io_s(FullAdder_195_io_s),
    .io_co(FullAdder_195_io_co)
  );
  FullAdder FullAdder_196 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_196_io_a),
    .io_b(FullAdder_196_io_b),
    .io_ci(FullAdder_196_io_ci),
    .io_s(FullAdder_196_io_s),
    .io_co(FullAdder_196_io_co)
  );
  FullAdder FullAdder_197 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_197_io_a),
    .io_b(FullAdder_197_io_b),
    .io_ci(FullAdder_197_io_ci),
    .io_s(FullAdder_197_io_s),
    .io_co(FullAdder_197_io_co)
  );
  HalfAdder HalfAdder_8 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_8_io_a),
    .io_b(HalfAdder_8_io_b),
    .io_s(HalfAdder_8_io_s),
    .io_co(HalfAdder_8_io_co)
  );
  FullAdder FullAdder_198 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_198_io_a),
    .io_b(FullAdder_198_io_b),
    .io_ci(FullAdder_198_io_ci),
    .io_s(FullAdder_198_io_s),
    .io_co(FullAdder_198_io_co)
  );
  FullAdder FullAdder_199 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_199_io_a),
    .io_b(FullAdder_199_io_b),
    .io_ci(FullAdder_199_io_ci),
    .io_s(FullAdder_199_io_s),
    .io_co(FullAdder_199_io_co)
  );
  FullAdder FullAdder_200 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_200_io_a),
    .io_b(FullAdder_200_io_b),
    .io_ci(FullAdder_200_io_ci),
    .io_s(FullAdder_200_io_s),
    .io_co(FullAdder_200_io_co)
  );
  FullAdder FullAdder_201 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_201_io_a),
    .io_b(FullAdder_201_io_b),
    .io_ci(FullAdder_201_io_ci),
    .io_s(FullAdder_201_io_s),
    .io_co(FullAdder_201_io_co)
  );
  FullAdder FullAdder_202 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_202_io_a),
    .io_b(FullAdder_202_io_b),
    .io_ci(FullAdder_202_io_ci),
    .io_s(FullAdder_202_io_s),
    .io_co(FullAdder_202_io_co)
  );
  FullAdder FullAdder_203 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_203_io_a),
    .io_b(FullAdder_203_io_b),
    .io_ci(FullAdder_203_io_ci),
    .io_s(FullAdder_203_io_s),
    .io_co(FullAdder_203_io_co)
  );
  FullAdder FullAdder_204 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_204_io_a),
    .io_b(FullAdder_204_io_b),
    .io_ci(FullAdder_204_io_ci),
    .io_s(FullAdder_204_io_s),
    .io_co(FullAdder_204_io_co)
  );
  FullAdder FullAdder_205 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_205_io_a),
    .io_b(FullAdder_205_io_b),
    .io_ci(FullAdder_205_io_ci),
    .io_s(FullAdder_205_io_s),
    .io_co(FullAdder_205_io_co)
  );
  FullAdder FullAdder_206 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_206_io_a),
    .io_b(FullAdder_206_io_b),
    .io_ci(FullAdder_206_io_ci),
    .io_s(FullAdder_206_io_s),
    .io_co(FullAdder_206_io_co)
  );
  FullAdder FullAdder_207 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_207_io_a),
    .io_b(FullAdder_207_io_b),
    .io_ci(FullAdder_207_io_ci),
    .io_s(FullAdder_207_io_s),
    .io_co(FullAdder_207_io_co)
  );
  FullAdder FullAdder_208 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_208_io_a),
    .io_b(FullAdder_208_io_b),
    .io_ci(FullAdder_208_io_ci),
    .io_s(FullAdder_208_io_s),
    .io_co(FullAdder_208_io_co)
  );
  FullAdder FullAdder_209 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_209_io_a),
    .io_b(FullAdder_209_io_b),
    .io_ci(FullAdder_209_io_ci),
    .io_s(FullAdder_209_io_s),
    .io_co(FullAdder_209_io_co)
  );
  FullAdder FullAdder_210 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_210_io_a),
    .io_b(FullAdder_210_io_b),
    .io_ci(FullAdder_210_io_ci),
    .io_s(FullAdder_210_io_s),
    .io_co(FullAdder_210_io_co)
  );
  FullAdder FullAdder_211 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_211_io_a),
    .io_b(FullAdder_211_io_b),
    .io_ci(FullAdder_211_io_ci),
    .io_s(FullAdder_211_io_s),
    .io_co(FullAdder_211_io_co)
  );
  FullAdder FullAdder_212 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_212_io_a),
    .io_b(FullAdder_212_io_b),
    .io_ci(FullAdder_212_io_ci),
    .io_s(FullAdder_212_io_s),
    .io_co(FullAdder_212_io_co)
  );
  FullAdder FullAdder_213 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_213_io_a),
    .io_b(FullAdder_213_io_b),
    .io_ci(FullAdder_213_io_ci),
    .io_s(FullAdder_213_io_s),
    .io_co(FullAdder_213_io_co)
  );
  FullAdder FullAdder_214 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_214_io_a),
    .io_b(FullAdder_214_io_b),
    .io_ci(FullAdder_214_io_ci),
    .io_s(FullAdder_214_io_s),
    .io_co(FullAdder_214_io_co)
  );
  FullAdder FullAdder_215 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_215_io_a),
    .io_b(FullAdder_215_io_b),
    .io_ci(FullAdder_215_io_ci),
    .io_s(FullAdder_215_io_s),
    .io_co(FullAdder_215_io_co)
  );
  FullAdder FullAdder_216 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_216_io_a),
    .io_b(FullAdder_216_io_b),
    .io_ci(FullAdder_216_io_ci),
    .io_s(FullAdder_216_io_s),
    .io_co(FullAdder_216_io_co)
  );
  FullAdder FullAdder_217 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_217_io_a),
    .io_b(FullAdder_217_io_b),
    .io_ci(FullAdder_217_io_ci),
    .io_s(FullAdder_217_io_s),
    .io_co(FullAdder_217_io_co)
  );
  FullAdder FullAdder_218 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_218_io_a),
    .io_b(FullAdder_218_io_b),
    .io_ci(FullAdder_218_io_ci),
    .io_s(FullAdder_218_io_s),
    .io_co(FullAdder_218_io_co)
  );
  FullAdder FullAdder_219 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_219_io_a),
    .io_b(FullAdder_219_io_b),
    .io_ci(FullAdder_219_io_ci),
    .io_s(FullAdder_219_io_s),
    .io_co(FullAdder_219_io_co)
  );
  FullAdder FullAdder_220 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_220_io_a),
    .io_b(FullAdder_220_io_b),
    .io_ci(FullAdder_220_io_ci),
    .io_s(FullAdder_220_io_s),
    .io_co(FullAdder_220_io_co)
  );
  FullAdder FullAdder_221 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_221_io_a),
    .io_b(FullAdder_221_io_b),
    .io_ci(FullAdder_221_io_ci),
    .io_s(FullAdder_221_io_s),
    .io_co(FullAdder_221_io_co)
  );
  FullAdder FullAdder_222 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_222_io_a),
    .io_b(FullAdder_222_io_b),
    .io_ci(FullAdder_222_io_ci),
    .io_s(FullAdder_222_io_s),
    .io_co(FullAdder_222_io_co)
  );
  FullAdder FullAdder_223 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_223_io_a),
    .io_b(FullAdder_223_io_b),
    .io_ci(FullAdder_223_io_ci),
    .io_s(FullAdder_223_io_s),
    .io_co(FullAdder_223_io_co)
  );
  FullAdder FullAdder_224 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_224_io_a),
    .io_b(FullAdder_224_io_b),
    .io_ci(FullAdder_224_io_ci),
    .io_s(FullAdder_224_io_s),
    .io_co(FullAdder_224_io_co)
  );
  FullAdder FullAdder_225 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_225_io_a),
    .io_b(FullAdder_225_io_b),
    .io_ci(FullAdder_225_io_ci),
    .io_s(FullAdder_225_io_s),
    .io_co(FullAdder_225_io_co)
  );
  FullAdder FullAdder_226 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_226_io_a),
    .io_b(FullAdder_226_io_b),
    .io_ci(FullAdder_226_io_ci),
    .io_s(FullAdder_226_io_s),
    .io_co(FullAdder_226_io_co)
  );
  FullAdder FullAdder_227 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_227_io_a),
    .io_b(FullAdder_227_io_b),
    .io_ci(FullAdder_227_io_ci),
    .io_s(FullAdder_227_io_s),
    .io_co(FullAdder_227_io_co)
  );
  FullAdder FullAdder_228 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_228_io_a),
    .io_b(FullAdder_228_io_b),
    .io_ci(FullAdder_228_io_ci),
    .io_s(FullAdder_228_io_s),
    .io_co(FullAdder_228_io_co)
  );
  FullAdder FullAdder_229 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_229_io_a),
    .io_b(FullAdder_229_io_b),
    .io_ci(FullAdder_229_io_ci),
    .io_s(FullAdder_229_io_s),
    .io_co(FullAdder_229_io_co)
  );
  FullAdder FullAdder_230 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_230_io_a),
    .io_b(FullAdder_230_io_b),
    .io_ci(FullAdder_230_io_ci),
    .io_s(FullAdder_230_io_s),
    .io_co(FullAdder_230_io_co)
  );
  FullAdder FullAdder_231 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_231_io_a),
    .io_b(FullAdder_231_io_b),
    .io_ci(FullAdder_231_io_ci),
    .io_s(FullAdder_231_io_s),
    .io_co(FullAdder_231_io_co)
  );
  FullAdder FullAdder_232 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_232_io_a),
    .io_b(FullAdder_232_io_b),
    .io_ci(FullAdder_232_io_ci),
    .io_s(FullAdder_232_io_s),
    .io_co(FullAdder_232_io_co)
  );
  FullAdder FullAdder_233 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_233_io_a),
    .io_b(FullAdder_233_io_b),
    .io_ci(FullAdder_233_io_ci),
    .io_s(FullAdder_233_io_s),
    .io_co(FullAdder_233_io_co)
  );
  HalfAdder HalfAdder_9 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_9_io_a),
    .io_b(HalfAdder_9_io_b),
    .io_s(HalfAdder_9_io_s),
    .io_co(HalfAdder_9_io_co)
  );
  FullAdder FullAdder_234 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_234_io_a),
    .io_b(FullAdder_234_io_b),
    .io_ci(FullAdder_234_io_ci),
    .io_s(FullAdder_234_io_s),
    .io_co(FullAdder_234_io_co)
  );
  FullAdder FullAdder_235 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_235_io_a),
    .io_b(FullAdder_235_io_b),
    .io_ci(FullAdder_235_io_ci),
    .io_s(FullAdder_235_io_s),
    .io_co(FullAdder_235_io_co)
  );
  FullAdder FullAdder_236 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_236_io_a),
    .io_b(FullAdder_236_io_b),
    .io_ci(FullAdder_236_io_ci),
    .io_s(FullAdder_236_io_s),
    .io_co(FullAdder_236_io_co)
  );
  FullAdder FullAdder_237 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_237_io_a),
    .io_b(FullAdder_237_io_b),
    .io_ci(FullAdder_237_io_ci),
    .io_s(FullAdder_237_io_s),
    .io_co(FullAdder_237_io_co)
  );
  FullAdder FullAdder_238 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_238_io_a),
    .io_b(FullAdder_238_io_b),
    .io_ci(FullAdder_238_io_ci),
    .io_s(FullAdder_238_io_s),
    .io_co(FullAdder_238_io_co)
  );
  FullAdder FullAdder_239 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_239_io_a),
    .io_b(FullAdder_239_io_b),
    .io_ci(FullAdder_239_io_ci),
    .io_s(FullAdder_239_io_s),
    .io_co(FullAdder_239_io_co)
  );
  FullAdder FullAdder_240 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_240_io_a),
    .io_b(FullAdder_240_io_b),
    .io_ci(FullAdder_240_io_ci),
    .io_s(FullAdder_240_io_s),
    .io_co(FullAdder_240_io_co)
  );
  FullAdder FullAdder_241 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_241_io_a),
    .io_b(FullAdder_241_io_b),
    .io_ci(FullAdder_241_io_ci),
    .io_s(FullAdder_241_io_s),
    .io_co(FullAdder_241_io_co)
  );
  FullAdder FullAdder_242 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_242_io_a),
    .io_b(FullAdder_242_io_b),
    .io_ci(FullAdder_242_io_ci),
    .io_s(FullAdder_242_io_s),
    .io_co(FullAdder_242_io_co)
  );
  FullAdder FullAdder_243 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_243_io_a),
    .io_b(FullAdder_243_io_b),
    .io_ci(FullAdder_243_io_ci),
    .io_s(FullAdder_243_io_s),
    .io_co(FullAdder_243_io_co)
  );
  FullAdder FullAdder_244 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_244_io_a),
    .io_b(FullAdder_244_io_b),
    .io_ci(FullAdder_244_io_ci),
    .io_s(FullAdder_244_io_s),
    .io_co(FullAdder_244_io_co)
  );
  FullAdder FullAdder_245 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_245_io_a),
    .io_b(FullAdder_245_io_b),
    .io_ci(FullAdder_245_io_ci),
    .io_s(FullAdder_245_io_s),
    .io_co(FullAdder_245_io_co)
  );
  FullAdder FullAdder_246 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_246_io_a),
    .io_b(FullAdder_246_io_b),
    .io_ci(FullAdder_246_io_ci),
    .io_s(FullAdder_246_io_s),
    .io_co(FullAdder_246_io_co)
  );
  FullAdder FullAdder_247 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_247_io_a),
    .io_b(FullAdder_247_io_b),
    .io_ci(FullAdder_247_io_ci),
    .io_s(FullAdder_247_io_s),
    .io_co(FullAdder_247_io_co)
  );
  FullAdder FullAdder_248 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_248_io_a),
    .io_b(FullAdder_248_io_b),
    .io_ci(FullAdder_248_io_ci),
    .io_s(FullAdder_248_io_s),
    .io_co(FullAdder_248_io_co)
  );
  FullAdder FullAdder_249 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_249_io_a),
    .io_b(FullAdder_249_io_b),
    .io_ci(FullAdder_249_io_ci),
    .io_s(FullAdder_249_io_s),
    .io_co(FullAdder_249_io_co)
  );
  FullAdder FullAdder_250 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_250_io_a),
    .io_b(FullAdder_250_io_b),
    .io_ci(FullAdder_250_io_ci),
    .io_s(FullAdder_250_io_s),
    .io_co(FullAdder_250_io_co)
  );
  FullAdder FullAdder_251 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_251_io_a),
    .io_b(FullAdder_251_io_b),
    .io_ci(FullAdder_251_io_ci),
    .io_s(FullAdder_251_io_s),
    .io_co(FullAdder_251_io_co)
  );
  FullAdder FullAdder_252 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_252_io_a),
    .io_b(FullAdder_252_io_b),
    .io_ci(FullAdder_252_io_ci),
    .io_s(FullAdder_252_io_s),
    .io_co(FullAdder_252_io_co)
  );
  FullAdder FullAdder_253 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_253_io_a),
    .io_b(FullAdder_253_io_b),
    .io_ci(FullAdder_253_io_ci),
    .io_s(FullAdder_253_io_s),
    .io_co(FullAdder_253_io_co)
  );
  FullAdder FullAdder_254 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_254_io_a),
    .io_b(FullAdder_254_io_b),
    .io_ci(FullAdder_254_io_ci),
    .io_s(FullAdder_254_io_s),
    .io_co(FullAdder_254_io_co)
  );
  FullAdder FullAdder_255 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_255_io_a),
    .io_b(FullAdder_255_io_b),
    .io_ci(FullAdder_255_io_ci),
    .io_s(FullAdder_255_io_s),
    .io_co(FullAdder_255_io_co)
  );
  FullAdder FullAdder_256 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_256_io_a),
    .io_b(FullAdder_256_io_b),
    .io_ci(FullAdder_256_io_ci),
    .io_s(FullAdder_256_io_s),
    .io_co(FullAdder_256_io_co)
  );
  FullAdder FullAdder_257 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_257_io_a),
    .io_b(FullAdder_257_io_b),
    .io_ci(FullAdder_257_io_ci),
    .io_s(FullAdder_257_io_s),
    .io_co(FullAdder_257_io_co)
  );
  FullAdder FullAdder_258 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_258_io_a),
    .io_b(FullAdder_258_io_b),
    .io_ci(FullAdder_258_io_ci),
    .io_s(FullAdder_258_io_s),
    .io_co(FullAdder_258_io_co)
  );
  FullAdder FullAdder_259 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_259_io_a),
    .io_b(FullAdder_259_io_b),
    .io_ci(FullAdder_259_io_ci),
    .io_s(FullAdder_259_io_s),
    .io_co(FullAdder_259_io_co)
  );
  FullAdder FullAdder_260 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_260_io_a),
    .io_b(FullAdder_260_io_b),
    .io_ci(FullAdder_260_io_ci),
    .io_s(FullAdder_260_io_s),
    .io_co(FullAdder_260_io_co)
  );
  FullAdder FullAdder_261 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_261_io_a),
    .io_b(FullAdder_261_io_b),
    .io_ci(FullAdder_261_io_ci),
    .io_s(FullAdder_261_io_s),
    .io_co(FullAdder_261_io_co)
  );
  FullAdder FullAdder_262 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_262_io_a),
    .io_b(FullAdder_262_io_b),
    .io_ci(FullAdder_262_io_ci),
    .io_s(FullAdder_262_io_s),
    .io_co(FullAdder_262_io_co)
  );
  FullAdder FullAdder_263 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_263_io_a),
    .io_b(FullAdder_263_io_b),
    .io_ci(FullAdder_263_io_ci),
    .io_s(FullAdder_263_io_s),
    .io_co(FullAdder_263_io_co)
  );
  FullAdder FullAdder_264 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_264_io_a),
    .io_b(FullAdder_264_io_b),
    .io_ci(FullAdder_264_io_ci),
    .io_s(FullAdder_264_io_s),
    .io_co(FullAdder_264_io_co)
  );
  FullAdder FullAdder_265 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_265_io_a),
    .io_b(FullAdder_265_io_b),
    .io_ci(FullAdder_265_io_ci),
    .io_s(FullAdder_265_io_s),
    .io_co(FullAdder_265_io_co)
  );
  FullAdder FullAdder_266 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_266_io_a),
    .io_b(FullAdder_266_io_b),
    .io_ci(FullAdder_266_io_ci),
    .io_s(FullAdder_266_io_s),
    .io_co(FullAdder_266_io_co)
  );
  FullAdder FullAdder_267 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_267_io_a),
    .io_b(FullAdder_267_io_b),
    .io_ci(FullAdder_267_io_ci),
    .io_s(FullAdder_267_io_s),
    .io_co(FullAdder_267_io_co)
  );
  FullAdder FullAdder_268 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_268_io_a),
    .io_b(FullAdder_268_io_b),
    .io_ci(FullAdder_268_io_ci),
    .io_s(FullAdder_268_io_s),
    .io_co(FullAdder_268_io_co)
  );
  FullAdder FullAdder_269 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_269_io_a),
    .io_b(FullAdder_269_io_b),
    .io_ci(FullAdder_269_io_ci),
    .io_s(FullAdder_269_io_s),
    .io_co(FullAdder_269_io_co)
  );
  FullAdder FullAdder_270 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_270_io_a),
    .io_b(FullAdder_270_io_b),
    .io_ci(FullAdder_270_io_ci),
    .io_s(FullAdder_270_io_s),
    .io_co(FullAdder_270_io_co)
  );
  FullAdder FullAdder_271 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_271_io_a),
    .io_b(FullAdder_271_io_b),
    .io_ci(FullAdder_271_io_ci),
    .io_s(FullAdder_271_io_s),
    .io_co(FullAdder_271_io_co)
  );
  FullAdder FullAdder_272 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_272_io_a),
    .io_b(FullAdder_272_io_b),
    .io_ci(FullAdder_272_io_ci),
    .io_s(FullAdder_272_io_s),
    .io_co(FullAdder_272_io_co)
  );
  HalfAdder HalfAdder_10 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_10_io_a),
    .io_b(HalfAdder_10_io_b),
    .io_s(HalfAdder_10_io_s),
    .io_co(HalfAdder_10_io_co)
  );
  FullAdder FullAdder_273 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_273_io_a),
    .io_b(FullAdder_273_io_b),
    .io_ci(FullAdder_273_io_ci),
    .io_s(FullAdder_273_io_s),
    .io_co(FullAdder_273_io_co)
  );
  FullAdder FullAdder_274 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_274_io_a),
    .io_b(FullAdder_274_io_b),
    .io_ci(FullAdder_274_io_ci),
    .io_s(FullAdder_274_io_s),
    .io_co(FullAdder_274_io_co)
  );
  FullAdder FullAdder_275 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_275_io_a),
    .io_b(FullAdder_275_io_b),
    .io_ci(FullAdder_275_io_ci),
    .io_s(FullAdder_275_io_s),
    .io_co(FullAdder_275_io_co)
  );
  FullAdder FullAdder_276 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_276_io_a),
    .io_b(FullAdder_276_io_b),
    .io_ci(FullAdder_276_io_ci),
    .io_s(FullAdder_276_io_s),
    .io_co(FullAdder_276_io_co)
  );
  FullAdder FullAdder_277 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_277_io_a),
    .io_b(FullAdder_277_io_b),
    .io_ci(FullAdder_277_io_ci),
    .io_s(FullAdder_277_io_s),
    .io_co(FullAdder_277_io_co)
  );
  FullAdder FullAdder_278 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_278_io_a),
    .io_b(FullAdder_278_io_b),
    .io_ci(FullAdder_278_io_ci),
    .io_s(FullAdder_278_io_s),
    .io_co(FullAdder_278_io_co)
  );
  FullAdder FullAdder_279 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_279_io_a),
    .io_b(FullAdder_279_io_b),
    .io_ci(FullAdder_279_io_ci),
    .io_s(FullAdder_279_io_s),
    .io_co(FullAdder_279_io_co)
  );
  FullAdder FullAdder_280 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_280_io_a),
    .io_b(FullAdder_280_io_b),
    .io_ci(FullAdder_280_io_ci),
    .io_s(FullAdder_280_io_s),
    .io_co(FullAdder_280_io_co)
  );
  FullAdder FullAdder_281 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_281_io_a),
    .io_b(FullAdder_281_io_b),
    .io_ci(FullAdder_281_io_ci),
    .io_s(FullAdder_281_io_s),
    .io_co(FullAdder_281_io_co)
  );
  FullAdder FullAdder_282 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_282_io_a),
    .io_b(FullAdder_282_io_b),
    .io_ci(FullAdder_282_io_ci),
    .io_s(FullAdder_282_io_s),
    .io_co(FullAdder_282_io_co)
  );
  FullAdder FullAdder_283 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_283_io_a),
    .io_b(FullAdder_283_io_b),
    .io_ci(FullAdder_283_io_ci),
    .io_s(FullAdder_283_io_s),
    .io_co(FullAdder_283_io_co)
  );
  FullAdder FullAdder_284 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_284_io_a),
    .io_b(FullAdder_284_io_b),
    .io_ci(FullAdder_284_io_ci),
    .io_s(FullAdder_284_io_s),
    .io_co(FullAdder_284_io_co)
  );
  FullAdder FullAdder_285 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_285_io_a),
    .io_b(FullAdder_285_io_b),
    .io_ci(FullAdder_285_io_ci),
    .io_s(FullAdder_285_io_s),
    .io_co(FullAdder_285_io_co)
  );
  FullAdder FullAdder_286 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_286_io_a),
    .io_b(FullAdder_286_io_b),
    .io_ci(FullAdder_286_io_ci),
    .io_s(FullAdder_286_io_s),
    .io_co(FullAdder_286_io_co)
  );
  FullAdder FullAdder_287 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_287_io_a),
    .io_b(FullAdder_287_io_b),
    .io_ci(FullAdder_287_io_ci),
    .io_s(FullAdder_287_io_s),
    .io_co(FullAdder_287_io_co)
  );
  FullAdder FullAdder_288 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_288_io_a),
    .io_b(FullAdder_288_io_b),
    .io_ci(FullAdder_288_io_ci),
    .io_s(FullAdder_288_io_s),
    .io_co(FullAdder_288_io_co)
  );
  FullAdder FullAdder_289 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_289_io_a),
    .io_b(FullAdder_289_io_b),
    .io_ci(FullAdder_289_io_ci),
    .io_s(FullAdder_289_io_s),
    .io_co(FullAdder_289_io_co)
  );
  FullAdder FullAdder_290 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_290_io_a),
    .io_b(FullAdder_290_io_b),
    .io_ci(FullAdder_290_io_ci),
    .io_s(FullAdder_290_io_s),
    .io_co(FullAdder_290_io_co)
  );
  FullAdder FullAdder_291 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_291_io_a),
    .io_b(FullAdder_291_io_b),
    .io_ci(FullAdder_291_io_ci),
    .io_s(FullAdder_291_io_s),
    .io_co(FullAdder_291_io_co)
  );
  FullAdder FullAdder_292 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_292_io_a),
    .io_b(FullAdder_292_io_b),
    .io_ci(FullAdder_292_io_ci),
    .io_s(FullAdder_292_io_s),
    .io_co(FullAdder_292_io_co)
  );
  FullAdder FullAdder_293 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_293_io_a),
    .io_b(FullAdder_293_io_b),
    .io_ci(FullAdder_293_io_ci),
    .io_s(FullAdder_293_io_s),
    .io_co(FullAdder_293_io_co)
  );
  FullAdder FullAdder_294 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_294_io_a),
    .io_b(FullAdder_294_io_b),
    .io_ci(FullAdder_294_io_ci),
    .io_s(FullAdder_294_io_s),
    .io_co(FullAdder_294_io_co)
  );
  FullAdder FullAdder_295 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_295_io_a),
    .io_b(FullAdder_295_io_b),
    .io_ci(FullAdder_295_io_ci),
    .io_s(FullAdder_295_io_s),
    .io_co(FullAdder_295_io_co)
  );
  FullAdder FullAdder_296 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_296_io_a),
    .io_b(FullAdder_296_io_b),
    .io_ci(FullAdder_296_io_ci),
    .io_s(FullAdder_296_io_s),
    .io_co(FullAdder_296_io_co)
  );
  FullAdder FullAdder_297 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_297_io_a),
    .io_b(FullAdder_297_io_b),
    .io_ci(FullAdder_297_io_ci),
    .io_s(FullAdder_297_io_s),
    .io_co(FullAdder_297_io_co)
  );
  FullAdder FullAdder_298 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_298_io_a),
    .io_b(FullAdder_298_io_b),
    .io_ci(FullAdder_298_io_ci),
    .io_s(FullAdder_298_io_s),
    .io_co(FullAdder_298_io_co)
  );
  FullAdder FullAdder_299 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_299_io_a),
    .io_b(FullAdder_299_io_b),
    .io_ci(FullAdder_299_io_ci),
    .io_s(FullAdder_299_io_s),
    .io_co(FullAdder_299_io_co)
  );
  FullAdder FullAdder_300 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_300_io_a),
    .io_b(FullAdder_300_io_b),
    .io_ci(FullAdder_300_io_ci),
    .io_s(FullAdder_300_io_s),
    .io_co(FullAdder_300_io_co)
  );
  FullAdder FullAdder_301 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_301_io_a),
    .io_b(FullAdder_301_io_b),
    .io_ci(FullAdder_301_io_ci),
    .io_s(FullAdder_301_io_s),
    .io_co(FullAdder_301_io_co)
  );
  FullAdder FullAdder_302 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_302_io_a),
    .io_b(FullAdder_302_io_b),
    .io_ci(FullAdder_302_io_ci),
    .io_s(FullAdder_302_io_s),
    .io_co(FullAdder_302_io_co)
  );
  FullAdder FullAdder_303 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_303_io_a),
    .io_b(FullAdder_303_io_b),
    .io_ci(FullAdder_303_io_ci),
    .io_s(FullAdder_303_io_s),
    .io_co(FullAdder_303_io_co)
  );
  FullAdder FullAdder_304 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_304_io_a),
    .io_b(FullAdder_304_io_b),
    .io_ci(FullAdder_304_io_ci),
    .io_s(FullAdder_304_io_s),
    .io_co(FullAdder_304_io_co)
  );
  FullAdder FullAdder_305 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_305_io_a),
    .io_b(FullAdder_305_io_b),
    .io_ci(FullAdder_305_io_ci),
    .io_s(FullAdder_305_io_s),
    .io_co(FullAdder_305_io_co)
  );
  FullAdder FullAdder_306 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_306_io_a),
    .io_b(FullAdder_306_io_b),
    .io_ci(FullAdder_306_io_ci),
    .io_s(FullAdder_306_io_s),
    .io_co(FullAdder_306_io_co)
  );
  FullAdder FullAdder_307 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_307_io_a),
    .io_b(FullAdder_307_io_b),
    .io_ci(FullAdder_307_io_ci),
    .io_s(FullAdder_307_io_s),
    .io_co(FullAdder_307_io_co)
  );
  FullAdder FullAdder_308 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_308_io_a),
    .io_b(FullAdder_308_io_b),
    .io_ci(FullAdder_308_io_ci),
    .io_s(FullAdder_308_io_s),
    .io_co(FullAdder_308_io_co)
  );
  FullAdder FullAdder_309 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_309_io_a),
    .io_b(FullAdder_309_io_b),
    .io_ci(FullAdder_309_io_ci),
    .io_s(FullAdder_309_io_s),
    .io_co(FullAdder_309_io_co)
  );
  FullAdder FullAdder_310 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_310_io_a),
    .io_b(FullAdder_310_io_b),
    .io_ci(FullAdder_310_io_ci),
    .io_s(FullAdder_310_io_s),
    .io_co(FullAdder_310_io_co)
  );
  FullAdder FullAdder_311 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_311_io_a),
    .io_b(FullAdder_311_io_b),
    .io_ci(FullAdder_311_io_ci),
    .io_s(FullAdder_311_io_s),
    .io_co(FullAdder_311_io_co)
  );
  FullAdder FullAdder_312 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_312_io_a),
    .io_b(FullAdder_312_io_b),
    .io_ci(FullAdder_312_io_ci),
    .io_s(FullAdder_312_io_s),
    .io_co(FullAdder_312_io_co)
  );
  FullAdder FullAdder_313 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_313_io_a),
    .io_b(FullAdder_313_io_b),
    .io_ci(FullAdder_313_io_ci),
    .io_s(FullAdder_313_io_s),
    .io_co(FullAdder_313_io_co)
  );
  FullAdder FullAdder_314 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_314_io_a),
    .io_b(FullAdder_314_io_b),
    .io_ci(FullAdder_314_io_ci),
    .io_s(FullAdder_314_io_s),
    .io_co(FullAdder_314_io_co)
  );
  HalfAdder HalfAdder_11 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_11_io_a),
    .io_b(HalfAdder_11_io_b),
    .io_s(HalfAdder_11_io_s),
    .io_co(HalfAdder_11_io_co)
  );
  FullAdder FullAdder_315 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_315_io_a),
    .io_b(FullAdder_315_io_b),
    .io_ci(FullAdder_315_io_ci),
    .io_s(FullAdder_315_io_s),
    .io_co(FullAdder_315_io_co)
  );
  FullAdder FullAdder_316 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_316_io_a),
    .io_b(FullAdder_316_io_b),
    .io_ci(FullAdder_316_io_ci),
    .io_s(FullAdder_316_io_s),
    .io_co(FullAdder_316_io_co)
  );
  FullAdder FullAdder_317 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_317_io_a),
    .io_b(FullAdder_317_io_b),
    .io_ci(FullAdder_317_io_ci),
    .io_s(FullAdder_317_io_s),
    .io_co(FullAdder_317_io_co)
  );
  FullAdder FullAdder_318 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_318_io_a),
    .io_b(FullAdder_318_io_b),
    .io_ci(FullAdder_318_io_ci),
    .io_s(FullAdder_318_io_s),
    .io_co(FullAdder_318_io_co)
  );
  FullAdder FullAdder_319 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_319_io_a),
    .io_b(FullAdder_319_io_b),
    .io_ci(FullAdder_319_io_ci),
    .io_s(FullAdder_319_io_s),
    .io_co(FullAdder_319_io_co)
  );
  FullAdder FullAdder_320 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_320_io_a),
    .io_b(FullAdder_320_io_b),
    .io_ci(FullAdder_320_io_ci),
    .io_s(FullAdder_320_io_s),
    .io_co(FullAdder_320_io_co)
  );
  FullAdder FullAdder_321 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_321_io_a),
    .io_b(FullAdder_321_io_b),
    .io_ci(FullAdder_321_io_ci),
    .io_s(FullAdder_321_io_s),
    .io_co(FullAdder_321_io_co)
  );
  FullAdder FullAdder_322 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_322_io_a),
    .io_b(FullAdder_322_io_b),
    .io_ci(FullAdder_322_io_ci),
    .io_s(FullAdder_322_io_s),
    .io_co(FullAdder_322_io_co)
  );
  FullAdder FullAdder_323 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_323_io_a),
    .io_b(FullAdder_323_io_b),
    .io_ci(FullAdder_323_io_ci),
    .io_s(FullAdder_323_io_s),
    .io_co(FullAdder_323_io_co)
  );
  FullAdder FullAdder_324 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_324_io_a),
    .io_b(FullAdder_324_io_b),
    .io_ci(FullAdder_324_io_ci),
    .io_s(FullAdder_324_io_s),
    .io_co(FullAdder_324_io_co)
  );
  FullAdder FullAdder_325 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_325_io_a),
    .io_b(FullAdder_325_io_b),
    .io_ci(FullAdder_325_io_ci),
    .io_s(FullAdder_325_io_s),
    .io_co(FullAdder_325_io_co)
  );
  FullAdder FullAdder_326 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_326_io_a),
    .io_b(FullAdder_326_io_b),
    .io_ci(FullAdder_326_io_ci),
    .io_s(FullAdder_326_io_s),
    .io_co(FullAdder_326_io_co)
  );
  FullAdder FullAdder_327 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_327_io_a),
    .io_b(FullAdder_327_io_b),
    .io_ci(FullAdder_327_io_ci),
    .io_s(FullAdder_327_io_s),
    .io_co(FullAdder_327_io_co)
  );
  FullAdder FullAdder_328 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_328_io_a),
    .io_b(FullAdder_328_io_b),
    .io_ci(FullAdder_328_io_ci),
    .io_s(FullAdder_328_io_s),
    .io_co(FullAdder_328_io_co)
  );
  FullAdder FullAdder_329 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_329_io_a),
    .io_b(FullAdder_329_io_b),
    .io_ci(FullAdder_329_io_ci),
    .io_s(FullAdder_329_io_s),
    .io_co(FullAdder_329_io_co)
  );
  FullAdder FullAdder_330 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_330_io_a),
    .io_b(FullAdder_330_io_b),
    .io_ci(FullAdder_330_io_ci),
    .io_s(FullAdder_330_io_s),
    .io_co(FullAdder_330_io_co)
  );
  FullAdder FullAdder_331 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_331_io_a),
    .io_b(FullAdder_331_io_b),
    .io_ci(FullAdder_331_io_ci),
    .io_s(FullAdder_331_io_s),
    .io_co(FullAdder_331_io_co)
  );
  FullAdder FullAdder_332 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_332_io_a),
    .io_b(FullAdder_332_io_b),
    .io_ci(FullAdder_332_io_ci),
    .io_s(FullAdder_332_io_s),
    .io_co(FullAdder_332_io_co)
  );
  FullAdder FullAdder_333 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_333_io_a),
    .io_b(FullAdder_333_io_b),
    .io_ci(FullAdder_333_io_ci),
    .io_s(FullAdder_333_io_s),
    .io_co(FullAdder_333_io_co)
  );
  FullAdder FullAdder_334 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_334_io_a),
    .io_b(FullAdder_334_io_b),
    .io_ci(FullAdder_334_io_ci),
    .io_s(FullAdder_334_io_s),
    .io_co(FullAdder_334_io_co)
  );
  FullAdder FullAdder_335 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_335_io_a),
    .io_b(FullAdder_335_io_b),
    .io_ci(FullAdder_335_io_ci),
    .io_s(FullAdder_335_io_s),
    .io_co(FullAdder_335_io_co)
  );
  FullAdder FullAdder_336 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_336_io_a),
    .io_b(FullAdder_336_io_b),
    .io_ci(FullAdder_336_io_ci),
    .io_s(FullAdder_336_io_s),
    .io_co(FullAdder_336_io_co)
  );
  FullAdder FullAdder_337 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_337_io_a),
    .io_b(FullAdder_337_io_b),
    .io_ci(FullAdder_337_io_ci),
    .io_s(FullAdder_337_io_s),
    .io_co(FullAdder_337_io_co)
  );
  FullAdder FullAdder_338 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_338_io_a),
    .io_b(FullAdder_338_io_b),
    .io_ci(FullAdder_338_io_ci),
    .io_s(FullAdder_338_io_s),
    .io_co(FullAdder_338_io_co)
  );
  FullAdder FullAdder_339 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_339_io_a),
    .io_b(FullAdder_339_io_b),
    .io_ci(FullAdder_339_io_ci),
    .io_s(FullAdder_339_io_s),
    .io_co(FullAdder_339_io_co)
  );
  FullAdder FullAdder_340 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_340_io_a),
    .io_b(FullAdder_340_io_b),
    .io_ci(FullAdder_340_io_ci),
    .io_s(FullAdder_340_io_s),
    .io_co(FullAdder_340_io_co)
  );
  FullAdder FullAdder_341 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_341_io_a),
    .io_b(FullAdder_341_io_b),
    .io_ci(FullAdder_341_io_ci),
    .io_s(FullAdder_341_io_s),
    .io_co(FullAdder_341_io_co)
  );
  FullAdder FullAdder_342 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_342_io_a),
    .io_b(FullAdder_342_io_b),
    .io_ci(FullAdder_342_io_ci),
    .io_s(FullAdder_342_io_s),
    .io_co(FullAdder_342_io_co)
  );
  FullAdder FullAdder_343 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_343_io_a),
    .io_b(FullAdder_343_io_b),
    .io_ci(FullAdder_343_io_ci),
    .io_s(FullAdder_343_io_s),
    .io_co(FullAdder_343_io_co)
  );
  FullAdder FullAdder_344 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_344_io_a),
    .io_b(FullAdder_344_io_b),
    .io_ci(FullAdder_344_io_ci),
    .io_s(FullAdder_344_io_s),
    .io_co(FullAdder_344_io_co)
  );
  FullAdder FullAdder_345 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_345_io_a),
    .io_b(FullAdder_345_io_b),
    .io_ci(FullAdder_345_io_ci),
    .io_s(FullAdder_345_io_s),
    .io_co(FullAdder_345_io_co)
  );
  FullAdder FullAdder_346 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_346_io_a),
    .io_b(FullAdder_346_io_b),
    .io_ci(FullAdder_346_io_ci),
    .io_s(FullAdder_346_io_s),
    .io_co(FullAdder_346_io_co)
  );
  FullAdder FullAdder_347 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_347_io_a),
    .io_b(FullAdder_347_io_b),
    .io_ci(FullAdder_347_io_ci),
    .io_s(FullAdder_347_io_s),
    .io_co(FullAdder_347_io_co)
  );
  FullAdder FullAdder_348 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_348_io_a),
    .io_b(FullAdder_348_io_b),
    .io_ci(FullAdder_348_io_ci),
    .io_s(FullAdder_348_io_s),
    .io_co(FullAdder_348_io_co)
  );
  FullAdder FullAdder_349 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_349_io_a),
    .io_b(FullAdder_349_io_b),
    .io_ci(FullAdder_349_io_ci),
    .io_s(FullAdder_349_io_s),
    .io_co(FullAdder_349_io_co)
  );
  FullAdder FullAdder_350 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_350_io_a),
    .io_b(FullAdder_350_io_b),
    .io_ci(FullAdder_350_io_ci),
    .io_s(FullAdder_350_io_s),
    .io_co(FullAdder_350_io_co)
  );
  FullAdder FullAdder_351 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_351_io_a),
    .io_b(FullAdder_351_io_b),
    .io_ci(FullAdder_351_io_ci),
    .io_s(FullAdder_351_io_s),
    .io_co(FullAdder_351_io_co)
  );
  FullAdder FullAdder_352 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_352_io_a),
    .io_b(FullAdder_352_io_b),
    .io_ci(FullAdder_352_io_ci),
    .io_s(FullAdder_352_io_s),
    .io_co(FullAdder_352_io_co)
  );
  FullAdder FullAdder_353 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_353_io_a),
    .io_b(FullAdder_353_io_b),
    .io_ci(FullAdder_353_io_ci),
    .io_s(FullAdder_353_io_s),
    .io_co(FullAdder_353_io_co)
  );
  FullAdder FullAdder_354 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_354_io_a),
    .io_b(FullAdder_354_io_b),
    .io_ci(FullAdder_354_io_ci),
    .io_s(FullAdder_354_io_s),
    .io_co(FullAdder_354_io_co)
  );
  FullAdder FullAdder_355 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_355_io_a),
    .io_b(FullAdder_355_io_b),
    .io_ci(FullAdder_355_io_ci),
    .io_s(FullAdder_355_io_s),
    .io_co(FullAdder_355_io_co)
  );
  FullAdder FullAdder_356 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_356_io_a),
    .io_b(FullAdder_356_io_b),
    .io_ci(FullAdder_356_io_ci),
    .io_s(FullAdder_356_io_s),
    .io_co(FullAdder_356_io_co)
  );
  FullAdder FullAdder_357 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_357_io_a),
    .io_b(FullAdder_357_io_b),
    .io_ci(FullAdder_357_io_ci),
    .io_s(FullAdder_357_io_s),
    .io_co(FullAdder_357_io_co)
  );
  FullAdder FullAdder_358 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_358_io_a),
    .io_b(FullAdder_358_io_b),
    .io_ci(FullAdder_358_io_ci),
    .io_s(FullAdder_358_io_s),
    .io_co(FullAdder_358_io_co)
  );
  FullAdder FullAdder_359 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_359_io_a),
    .io_b(FullAdder_359_io_b),
    .io_ci(FullAdder_359_io_ci),
    .io_s(FullAdder_359_io_s),
    .io_co(FullAdder_359_io_co)
  );
  HalfAdder HalfAdder_12 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_12_io_a),
    .io_b(HalfAdder_12_io_b),
    .io_s(HalfAdder_12_io_s),
    .io_co(HalfAdder_12_io_co)
  );
  FullAdder FullAdder_360 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_360_io_a),
    .io_b(FullAdder_360_io_b),
    .io_ci(FullAdder_360_io_ci),
    .io_s(FullAdder_360_io_s),
    .io_co(FullAdder_360_io_co)
  );
  FullAdder FullAdder_361 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_361_io_a),
    .io_b(FullAdder_361_io_b),
    .io_ci(FullAdder_361_io_ci),
    .io_s(FullAdder_361_io_s),
    .io_co(FullAdder_361_io_co)
  );
  FullAdder FullAdder_362 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_362_io_a),
    .io_b(FullAdder_362_io_b),
    .io_ci(FullAdder_362_io_ci),
    .io_s(FullAdder_362_io_s),
    .io_co(FullAdder_362_io_co)
  );
  FullAdder FullAdder_363 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_363_io_a),
    .io_b(FullAdder_363_io_b),
    .io_ci(FullAdder_363_io_ci),
    .io_s(FullAdder_363_io_s),
    .io_co(FullAdder_363_io_co)
  );
  FullAdder FullAdder_364 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_364_io_a),
    .io_b(FullAdder_364_io_b),
    .io_ci(FullAdder_364_io_ci),
    .io_s(FullAdder_364_io_s),
    .io_co(FullAdder_364_io_co)
  );
  FullAdder FullAdder_365 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_365_io_a),
    .io_b(FullAdder_365_io_b),
    .io_ci(FullAdder_365_io_ci),
    .io_s(FullAdder_365_io_s),
    .io_co(FullAdder_365_io_co)
  );
  FullAdder FullAdder_366 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_366_io_a),
    .io_b(FullAdder_366_io_b),
    .io_ci(FullAdder_366_io_ci),
    .io_s(FullAdder_366_io_s),
    .io_co(FullAdder_366_io_co)
  );
  FullAdder FullAdder_367 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_367_io_a),
    .io_b(FullAdder_367_io_b),
    .io_ci(FullAdder_367_io_ci),
    .io_s(FullAdder_367_io_s),
    .io_co(FullAdder_367_io_co)
  );
  FullAdder FullAdder_368 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_368_io_a),
    .io_b(FullAdder_368_io_b),
    .io_ci(FullAdder_368_io_ci),
    .io_s(FullAdder_368_io_s),
    .io_co(FullAdder_368_io_co)
  );
  FullAdder FullAdder_369 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_369_io_a),
    .io_b(FullAdder_369_io_b),
    .io_ci(FullAdder_369_io_ci),
    .io_s(FullAdder_369_io_s),
    .io_co(FullAdder_369_io_co)
  );
  FullAdder FullAdder_370 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_370_io_a),
    .io_b(FullAdder_370_io_b),
    .io_ci(FullAdder_370_io_ci),
    .io_s(FullAdder_370_io_s),
    .io_co(FullAdder_370_io_co)
  );
  FullAdder FullAdder_371 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_371_io_a),
    .io_b(FullAdder_371_io_b),
    .io_ci(FullAdder_371_io_ci),
    .io_s(FullAdder_371_io_s),
    .io_co(FullAdder_371_io_co)
  );
  FullAdder FullAdder_372 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_372_io_a),
    .io_b(FullAdder_372_io_b),
    .io_ci(FullAdder_372_io_ci),
    .io_s(FullAdder_372_io_s),
    .io_co(FullAdder_372_io_co)
  );
  FullAdder FullAdder_373 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_373_io_a),
    .io_b(FullAdder_373_io_b),
    .io_ci(FullAdder_373_io_ci),
    .io_s(FullAdder_373_io_s),
    .io_co(FullAdder_373_io_co)
  );
  FullAdder FullAdder_374 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_374_io_a),
    .io_b(FullAdder_374_io_b),
    .io_ci(FullAdder_374_io_ci),
    .io_s(FullAdder_374_io_s),
    .io_co(FullAdder_374_io_co)
  );
  FullAdder FullAdder_375 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_375_io_a),
    .io_b(FullAdder_375_io_b),
    .io_ci(FullAdder_375_io_ci),
    .io_s(FullAdder_375_io_s),
    .io_co(FullAdder_375_io_co)
  );
  FullAdder FullAdder_376 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_376_io_a),
    .io_b(FullAdder_376_io_b),
    .io_ci(FullAdder_376_io_ci),
    .io_s(FullAdder_376_io_s),
    .io_co(FullAdder_376_io_co)
  );
  FullAdder FullAdder_377 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_377_io_a),
    .io_b(FullAdder_377_io_b),
    .io_ci(FullAdder_377_io_ci),
    .io_s(FullAdder_377_io_s),
    .io_co(FullAdder_377_io_co)
  );
  FullAdder FullAdder_378 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_378_io_a),
    .io_b(FullAdder_378_io_b),
    .io_ci(FullAdder_378_io_ci),
    .io_s(FullAdder_378_io_s),
    .io_co(FullAdder_378_io_co)
  );
  FullAdder FullAdder_379 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_379_io_a),
    .io_b(FullAdder_379_io_b),
    .io_ci(FullAdder_379_io_ci),
    .io_s(FullAdder_379_io_s),
    .io_co(FullAdder_379_io_co)
  );
  FullAdder FullAdder_380 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_380_io_a),
    .io_b(FullAdder_380_io_b),
    .io_ci(FullAdder_380_io_ci),
    .io_s(FullAdder_380_io_s),
    .io_co(FullAdder_380_io_co)
  );
  FullAdder FullAdder_381 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_381_io_a),
    .io_b(FullAdder_381_io_b),
    .io_ci(FullAdder_381_io_ci),
    .io_s(FullAdder_381_io_s),
    .io_co(FullAdder_381_io_co)
  );
  FullAdder FullAdder_382 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_382_io_a),
    .io_b(FullAdder_382_io_b),
    .io_ci(FullAdder_382_io_ci),
    .io_s(FullAdder_382_io_s),
    .io_co(FullAdder_382_io_co)
  );
  FullAdder FullAdder_383 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_383_io_a),
    .io_b(FullAdder_383_io_b),
    .io_ci(FullAdder_383_io_ci),
    .io_s(FullAdder_383_io_s),
    .io_co(FullAdder_383_io_co)
  );
  FullAdder FullAdder_384 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_384_io_a),
    .io_b(FullAdder_384_io_b),
    .io_ci(FullAdder_384_io_ci),
    .io_s(FullAdder_384_io_s),
    .io_co(FullAdder_384_io_co)
  );
  FullAdder FullAdder_385 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_385_io_a),
    .io_b(FullAdder_385_io_b),
    .io_ci(FullAdder_385_io_ci),
    .io_s(FullAdder_385_io_s),
    .io_co(FullAdder_385_io_co)
  );
  FullAdder FullAdder_386 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_386_io_a),
    .io_b(FullAdder_386_io_b),
    .io_ci(FullAdder_386_io_ci),
    .io_s(FullAdder_386_io_s),
    .io_co(FullAdder_386_io_co)
  );
  FullAdder FullAdder_387 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_387_io_a),
    .io_b(FullAdder_387_io_b),
    .io_ci(FullAdder_387_io_ci),
    .io_s(FullAdder_387_io_s),
    .io_co(FullAdder_387_io_co)
  );
  FullAdder FullAdder_388 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_388_io_a),
    .io_b(FullAdder_388_io_b),
    .io_ci(FullAdder_388_io_ci),
    .io_s(FullAdder_388_io_s),
    .io_co(FullAdder_388_io_co)
  );
  FullAdder FullAdder_389 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_389_io_a),
    .io_b(FullAdder_389_io_b),
    .io_ci(FullAdder_389_io_ci),
    .io_s(FullAdder_389_io_s),
    .io_co(FullAdder_389_io_co)
  );
  FullAdder FullAdder_390 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_390_io_a),
    .io_b(FullAdder_390_io_b),
    .io_ci(FullAdder_390_io_ci),
    .io_s(FullAdder_390_io_s),
    .io_co(FullAdder_390_io_co)
  );
  FullAdder FullAdder_391 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_391_io_a),
    .io_b(FullAdder_391_io_b),
    .io_ci(FullAdder_391_io_ci),
    .io_s(FullAdder_391_io_s),
    .io_co(FullAdder_391_io_co)
  );
  FullAdder FullAdder_392 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_392_io_a),
    .io_b(FullAdder_392_io_b),
    .io_ci(FullAdder_392_io_ci),
    .io_s(FullAdder_392_io_s),
    .io_co(FullAdder_392_io_co)
  );
  FullAdder FullAdder_393 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_393_io_a),
    .io_b(FullAdder_393_io_b),
    .io_ci(FullAdder_393_io_ci),
    .io_s(FullAdder_393_io_s),
    .io_co(FullAdder_393_io_co)
  );
  FullAdder FullAdder_394 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_394_io_a),
    .io_b(FullAdder_394_io_b),
    .io_ci(FullAdder_394_io_ci),
    .io_s(FullAdder_394_io_s),
    .io_co(FullAdder_394_io_co)
  );
  FullAdder FullAdder_395 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_395_io_a),
    .io_b(FullAdder_395_io_b),
    .io_ci(FullAdder_395_io_ci),
    .io_s(FullAdder_395_io_s),
    .io_co(FullAdder_395_io_co)
  );
  FullAdder FullAdder_396 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_396_io_a),
    .io_b(FullAdder_396_io_b),
    .io_ci(FullAdder_396_io_ci),
    .io_s(FullAdder_396_io_s),
    .io_co(FullAdder_396_io_co)
  );
  FullAdder FullAdder_397 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_397_io_a),
    .io_b(FullAdder_397_io_b),
    .io_ci(FullAdder_397_io_ci),
    .io_s(FullAdder_397_io_s),
    .io_co(FullAdder_397_io_co)
  );
  FullAdder FullAdder_398 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_398_io_a),
    .io_b(FullAdder_398_io_b),
    .io_ci(FullAdder_398_io_ci),
    .io_s(FullAdder_398_io_s),
    .io_co(FullAdder_398_io_co)
  );
  FullAdder FullAdder_399 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_399_io_a),
    .io_b(FullAdder_399_io_b),
    .io_ci(FullAdder_399_io_ci),
    .io_s(FullAdder_399_io_s),
    .io_co(FullAdder_399_io_co)
  );
  FullAdder FullAdder_400 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_400_io_a),
    .io_b(FullAdder_400_io_b),
    .io_ci(FullAdder_400_io_ci),
    .io_s(FullAdder_400_io_s),
    .io_co(FullAdder_400_io_co)
  );
  FullAdder FullAdder_401 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_401_io_a),
    .io_b(FullAdder_401_io_b),
    .io_ci(FullAdder_401_io_ci),
    .io_s(FullAdder_401_io_s),
    .io_co(FullAdder_401_io_co)
  );
  FullAdder FullAdder_402 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_402_io_a),
    .io_b(FullAdder_402_io_b),
    .io_ci(FullAdder_402_io_ci),
    .io_s(FullAdder_402_io_s),
    .io_co(FullAdder_402_io_co)
  );
  FullAdder FullAdder_403 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_403_io_a),
    .io_b(FullAdder_403_io_b),
    .io_ci(FullAdder_403_io_ci),
    .io_s(FullAdder_403_io_s),
    .io_co(FullAdder_403_io_co)
  );
  FullAdder FullAdder_404 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_404_io_a),
    .io_b(FullAdder_404_io_b),
    .io_ci(FullAdder_404_io_ci),
    .io_s(FullAdder_404_io_s),
    .io_co(FullAdder_404_io_co)
  );
  FullAdder FullAdder_405 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_405_io_a),
    .io_b(FullAdder_405_io_b),
    .io_ci(FullAdder_405_io_ci),
    .io_s(FullAdder_405_io_s),
    .io_co(FullAdder_405_io_co)
  );
  FullAdder FullAdder_406 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_406_io_a),
    .io_b(FullAdder_406_io_b),
    .io_ci(FullAdder_406_io_ci),
    .io_s(FullAdder_406_io_s),
    .io_co(FullAdder_406_io_co)
  );
  FullAdder FullAdder_407 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_407_io_a),
    .io_b(FullAdder_407_io_b),
    .io_ci(FullAdder_407_io_ci),
    .io_s(FullAdder_407_io_s),
    .io_co(FullAdder_407_io_co)
  );
  HalfAdder HalfAdder_13 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_13_io_a),
    .io_b(HalfAdder_13_io_b),
    .io_s(HalfAdder_13_io_s),
    .io_co(HalfAdder_13_io_co)
  );
  FullAdder FullAdder_408 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_408_io_a),
    .io_b(FullAdder_408_io_b),
    .io_ci(FullAdder_408_io_ci),
    .io_s(FullAdder_408_io_s),
    .io_co(FullAdder_408_io_co)
  );
  FullAdder FullAdder_409 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_409_io_a),
    .io_b(FullAdder_409_io_b),
    .io_ci(FullAdder_409_io_ci),
    .io_s(FullAdder_409_io_s),
    .io_co(FullAdder_409_io_co)
  );
  FullAdder FullAdder_410 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_410_io_a),
    .io_b(FullAdder_410_io_b),
    .io_ci(FullAdder_410_io_ci),
    .io_s(FullAdder_410_io_s),
    .io_co(FullAdder_410_io_co)
  );
  FullAdder FullAdder_411 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_411_io_a),
    .io_b(FullAdder_411_io_b),
    .io_ci(FullAdder_411_io_ci),
    .io_s(FullAdder_411_io_s),
    .io_co(FullAdder_411_io_co)
  );
  FullAdder FullAdder_412 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_412_io_a),
    .io_b(FullAdder_412_io_b),
    .io_ci(FullAdder_412_io_ci),
    .io_s(FullAdder_412_io_s),
    .io_co(FullAdder_412_io_co)
  );
  FullAdder FullAdder_413 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_413_io_a),
    .io_b(FullAdder_413_io_b),
    .io_ci(FullAdder_413_io_ci),
    .io_s(FullAdder_413_io_s),
    .io_co(FullAdder_413_io_co)
  );
  FullAdder FullAdder_414 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_414_io_a),
    .io_b(FullAdder_414_io_b),
    .io_ci(FullAdder_414_io_ci),
    .io_s(FullAdder_414_io_s),
    .io_co(FullAdder_414_io_co)
  );
  FullAdder FullAdder_415 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_415_io_a),
    .io_b(FullAdder_415_io_b),
    .io_ci(FullAdder_415_io_ci),
    .io_s(FullAdder_415_io_s),
    .io_co(FullAdder_415_io_co)
  );
  FullAdder FullAdder_416 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_416_io_a),
    .io_b(FullAdder_416_io_b),
    .io_ci(FullAdder_416_io_ci),
    .io_s(FullAdder_416_io_s),
    .io_co(FullAdder_416_io_co)
  );
  FullAdder FullAdder_417 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_417_io_a),
    .io_b(FullAdder_417_io_b),
    .io_ci(FullAdder_417_io_ci),
    .io_s(FullAdder_417_io_s),
    .io_co(FullAdder_417_io_co)
  );
  FullAdder FullAdder_418 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_418_io_a),
    .io_b(FullAdder_418_io_b),
    .io_ci(FullAdder_418_io_ci),
    .io_s(FullAdder_418_io_s),
    .io_co(FullAdder_418_io_co)
  );
  FullAdder FullAdder_419 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_419_io_a),
    .io_b(FullAdder_419_io_b),
    .io_ci(FullAdder_419_io_ci),
    .io_s(FullAdder_419_io_s),
    .io_co(FullAdder_419_io_co)
  );
  FullAdder FullAdder_420 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_420_io_a),
    .io_b(FullAdder_420_io_b),
    .io_ci(FullAdder_420_io_ci),
    .io_s(FullAdder_420_io_s),
    .io_co(FullAdder_420_io_co)
  );
  FullAdder FullAdder_421 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_421_io_a),
    .io_b(FullAdder_421_io_b),
    .io_ci(FullAdder_421_io_ci),
    .io_s(FullAdder_421_io_s),
    .io_co(FullAdder_421_io_co)
  );
  FullAdder FullAdder_422 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_422_io_a),
    .io_b(FullAdder_422_io_b),
    .io_ci(FullAdder_422_io_ci),
    .io_s(FullAdder_422_io_s),
    .io_co(FullAdder_422_io_co)
  );
  FullAdder FullAdder_423 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_423_io_a),
    .io_b(FullAdder_423_io_b),
    .io_ci(FullAdder_423_io_ci),
    .io_s(FullAdder_423_io_s),
    .io_co(FullAdder_423_io_co)
  );
  FullAdder FullAdder_424 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_424_io_a),
    .io_b(FullAdder_424_io_b),
    .io_ci(FullAdder_424_io_ci),
    .io_s(FullAdder_424_io_s),
    .io_co(FullAdder_424_io_co)
  );
  FullAdder FullAdder_425 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_425_io_a),
    .io_b(FullAdder_425_io_b),
    .io_ci(FullAdder_425_io_ci),
    .io_s(FullAdder_425_io_s),
    .io_co(FullAdder_425_io_co)
  );
  FullAdder FullAdder_426 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_426_io_a),
    .io_b(FullAdder_426_io_b),
    .io_ci(FullAdder_426_io_ci),
    .io_s(FullAdder_426_io_s),
    .io_co(FullAdder_426_io_co)
  );
  FullAdder FullAdder_427 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_427_io_a),
    .io_b(FullAdder_427_io_b),
    .io_ci(FullAdder_427_io_ci),
    .io_s(FullAdder_427_io_s),
    .io_co(FullAdder_427_io_co)
  );
  FullAdder FullAdder_428 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_428_io_a),
    .io_b(FullAdder_428_io_b),
    .io_ci(FullAdder_428_io_ci),
    .io_s(FullAdder_428_io_s),
    .io_co(FullAdder_428_io_co)
  );
  FullAdder FullAdder_429 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_429_io_a),
    .io_b(FullAdder_429_io_b),
    .io_ci(FullAdder_429_io_ci),
    .io_s(FullAdder_429_io_s),
    .io_co(FullAdder_429_io_co)
  );
  FullAdder FullAdder_430 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_430_io_a),
    .io_b(FullAdder_430_io_b),
    .io_ci(FullAdder_430_io_ci),
    .io_s(FullAdder_430_io_s),
    .io_co(FullAdder_430_io_co)
  );
  FullAdder FullAdder_431 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_431_io_a),
    .io_b(FullAdder_431_io_b),
    .io_ci(FullAdder_431_io_ci),
    .io_s(FullAdder_431_io_s),
    .io_co(FullAdder_431_io_co)
  );
  FullAdder FullAdder_432 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_432_io_a),
    .io_b(FullAdder_432_io_b),
    .io_ci(FullAdder_432_io_ci),
    .io_s(FullAdder_432_io_s),
    .io_co(FullAdder_432_io_co)
  );
  FullAdder FullAdder_433 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_433_io_a),
    .io_b(FullAdder_433_io_b),
    .io_ci(FullAdder_433_io_ci),
    .io_s(FullAdder_433_io_s),
    .io_co(FullAdder_433_io_co)
  );
  FullAdder FullAdder_434 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_434_io_a),
    .io_b(FullAdder_434_io_b),
    .io_ci(FullAdder_434_io_ci),
    .io_s(FullAdder_434_io_s),
    .io_co(FullAdder_434_io_co)
  );
  FullAdder FullAdder_435 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_435_io_a),
    .io_b(FullAdder_435_io_b),
    .io_ci(FullAdder_435_io_ci),
    .io_s(FullAdder_435_io_s),
    .io_co(FullAdder_435_io_co)
  );
  FullAdder FullAdder_436 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_436_io_a),
    .io_b(FullAdder_436_io_b),
    .io_ci(FullAdder_436_io_ci),
    .io_s(FullAdder_436_io_s),
    .io_co(FullAdder_436_io_co)
  );
  FullAdder FullAdder_437 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_437_io_a),
    .io_b(FullAdder_437_io_b),
    .io_ci(FullAdder_437_io_ci),
    .io_s(FullAdder_437_io_s),
    .io_co(FullAdder_437_io_co)
  );
  FullAdder FullAdder_438 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_438_io_a),
    .io_b(FullAdder_438_io_b),
    .io_ci(FullAdder_438_io_ci),
    .io_s(FullAdder_438_io_s),
    .io_co(FullAdder_438_io_co)
  );
  FullAdder FullAdder_439 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_439_io_a),
    .io_b(FullAdder_439_io_b),
    .io_ci(FullAdder_439_io_ci),
    .io_s(FullAdder_439_io_s),
    .io_co(FullAdder_439_io_co)
  );
  FullAdder FullAdder_440 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_440_io_a),
    .io_b(FullAdder_440_io_b),
    .io_ci(FullAdder_440_io_ci),
    .io_s(FullAdder_440_io_s),
    .io_co(FullAdder_440_io_co)
  );
  FullAdder FullAdder_441 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_441_io_a),
    .io_b(FullAdder_441_io_b),
    .io_ci(FullAdder_441_io_ci),
    .io_s(FullAdder_441_io_s),
    .io_co(FullAdder_441_io_co)
  );
  FullAdder FullAdder_442 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_442_io_a),
    .io_b(FullAdder_442_io_b),
    .io_ci(FullAdder_442_io_ci),
    .io_s(FullAdder_442_io_s),
    .io_co(FullAdder_442_io_co)
  );
  FullAdder FullAdder_443 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_443_io_a),
    .io_b(FullAdder_443_io_b),
    .io_ci(FullAdder_443_io_ci),
    .io_s(FullAdder_443_io_s),
    .io_co(FullAdder_443_io_co)
  );
  FullAdder FullAdder_444 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_444_io_a),
    .io_b(FullAdder_444_io_b),
    .io_ci(FullAdder_444_io_ci),
    .io_s(FullAdder_444_io_s),
    .io_co(FullAdder_444_io_co)
  );
  FullAdder FullAdder_445 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_445_io_a),
    .io_b(FullAdder_445_io_b),
    .io_ci(FullAdder_445_io_ci),
    .io_s(FullAdder_445_io_s),
    .io_co(FullAdder_445_io_co)
  );
  FullAdder FullAdder_446 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_446_io_a),
    .io_b(FullAdder_446_io_b),
    .io_ci(FullAdder_446_io_ci),
    .io_s(FullAdder_446_io_s),
    .io_co(FullAdder_446_io_co)
  );
  FullAdder FullAdder_447 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_447_io_a),
    .io_b(FullAdder_447_io_b),
    .io_ci(FullAdder_447_io_ci),
    .io_s(FullAdder_447_io_s),
    .io_co(FullAdder_447_io_co)
  );
  FullAdder FullAdder_448 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_448_io_a),
    .io_b(FullAdder_448_io_b),
    .io_ci(FullAdder_448_io_ci),
    .io_s(FullAdder_448_io_s),
    .io_co(FullAdder_448_io_co)
  );
  FullAdder FullAdder_449 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_449_io_a),
    .io_b(FullAdder_449_io_b),
    .io_ci(FullAdder_449_io_ci),
    .io_s(FullAdder_449_io_s),
    .io_co(FullAdder_449_io_co)
  );
  FullAdder FullAdder_450 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_450_io_a),
    .io_b(FullAdder_450_io_b),
    .io_ci(FullAdder_450_io_ci),
    .io_s(FullAdder_450_io_s),
    .io_co(FullAdder_450_io_co)
  );
  FullAdder FullAdder_451 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_451_io_a),
    .io_b(FullAdder_451_io_b),
    .io_ci(FullAdder_451_io_ci),
    .io_s(FullAdder_451_io_s),
    .io_co(FullAdder_451_io_co)
  );
  FullAdder FullAdder_452 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_452_io_a),
    .io_b(FullAdder_452_io_b),
    .io_ci(FullAdder_452_io_ci),
    .io_s(FullAdder_452_io_s),
    .io_co(FullAdder_452_io_co)
  );
  FullAdder FullAdder_453 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_453_io_a),
    .io_b(FullAdder_453_io_b),
    .io_ci(FullAdder_453_io_ci),
    .io_s(FullAdder_453_io_s),
    .io_co(FullAdder_453_io_co)
  );
  FullAdder FullAdder_454 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_454_io_a),
    .io_b(FullAdder_454_io_b),
    .io_ci(FullAdder_454_io_ci),
    .io_s(FullAdder_454_io_s),
    .io_co(FullAdder_454_io_co)
  );
  FullAdder FullAdder_455 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_455_io_a),
    .io_b(FullAdder_455_io_b),
    .io_ci(FullAdder_455_io_ci),
    .io_s(FullAdder_455_io_s),
    .io_co(FullAdder_455_io_co)
  );
  FullAdder FullAdder_456 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_456_io_a),
    .io_b(FullAdder_456_io_b),
    .io_ci(FullAdder_456_io_ci),
    .io_s(FullAdder_456_io_s),
    .io_co(FullAdder_456_io_co)
  );
  FullAdder FullAdder_457 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_457_io_a),
    .io_b(FullAdder_457_io_b),
    .io_ci(FullAdder_457_io_ci),
    .io_s(FullAdder_457_io_s),
    .io_co(FullAdder_457_io_co)
  );
  FullAdder FullAdder_458 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_458_io_a),
    .io_b(FullAdder_458_io_b),
    .io_ci(FullAdder_458_io_ci),
    .io_s(FullAdder_458_io_s),
    .io_co(FullAdder_458_io_co)
  );
  HalfAdder HalfAdder_14 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_14_io_a),
    .io_b(HalfAdder_14_io_b),
    .io_s(HalfAdder_14_io_s),
    .io_co(HalfAdder_14_io_co)
  );
  FullAdder FullAdder_459 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_459_io_a),
    .io_b(FullAdder_459_io_b),
    .io_ci(FullAdder_459_io_ci),
    .io_s(FullAdder_459_io_s),
    .io_co(FullAdder_459_io_co)
  );
  FullAdder FullAdder_460 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_460_io_a),
    .io_b(FullAdder_460_io_b),
    .io_ci(FullAdder_460_io_ci),
    .io_s(FullAdder_460_io_s),
    .io_co(FullAdder_460_io_co)
  );
  FullAdder FullAdder_461 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_461_io_a),
    .io_b(FullAdder_461_io_b),
    .io_ci(FullAdder_461_io_ci),
    .io_s(FullAdder_461_io_s),
    .io_co(FullAdder_461_io_co)
  );
  FullAdder FullAdder_462 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_462_io_a),
    .io_b(FullAdder_462_io_b),
    .io_ci(FullAdder_462_io_ci),
    .io_s(FullAdder_462_io_s),
    .io_co(FullAdder_462_io_co)
  );
  FullAdder FullAdder_463 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_463_io_a),
    .io_b(FullAdder_463_io_b),
    .io_ci(FullAdder_463_io_ci),
    .io_s(FullAdder_463_io_s),
    .io_co(FullAdder_463_io_co)
  );
  FullAdder FullAdder_464 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_464_io_a),
    .io_b(FullAdder_464_io_b),
    .io_ci(FullAdder_464_io_ci),
    .io_s(FullAdder_464_io_s),
    .io_co(FullAdder_464_io_co)
  );
  FullAdder FullAdder_465 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_465_io_a),
    .io_b(FullAdder_465_io_b),
    .io_ci(FullAdder_465_io_ci),
    .io_s(FullAdder_465_io_s),
    .io_co(FullAdder_465_io_co)
  );
  FullAdder FullAdder_466 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_466_io_a),
    .io_b(FullAdder_466_io_b),
    .io_ci(FullAdder_466_io_ci),
    .io_s(FullAdder_466_io_s),
    .io_co(FullAdder_466_io_co)
  );
  FullAdder FullAdder_467 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_467_io_a),
    .io_b(FullAdder_467_io_b),
    .io_ci(FullAdder_467_io_ci),
    .io_s(FullAdder_467_io_s),
    .io_co(FullAdder_467_io_co)
  );
  FullAdder FullAdder_468 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_468_io_a),
    .io_b(FullAdder_468_io_b),
    .io_ci(FullAdder_468_io_ci),
    .io_s(FullAdder_468_io_s),
    .io_co(FullAdder_468_io_co)
  );
  FullAdder FullAdder_469 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_469_io_a),
    .io_b(FullAdder_469_io_b),
    .io_ci(FullAdder_469_io_ci),
    .io_s(FullAdder_469_io_s),
    .io_co(FullAdder_469_io_co)
  );
  FullAdder FullAdder_470 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_470_io_a),
    .io_b(FullAdder_470_io_b),
    .io_ci(FullAdder_470_io_ci),
    .io_s(FullAdder_470_io_s),
    .io_co(FullAdder_470_io_co)
  );
  FullAdder FullAdder_471 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_471_io_a),
    .io_b(FullAdder_471_io_b),
    .io_ci(FullAdder_471_io_ci),
    .io_s(FullAdder_471_io_s),
    .io_co(FullAdder_471_io_co)
  );
  FullAdder FullAdder_472 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_472_io_a),
    .io_b(FullAdder_472_io_b),
    .io_ci(FullAdder_472_io_ci),
    .io_s(FullAdder_472_io_s),
    .io_co(FullAdder_472_io_co)
  );
  FullAdder FullAdder_473 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_473_io_a),
    .io_b(FullAdder_473_io_b),
    .io_ci(FullAdder_473_io_ci),
    .io_s(FullAdder_473_io_s),
    .io_co(FullAdder_473_io_co)
  );
  FullAdder FullAdder_474 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_474_io_a),
    .io_b(FullAdder_474_io_b),
    .io_ci(FullAdder_474_io_ci),
    .io_s(FullAdder_474_io_s),
    .io_co(FullAdder_474_io_co)
  );
  FullAdder FullAdder_475 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_475_io_a),
    .io_b(FullAdder_475_io_b),
    .io_ci(FullAdder_475_io_ci),
    .io_s(FullAdder_475_io_s),
    .io_co(FullAdder_475_io_co)
  );
  FullAdder FullAdder_476 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_476_io_a),
    .io_b(FullAdder_476_io_b),
    .io_ci(FullAdder_476_io_ci),
    .io_s(FullAdder_476_io_s),
    .io_co(FullAdder_476_io_co)
  );
  FullAdder FullAdder_477 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_477_io_a),
    .io_b(FullAdder_477_io_b),
    .io_ci(FullAdder_477_io_ci),
    .io_s(FullAdder_477_io_s),
    .io_co(FullAdder_477_io_co)
  );
  FullAdder FullAdder_478 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_478_io_a),
    .io_b(FullAdder_478_io_b),
    .io_ci(FullAdder_478_io_ci),
    .io_s(FullAdder_478_io_s),
    .io_co(FullAdder_478_io_co)
  );
  FullAdder FullAdder_479 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_479_io_a),
    .io_b(FullAdder_479_io_b),
    .io_ci(FullAdder_479_io_ci),
    .io_s(FullAdder_479_io_s),
    .io_co(FullAdder_479_io_co)
  );
  FullAdder FullAdder_480 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_480_io_a),
    .io_b(FullAdder_480_io_b),
    .io_ci(FullAdder_480_io_ci),
    .io_s(FullAdder_480_io_s),
    .io_co(FullAdder_480_io_co)
  );
  FullAdder FullAdder_481 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_481_io_a),
    .io_b(FullAdder_481_io_b),
    .io_ci(FullAdder_481_io_ci),
    .io_s(FullAdder_481_io_s),
    .io_co(FullAdder_481_io_co)
  );
  FullAdder FullAdder_482 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_482_io_a),
    .io_b(FullAdder_482_io_b),
    .io_ci(FullAdder_482_io_ci),
    .io_s(FullAdder_482_io_s),
    .io_co(FullAdder_482_io_co)
  );
  FullAdder FullAdder_483 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_483_io_a),
    .io_b(FullAdder_483_io_b),
    .io_ci(FullAdder_483_io_ci),
    .io_s(FullAdder_483_io_s),
    .io_co(FullAdder_483_io_co)
  );
  FullAdder FullAdder_484 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_484_io_a),
    .io_b(FullAdder_484_io_b),
    .io_ci(FullAdder_484_io_ci),
    .io_s(FullAdder_484_io_s),
    .io_co(FullAdder_484_io_co)
  );
  FullAdder FullAdder_485 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_485_io_a),
    .io_b(FullAdder_485_io_b),
    .io_ci(FullAdder_485_io_ci),
    .io_s(FullAdder_485_io_s),
    .io_co(FullAdder_485_io_co)
  );
  FullAdder FullAdder_486 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_486_io_a),
    .io_b(FullAdder_486_io_b),
    .io_ci(FullAdder_486_io_ci),
    .io_s(FullAdder_486_io_s),
    .io_co(FullAdder_486_io_co)
  );
  FullAdder FullAdder_487 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_487_io_a),
    .io_b(FullAdder_487_io_b),
    .io_ci(FullAdder_487_io_ci),
    .io_s(FullAdder_487_io_s),
    .io_co(FullAdder_487_io_co)
  );
  FullAdder FullAdder_488 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_488_io_a),
    .io_b(FullAdder_488_io_b),
    .io_ci(FullAdder_488_io_ci),
    .io_s(FullAdder_488_io_s),
    .io_co(FullAdder_488_io_co)
  );
  FullAdder FullAdder_489 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_489_io_a),
    .io_b(FullAdder_489_io_b),
    .io_ci(FullAdder_489_io_ci),
    .io_s(FullAdder_489_io_s),
    .io_co(FullAdder_489_io_co)
  );
  FullAdder FullAdder_490 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_490_io_a),
    .io_b(FullAdder_490_io_b),
    .io_ci(FullAdder_490_io_ci),
    .io_s(FullAdder_490_io_s),
    .io_co(FullAdder_490_io_co)
  );
  FullAdder FullAdder_491 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_491_io_a),
    .io_b(FullAdder_491_io_b),
    .io_ci(FullAdder_491_io_ci),
    .io_s(FullAdder_491_io_s),
    .io_co(FullAdder_491_io_co)
  );
  FullAdder FullAdder_492 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_492_io_a),
    .io_b(FullAdder_492_io_b),
    .io_ci(FullAdder_492_io_ci),
    .io_s(FullAdder_492_io_s),
    .io_co(FullAdder_492_io_co)
  );
  FullAdder FullAdder_493 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_493_io_a),
    .io_b(FullAdder_493_io_b),
    .io_ci(FullAdder_493_io_ci),
    .io_s(FullAdder_493_io_s),
    .io_co(FullAdder_493_io_co)
  );
  FullAdder FullAdder_494 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_494_io_a),
    .io_b(FullAdder_494_io_b),
    .io_ci(FullAdder_494_io_ci),
    .io_s(FullAdder_494_io_s),
    .io_co(FullAdder_494_io_co)
  );
  FullAdder FullAdder_495 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_495_io_a),
    .io_b(FullAdder_495_io_b),
    .io_ci(FullAdder_495_io_ci),
    .io_s(FullAdder_495_io_s),
    .io_co(FullAdder_495_io_co)
  );
  FullAdder FullAdder_496 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_496_io_a),
    .io_b(FullAdder_496_io_b),
    .io_ci(FullAdder_496_io_ci),
    .io_s(FullAdder_496_io_s),
    .io_co(FullAdder_496_io_co)
  );
  FullAdder FullAdder_497 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_497_io_a),
    .io_b(FullAdder_497_io_b),
    .io_ci(FullAdder_497_io_ci),
    .io_s(FullAdder_497_io_s),
    .io_co(FullAdder_497_io_co)
  );
  FullAdder FullAdder_498 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_498_io_a),
    .io_b(FullAdder_498_io_b),
    .io_ci(FullAdder_498_io_ci),
    .io_s(FullAdder_498_io_s),
    .io_co(FullAdder_498_io_co)
  );
  FullAdder FullAdder_499 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_499_io_a),
    .io_b(FullAdder_499_io_b),
    .io_ci(FullAdder_499_io_ci),
    .io_s(FullAdder_499_io_s),
    .io_co(FullAdder_499_io_co)
  );
  FullAdder FullAdder_500 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_500_io_a),
    .io_b(FullAdder_500_io_b),
    .io_ci(FullAdder_500_io_ci),
    .io_s(FullAdder_500_io_s),
    .io_co(FullAdder_500_io_co)
  );
  FullAdder FullAdder_501 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_501_io_a),
    .io_b(FullAdder_501_io_b),
    .io_ci(FullAdder_501_io_ci),
    .io_s(FullAdder_501_io_s),
    .io_co(FullAdder_501_io_co)
  );
  FullAdder FullAdder_502 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_502_io_a),
    .io_b(FullAdder_502_io_b),
    .io_ci(FullAdder_502_io_ci),
    .io_s(FullAdder_502_io_s),
    .io_co(FullAdder_502_io_co)
  );
  FullAdder FullAdder_503 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_503_io_a),
    .io_b(FullAdder_503_io_b),
    .io_ci(FullAdder_503_io_ci),
    .io_s(FullAdder_503_io_s),
    .io_co(FullAdder_503_io_co)
  );
  FullAdder FullAdder_504 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_504_io_a),
    .io_b(FullAdder_504_io_b),
    .io_ci(FullAdder_504_io_ci),
    .io_s(FullAdder_504_io_s),
    .io_co(FullAdder_504_io_co)
  );
  FullAdder FullAdder_505 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_505_io_a),
    .io_b(FullAdder_505_io_b),
    .io_ci(FullAdder_505_io_ci),
    .io_s(FullAdder_505_io_s),
    .io_co(FullAdder_505_io_co)
  );
  FullAdder FullAdder_506 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_506_io_a),
    .io_b(FullAdder_506_io_b),
    .io_ci(FullAdder_506_io_ci),
    .io_s(FullAdder_506_io_s),
    .io_co(FullAdder_506_io_co)
  );
  FullAdder FullAdder_507 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_507_io_a),
    .io_b(FullAdder_507_io_b),
    .io_ci(FullAdder_507_io_ci),
    .io_s(FullAdder_507_io_s),
    .io_co(FullAdder_507_io_co)
  );
  FullAdder FullAdder_508 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_508_io_a),
    .io_b(FullAdder_508_io_b),
    .io_ci(FullAdder_508_io_ci),
    .io_s(FullAdder_508_io_s),
    .io_co(FullAdder_508_io_co)
  );
  FullAdder FullAdder_509 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_509_io_a),
    .io_b(FullAdder_509_io_b),
    .io_ci(FullAdder_509_io_ci),
    .io_s(FullAdder_509_io_s),
    .io_co(FullAdder_509_io_co)
  );
  FullAdder FullAdder_510 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_510_io_a),
    .io_b(FullAdder_510_io_b),
    .io_ci(FullAdder_510_io_ci),
    .io_s(FullAdder_510_io_s),
    .io_co(FullAdder_510_io_co)
  );
  FullAdder FullAdder_511 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_511_io_a),
    .io_b(FullAdder_511_io_b),
    .io_ci(FullAdder_511_io_ci),
    .io_s(FullAdder_511_io_s),
    .io_co(FullAdder_511_io_co)
  );
  FullAdder FullAdder_512 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_512_io_a),
    .io_b(FullAdder_512_io_b),
    .io_ci(FullAdder_512_io_ci),
    .io_s(FullAdder_512_io_s),
    .io_co(FullAdder_512_io_co)
  );
  HalfAdder HalfAdder_15 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_15_io_a),
    .io_b(HalfAdder_15_io_b),
    .io_s(HalfAdder_15_io_s),
    .io_co(HalfAdder_15_io_co)
  );
  FullAdder FullAdder_513 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_513_io_a),
    .io_b(FullAdder_513_io_b),
    .io_ci(FullAdder_513_io_ci),
    .io_s(FullAdder_513_io_s),
    .io_co(FullAdder_513_io_co)
  );
  FullAdder FullAdder_514 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_514_io_a),
    .io_b(FullAdder_514_io_b),
    .io_ci(FullAdder_514_io_ci),
    .io_s(FullAdder_514_io_s),
    .io_co(FullAdder_514_io_co)
  );
  FullAdder FullAdder_515 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_515_io_a),
    .io_b(FullAdder_515_io_b),
    .io_ci(FullAdder_515_io_ci),
    .io_s(FullAdder_515_io_s),
    .io_co(FullAdder_515_io_co)
  );
  FullAdder FullAdder_516 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_516_io_a),
    .io_b(FullAdder_516_io_b),
    .io_ci(FullAdder_516_io_ci),
    .io_s(FullAdder_516_io_s),
    .io_co(FullAdder_516_io_co)
  );
  FullAdder FullAdder_517 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_517_io_a),
    .io_b(FullAdder_517_io_b),
    .io_ci(FullAdder_517_io_ci),
    .io_s(FullAdder_517_io_s),
    .io_co(FullAdder_517_io_co)
  );
  FullAdder FullAdder_518 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_518_io_a),
    .io_b(FullAdder_518_io_b),
    .io_ci(FullAdder_518_io_ci),
    .io_s(FullAdder_518_io_s),
    .io_co(FullAdder_518_io_co)
  );
  FullAdder FullAdder_519 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_519_io_a),
    .io_b(FullAdder_519_io_b),
    .io_ci(FullAdder_519_io_ci),
    .io_s(FullAdder_519_io_s),
    .io_co(FullAdder_519_io_co)
  );
  FullAdder FullAdder_520 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_520_io_a),
    .io_b(FullAdder_520_io_b),
    .io_ci(FullAdder_520_io_ci),
    .io_s(FullAdder_520_io_s),
    .io_co(FullAdder_520_io_co)
  );
  FullAdder FullAdder_521 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_521_io_a),
    .io_b(FullAdder_521_io_b),
    .io_ci(FullAdder_521_io_ci),
    .io_s(FullAdder_521_io_s),
    .io_co(FullAdder_521_io_co)
  );
  FullAdder FullAdder_522 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_522_io_a),
    .io_b(FullAdder_522_io_b),
    .io_ci(FullAdder_522_io_ci),
    .io_s(FullAdder_522_io_s),
    .io_co(FullAdder_522_io_co)
  );
  FullAdder FullAdder_523 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_523_io_a),
    .io_b(FullAdder_523_io_b),
    .io_ci(FullAdder_523_io_ci),
    .io_s(FullAdder_523_io_s),
    .io_co(FullAdder_523_io_co)
  );
  FullAdder FullAdder_524 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_524_io_a),
    .io_b(FullAdder_524_io_b),
    .io_ci(FullAdder_524_io_ci),
    .io_s(FullAdder_524_io_s),
    .io_co(FullAdder_524_io_co)
  );
  FullAdder FullAdder_525 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_525_io_a),
    .io_b(FullAdder_525_io_b),
    .io_ci(FullAdder_525_io_ci),
    .io_s(FullAdder_525_io_s),
    .io_co(FullAdder_525_io_co)
  );
  FullAdder FullAdder_526 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_526_io_a),
    .io_b(FullAdder_526_io_b),
    .io_ci(FullAdder_526_io_ci),
    .io_s(FullAdder_526_io_s),
    .io_co(FullAdder_526_io_co)
  );
  FullAdder FullAdder_527 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_527_io_a),
    .io_b(FullAdder_527_io_b),
    .io_ci(FullAdder_527_io_ci),
    .io_s(FullAdder_527_io_s),
    .io_co(FullAdder_527_io_co)
  );
  FullAdder FullAdder_528 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_528_io_a),
    .io_b(FullAdder_528_io_b),
    .io_ci(FullAdder_528_io_ci),
    .io_s(FullAdder_528_io_s),
    .io_co(FullAdder_528_io_co)
  );
  FullAdder FullAdder_529 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_529_io_a),
    .io_b(FullAdder_529_io_b),
    .io_ci(FullAdder_529_io_ci),
    .io_s(FullAdder_529_io_s),
    .io_co(FullAdder_529_io_co)
  );
  FullAdder FullAdder_530 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_530_io_a),
    .io_b(FullAdder_530_io_b),
    .io_ci(FullAdder_530_io_ci),
    .io_s(FullAdder_530_io_s),
    .io_co(FullAdder_530_io_co)
  );
  FullAdder FullAdder_531 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_531_io_a),
    .io_b(FullAdder_531_io_b),
    .io_ci(FullAdder_531_io_ci),
    .io_s(FullAdder_531_io_s),
    .io_co(FullAdder_531_io_co)
  );
  FullAdder FullAdder_532 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_532_io_a),
    .io_b(FullAdder_532_io_b),
    .io_ci(FullAdder_532_io_ci),
    .io_s(FullAdder_532_io_s),
    .io_co(FullAdder_532_io_co)
  );
  FullAdder FullAdder_533 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_533_io_a),
    .io_b(FullAdder_533_io_b),
    .io_ci(FullAdder_533_io_ci),
    .io_s(FullAdder_533_io_s),
    .io_co(FullAdder_533_io_co)
  );
  FullAdder FullAdder_534 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_534_io_a),
    .io_b(FullAdder_534_io_b),
    .io_ci(FullAdder_534_io_ci),
    .io_s(FullAdder_534_io_s),
    .io_co(FullAdder_534_io_co)
  );
  FullAdder FullAdder_535 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_535_io_a),
    .io_b(FullAdder_535_io_b),
    .io_ci(FullAdder_535_io_ci),
    .io_s(FullAdder_535_io_s),
    .io_co(FullAdder_535_io_co)
  );
  FullAdder FullAdder_536 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_536_io_a),
    .io_b(FullAdder_536_io_b),
    .io_ci(FullAdder_536_io_ci),
    .io_s(FullAdder_536_io_s),
    .io_co(FullAdder_536_io_co)
  );
  FullAdder FullAdder_537 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_537_io_a),
    .io_b(FullAdder_537_io_b),
    .io_ci(FullAdder_537_io_ci),
    .io_s(FullAdder_537_io_s),
    .io_co(FullAdder_537_io_co)
  );
  FullAdder FullAdder_538 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_538_io_a),
    .io_b(FullAdder_538_io_b),
    .io_ci(FullAdder_538_io_ci),
    .io_s(FullAdder_538_io_s),
    .io_co(FullAdder_538_io_co)
  );
  FullAdder FullAdder_539 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_539_io_a),
    .io_b(FullAdder_539_io_b),
    .io_ci(FullAdder_539_io_ci),
    .io_s(FullAdder_539_io_s),
    .io_co(FullAdder_539_io_co)
  );
  FullAdder FullAdder_540 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_540_io_a),
    .io_b(FullAdder_540_io_b),
    .io_ci(FullAdder_540_io_ci),
    .io_s(FullAdder_540_io_s),
    .io_co(FullAdder_540_io_co)
  );
  FullAdder FullAdder_541 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_541_io_a),
    .io_b(FullAdder_541_io_b),
    .io_ci(FullAdder_541_io_ci),
    .io_s(FullAdder_541_io_s),
    .io_co(FullAdder_541_io_co)
  );
  FullAdder FullAdder_542 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_542_io_a),
    .io_b(FullAdder_542_io_b),
    .io_ci(FullAdder_542_io_ci),
    .io_s(FullAdder_542_io_s),
    .io_co(FullAdder_542_io_co)
  );
  FullAdder FullAdder_543 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_543_io_a),
    .io_b(FullAdder_543_io_b),
    .io_ci(FullAdder_543_io_ci),
    .io_s(FullAdder_543_io_s),
    .io_co(FullAdder_543_io_co)
  );
  FullAdder FullAdder_544 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_544_io_a),
    .io_b(FullAdder_544_io_b),
    .io_ci(FullAdder_544_io_ci),
    .io_s(FullAdder_544_io_s),
    .io_co(FullAdder_544_io_co)
  );
  FullAdder FullAdder_545 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_545_io_a),
    .io_b(FullAdder_545_io_b),
    .io_ci(FullAdder_545_io_ci),
    .io_s(FullAdder_545_io_s),
    .io_co(FullAdder_545_io_co)
  );
  FullAdder FullAdder_546 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_546_io_a),
    .io_b(FullAdder_546_io_b),
    .io_ci(FullAdder_546_io_ci),
    .io_s(FullAdder_546_io_s),
    .io_co(FullAdder_546_io_co)
  );
  FullAdder FullAdder_547 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_547_io_a),
    .io_b(FullAdder_547_io_b),
    .io_ci(FullAdder_547_io_ci),
    .io_s(FullAdder_547_io_s),
    .io_co(FullAdder_547_io_co)
  );
  FullAdder FullAdder_548 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_548_io_a),
    .io_b(FullAdder_548_io_b),
    .io_ci(FullAdder_548_io_ci),
    .io_s(FullAdder_548_io_s),
    .io_co(FullAdder_548_io_co)
  );
  FullAdder FullAdder_549 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_549_io_a),
    .io_b(FullAdder_549_io_b),
    .io_ci(FullAdder_549_io_ci),
    .io_s(FullAdder_549_io_s),
    .io_co(FullAdder_549_io_co)
  );
  FullAdder FullAdder_550 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_550_io_a),
    .io_b(FullAdder_550_io_b),
    .io_ci(FullAdder_550_io_ci),
    .io_s(FullAdder_550_io_s),
    .io_co(FullAdder_550_io_co)
  );
  FullAdder FullAdder_551 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_551_io_a),
    .io_b(FullAdder_551_io_b),
    .io_ci(FullAdder_551_io_ci),
    .io_s(FullAdder_551_io_s),
    .io_co(FullAdder_551_io_co)
  );
  FullAdder FullAdder_552 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_552_io_a),
    .io_b(FullAdder_552_io_b),
    .io_ci(FullAdder_552_io_ci),
    .io_s(FullAdder_552_io_s),
    .io_co(FullAdder_552_io_co)
  );
  FullAdder FullAdder_553 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_553_io_a),
    .io_b(FullAdder_553_io_b),
    .io_ci(FullAdder_553_io_ci),
    .io_s(FullAdder_553_io_s),
    .io_co(FullAdder_553_io_co)
  );
  FullAdder FullAdder_554 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_554_io_a),
    .io_b(FullAdder_554_io_b),
    .io_ci(FullAdder_554_io_ci),
    .io_s(FullAdder_554_io_s),
    .io_co(FullAdder_554_io_co)
  );
  FullAdder FullAdder_555 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_555_io_a),
    .io_b(FullAdder_555_io_b),
    .io_ci(FullAdder_555_io_ci),
    .io_s(FullAdder_555_io_s),
    .io_co(FullAdder_555_io_co)
  );
  FullAdder FullAdder_556 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_556_io_a),
    .io_b(FullAdder_556_io_b),
    .io_ci(FullAdder_556_io_ci),
    .io_s(FullAdder_556_io_s),
    .io_co(FullAdder_556_io_co)
  );
  FullAdder FullAdder_557 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_557_io_a),
    .io_b(FullAdder_557_io_b),
    .io_ci(FullAdder_557_io_ci),
    .io_s(FullAdder_557_io_s),
    .io_co(FullAdder_557_io_co)
  );
  FullAdder FullAdder_558 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_558_io_a),
    .io_b(FullAdder_558_io_b),
    .io_ci(FullAdder_558_io_ci),
    .io_s(FullAdder_558_io_s),
    .io_co(FullAdder_558_io_co)
  );
  FullAdder FullAdder_559 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_559_io_a),
    .io_b(FullAdder_559_io_b),
    .io_ci(FullAdder_559_io_ci),
    .io_s(FullAdder_559_io_s),
    .io_co(FullAdder_559_io_co)
  );
  FullAdder FullAdder_560 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_560_io_a),
    .io_b(FullAdder_560_io_b),
    .io_ci(FullAdder_560_io_ci),
    .io_s(FullAdder_560_io_s),
    .io_co(FullAdder_560_io_co)
  );
  FullAdder FullAdder_561 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_561_io_a),
    .io_b(FullAdder_561_io_b),
    .io_ci(FullAdder_561_io_ci),
    .io_s(FullAdder_561_io_s),
    .io_co(FullAdder_561_io_co)
  );
  FullAdder FullAdder_562 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_562_io_a),
    .io_b(FullAdder_562_io_b),
    .io_ci(FullAdder_562_io_ci),
    .io_s(FullAdder_562_io_s),
    .io_co(FullAdder_562_io_co)
  );
  FullAdder FullAdder_563 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_563_io_a),
    .io_b(FullAdder_563_io_b),
    .io_ci(FullAdder_563_io_ci),
    .io_s(FullAdder_563_io_s),
    .io_co(FullAdder_563_io_co)
  );
  FullAdder FullAdder_564 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_564_io_a),
    .io_b(FullAdder_564_io_b),
    .io_ci(FullAdder_564_io_ci),
    .io_s(FullAdder_564_io_s),
    .io_co(FullAdder_564_io_co)
  );
  FullAdder FullAdder_565 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_565_io_a),
    .io_b(FullAdder_565_io_b),
    .io_ci(FullAdder_565_io_ci),
    .io_s(FullAdder_565_io_s),
    .io_co(FullAdder_565_io_co)
  );
  FullAdder FullAdder_566 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_566_io_a),
    .io_b(FullAdder_566_io_b),
    .io_ci(FullAdder_566_io_ci),
    .io_s(FullAdder_566_io_s),
    .io_co(FullAdder_566_io_co)
  );
  FullAdder FullAdder_567 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_567_io_a),
    .io_b(FullAdder_567_io_b),
    .io_ci(FullAdder_567_io_ci),
    .io_s(FullAdder_567_io_s),
    .io_co(FullAdder_567_io_co)
  );
  FullAdder FullAdder_568 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_568_io_a),
    .io_b(FullAdder_568_io_b),
    .io_ci(FullAdder_568_io_ci),
    .io_s(FullAdder_568_io_s),
    .io_co(FullAdder_568_io_co)
  );
  FullAdder FullAdder_569 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_569_io_a),
    .io_b(FullAdder_569_io_b),
    .io_ci(FullAdder_569_io_ci),
    .io_s(FullAdder_569_io_s),
    .io_co(FullAdder_569_io_co)
  );
  HalfAdder HalfAdder_16 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_16_io_a),
    .io_b(HalfAdder_16_io_b),
    .io_s(HalfAdder_16_io_s),
    .io_co(HalfAdder_16_io_co)
  );
  FullAdder FullAdder_570 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_570_io_a),
    .io_b(FullAdder_570_io_b),
    .io_ci(FullAdder_570_io_ci),
    .io_s(FullAdder_570_io_s),
    .io_co(FullAdder_570_io_co)
  );
  FullAdder FullAdder_571 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_571_io_a),
    .io_b(FullAdder_571_io_b),
    .io_ci(FullAdder_571_io_ci),
    .io_s(FullAdder_571_io_s),
    .io_co(FullAdder_571_io_co)
  );
  FullAdder FullAdder_572 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_572_io_a),
    .io_b(FullAdder_572_io_b),
    .io_ci(FullAdder_572_io_ci),
    .io_s(FullAdder_572_io_s),
    .io_co(FullAdder_572_io_co)
  );
  FullAdder FullAdder_573 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_573_io_a),
    .io_b(FullAdder_573_io_b),
    .io_ci(FullAdder_573_io_ci),
    .io_s(FullAdder_573_io_s),
    .io_co(FullAdder_573_io_co)
  );
  FullAdder FullAdder_574 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_574_io_a),
    .io_b(FullAdder_574_io_b),
    .io_ci(FullAdder_574_io_ci),
    .io_s(FullAdder_574_io_s),
    .io_co(FullAdder_574_io_co)
  );
  FullAdder FullAdder_575 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_575_io_a),
    .io_b(FullAdder_575_io_b),
    .io_ci(FullAdder_575_io_ci),
    .io_s(FullAdder_575_io_s),
    .io_co(FullAdder_575_io_co)
  );
  FullAdder FullAdder_576 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_576_io_a),
    .io_b(FullAdder_576_io_b),
    .io_ci(FullAdder_576_io_ci),
    .io_s(FullAdder_576_io_s),
    .io_co(FullAdder_576_io_co)
  );
  FullAdder FullAdder_577 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_577_io_a),
    .io_b(FullAdder_577_io_b),
    .io_ci(FullAdder_577_io_ci),
    .io_s(FullAdder_577_io_s),
    .io_co(FullAdder_577_io_co)
  );
  FullAdder FullAdder_578 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_578_io_a),
    .io_b(FullAdder_578_io_b),
    .io_ci(FullAdder_578_io_ci),
    .io_s(FullAdder_578_io_s),
    .io_co(FullAdder_578_io_co)
  );
  FullAdder FullAdder_579 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_579_io_a),
    .io_b(FullAdder_579_io_b),
    .io_ci(FullAdder_579_io_ci),
    .io_s(FullAdder_579_io_s),
    .io_co(FullAdder_579_io_co)
  );
  FullAdder FullAdder_580 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_580_io_a),
    .io_b(FullAdder_580_io_b),
    .io_ci(FullAdder_580_io_ci),
    .io_s(FullAdder_580_io_s),
    .io_co(FullAdder_580_io_co)
  );
  FullAdder FullAdder_581 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_581_io_a),
    .io_b(FullAdder_581_io_b),
    .io_ci(FullAdder_581_io_ci),
    .io_s(FullAdder_581_io_s),
    .io_co(FullAdder_581_io_co)
  );
  FullAdder FullAdder_582 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_582_io_a),
    .io_b(FullAdder_582_io_b),
    .io_ci(FullAdder_582_io_ci),
    .io_s(FullAdder_582_io_s),
    .io_co(FullAdder_582_io_co)
  );
  FullAdder FullAdder_583 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_583_io_a),
    .io_b(FullAdder_583_io_b),
    .io_ci(FullAdder_583_io_ci),
    .io_s(FullAdder_583_io_s),
    .io_co(FullAdder_583_io_co)
  );
  FullAdder FullAdder_584 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_584_io_a),
    .io_b(FullAdder_584_io_b),
    .io_ci(FullAdder_584_io_ci),
    .io_s(FullAdder_584_io_s),
    .io_co(FullAdder_584_io_co)
  );
  FullAdder FullAdder_585 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_585_io_a),
    .io_b(FullAdder_585_io_b),
    .io_ci(FullAdder_585_io_ci),
    .io_s(FullAdder_585_io_s),
    .io_co(FullAdder_585_io_co)
  );
  FullAdder FullAdder_586 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_586_io_a),
    .io_b(FullAdder_586_io_b),
    .io_ci(FullAdder_586_io_ci),
    .io_s(FullAdder_586_io_s),
    .io_co(FullAdder_586_io_co)
  );
  FullAdder FullAdder_587 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_587_io_a),
    .io_b(FullAdder_587_io_b),
    .io_ci(FullAdder_587_io_ci),
    .io_s(FullAdder_587_io_s),
    .io_co(FullAdder_587_io_co)
  );
  FullAdder FullAdder_588 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_588_io_a),
    .io_b(FullAdder_588_io_b),
    .io_ci(FullAdder_588_io_ci),
    .io_s(FullAdder_588_io_s),
    .io_co(FullAdder_588_io_co)
  );
  FullAdder FullAdder_589 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_589_io_a),
    .io_b(FullAdder_589_io_b),
    .io_ci(FullAdder_589_io_ci),
    .io_s(FullAdder_589_io_s),
    .io_co(FullAdder_589_io_co)
  );
  FullAdder FullAdder_590 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_590_io_a),
    .io_b(FullAdder_590_io_b),
    .io_ci(FullAdder_590_io_ci),
    .io_s(FullAdder_590_io_s),
    .io_co(FullAdder_590_io_co)
  );
  FullAdder FullAdder_591 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_591_io_a),
    .io_b(FullAdder_591_io_b),
    .io_ci(FullAdder_591_io_ci),
    .io_s(FullAdder_591_io_s),
    .io_co(FullAdder_591_io_co)
  );
  FullAdder FullAdder_592 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_592_io_a),
    .io_b(FullAdder_592_io_b),
    .io_ci(FullAdder_592_io_ci),
    .io_s(FullAdder_592_io_s),
    .io_co(FullAdder_592_io_co)
  );
  FullAdder FullAdder_593 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_593_io_a),
    .io_b(FullAdder_593_io_b),
    .io_ci(FullAdder_593_io_ci),
    .io_s(FullAdder_593_io_s),
    .io_co(FullAdder_593_io_co)
  );
  FullAdder FullAdder_594 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_594_io_a),
    .io_b(FullAdder_594_io_b),
    .io_ci(FullAdder_594_io_ci),
    .io_s(FullAdder_594_io_s),
    .io_co(FullAdder_594_io_co)
  );
  FullAdder FullAdder_595 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_595_io_a),
    .io_b(FullAdder_595_io_b),
    .io_ci(FullAdder_595_io_ci),
    .io_s(FullAdder_595_io_s),
    .io_co(FullAdder_595_io_co)
  );
  FullAdder FullAdder_596 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_596_io_a),
    .io_b(FullAdder_596_io_b),
    .io_ci(FullAdder_596_io_ci),
    .io_s(FullAdder_596_io_s),
    .io_co(FullAdder_596_io_co)
  );
  FullAdder FullAdder_597 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_597_io_a),
    .io_b(FullAdder_597_io_b),
    .io_ci(FullAdder_597_io_ci),
    .io_s(FullAdder_597_io_s),
    .io_co(FullAdder_597_io_co)
  );
  FullAdder FullAdder_598 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_598_io_a),
    .io_b(FullAdder_598_io_b),
    .io_ci(FullAdder_598_io_ci),
    .io_s(FullAdder_598_io_s),
    .io_co(FullAdder_598_io_co)
  );
  FullAdder FullAdder_599 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_599_io_a),
    .io_b(FullAdder_599_io_b),
    .io_ci(FullAdder_599_io_ci),
    .io_s(FullAdder_599_io_s),
    .io_co(FullAdder_599_io_co)
  );
  FullAdder FullAdder_600 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_600_io_a),
    .io_b(FullAdder_600_io_b),
    .io_ci(FullAdder_600_io_ci),
    .io_s(FullAdder_600_io_s),
    .io_co(FullAdder_600_io_co)
  );
  FullAdder FullAdder_601 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_601_io_a),
    .io_b(FullAdder_601_io_b),
    .io_ci(FullAdder_601_io_ci),
    .io_s(FullAdder_601_io_s),
    .io_co(FullAdder_601_io_co)
  );
  FullAdder FullAdder_602 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_602_io_a),
    .io_b(FullAdder_602_io_b),
    .io_ci(FullAdder_602_io_ci),
    .io_s(FullAdder_602_io_s),
    .io_co(FullAdder_602_io_co)
  );
  FullAdder FullAdder_603 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_603_io_a),
    .io_b(FullAdder_603_io_b),
    .io_ci(FullAdder_603_io_ci),
    .io_s(FullAdder_603_io_s),
    .io_co(FullAdder_603_io_co)
  );
  FullAdder FullAdder_604 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_604_io_a),
    .io_b(FullAdder_604_io_b),
    .io_ci(FullAdder_604_io_ci),
    .io_s(FullAdder_604_io_s),
    .io_co(FullAdder_604_io_co)
  );
  FullAdder FullAdder_605 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_605_io_a),
    .io_b(FullAdder_605_io_b),
    .io_ci(FullAdder_605_io_ci),
    .io_s(FullAdder_605_io_s),
    .io_co(FullAdder_605_io_co)
  );
  FullAdder FullAdder_606 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_606_io_a),
    .io_b(FullAdder_606_io_b),
    .io_ci(FullAdder_606_io_ci),
    .io_s(FullAdder_606_io_s),
    .io_co(FullAdder_606_io_co)
  );
  FullAdder FullAdder_607 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_607_io_a),
    .io_b(FullAdder_607_io_b),
    .io_ci(FullAdder_607_io_ci),
    .io_s(FullAdder_607_io_s),
    .io_co(FullAdder_607_io_co)
  );
  FullAdder FullAdder_608 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_608_io_a),
    .io_b(FullAdder_608_io_b),
    .io_ci(FullAdder_608_io_ci),
    .io_s(FullAdder_608_io_s),
    .io_co(FullAdder_608_io_co)
  );
  FullAdder FullAdder_609 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_609_io_a),
    .io_b(FullAdder_609_io_b),
    .io_ci(FullAdder_609_io_ci),
    .io_s(FullAdder_609_io_s),
    .io_co(FullAdder_609_io_co)
  );
  FullAdder FullAdder_610 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_610_io_a),
    .io_b(FullAdder_610_io_b),
    .io_ci(FullAdder_610_io_ci),
    .io_s(FullAdder_610_io_s),
    .io_co(FullAdder_610_io_co)
  );
  FullAdder FullAdder_611 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_611_io_a),
    .io_b(FullAdder_611_io_b),
    .io_ci(FullAdder_611_io_ci),
    .io_s(FullAdder_611_io_s),
    .io_co(FullAdder_611_io_co)
  );
  FullAdder FullAdder_612 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_612_io_a),
    .io_b(FullAdder_612_io_b),
    .io_ci(FullAdder_612_io_ci),
    .io_s(FullAdder_612_io_s),
    .io_co(FullAdder_612_io_co)
  );
  FullAdder FullAdder_613 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_613_io_a),
    .io_b(FullAdder_613_io_b),
    .io_ci(FullAdder_613_io_ci),
    .io_s(FullAdder_613_io_s),
    .io_co(FullAdder_613_io_co)
  );
  FullAdder FullAdder_614 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_614_io_a),
    .io_b(FullAdder_614_io_b),
    .io_ci(FullAdder_614_io_ci),
    .io_s(FullAdder_614_io_s),
    .io_co(FullAdder_614_io_co)
  );
  FullAdder FullAdder_615 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_615_io_a),
    .io_b(FullAdder_615_io_b),
    .io_ci(FullAdder_615_io_ci),
    .io_s(FullAdder_615_io_s),
    .io_co(FullAdder_615_io_co)
  );
  FullAdder FullAdder_616 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_616_io_a),
    .io_b(FullAdder_616_io_b),
    .io_ci(FullAdder_616_io_ci),
    .io_s(FullAdder_616_io_s),
    .io_co(FullAdder_616_io_co)
  );
  FullAdder FullAdder_617 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_617_io_a),
    .io_b(FullAdder_617_io_b),
    .io_ci(FullAdder_617_io_ci),
    .io_s(FullAdder_617_io_s),
    .io_co(FullAdder_617_io_co)
  );
  FullAdder FullAdder_618 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_618_io_a),
    .io_b(FullAdder_618_io_b),
    .io_ci(FullAdder_618_io_ci),
    .io_s(FullAdder_618_io_s),
    .io_co(FullAdder_618_io_co)
  );
  FullAdder FullAdder_619 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_619_io_a),
    .io_b(FullAdder_619_io_b),
    .io_ci(FullAdder_619_io_ci),
    .io_s(FullAdder_619_io_s),
    .io_co(FullAdder_619_io_co)
  );
  FullAdder FullAdder_620 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_620_io_a),
    .io_b(FullAdder_620_io_b),
    .io_ci(FullAdder_620_io_ci),
    .io_s(FullAdder_620_io_s),
    .io_co(FullAdder_620_io_co)
  );
  FullAdder FullAdder_621 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_621_io_a),
    .io_b(FullAdder_621_io_b),
    .io_ci(FullAdder_621_io_ci),
    .io_s(FullAdder_621_io_s),
    .io_co(FullAdder_621_io_co)
  );
  FullAdder FullAdder_622 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_622_io_a),
    .io_b(FullAdder_622_io_b),
    .io_ci(FullAdder_622_io_ci),
    .io_s(FullAdder_622_io_s),
    .io_co(FullAdder_622_io_co)
  );
  FullAdder FullAdder_623 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_623_io_a),
    .io_b(FullAdder_623_io_b),
    .io_ci(FullAdder_623_io_ci),
    .io_s(FullAdder_623_io_s),
    .io_co(FullAdder_623_io_co)
  );
  FullAdder FullAdder_624 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_624_io_a),
    .io_b(FullAdder_624_io_b),
    .io_ci(FullAdder_624_io_ci),
    .io_s(FullAdder_624_io_s),
    .io_co(FullAdder_624_io_co)
  );
  FullAdder FullAdder_625 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_625_io_a),
    .io_b(FullAdder_625_io_b),
    .io_ci(FullAdder_625_io_ci),
    .io_s(FullAdder_625_io_s),
    .io_co(FullAdder_625_io_co)
  );
  FullAdder FullAdder_626 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_626_io_a),
    .io_b(FullAdder_626_io_b),
    .io_ci(FullAdder_626_io_ci),
    .io_s(FullAdder_626_io_s),
    .io_co(FullAdder_626_io_co)
  );
  FullAdder FullAdder_627 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_627_io_a),
    .io_b(FullAdder_627_io_b),
    .io_ci(FullAdder_627_io_ci),
    .io_s(FullAdder_627_io_s),
    .io_co(FullAdder_627_io_co)
  );
  FullAdder FullAdder_628 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_628_io_a),
    .io_b(FullAdder_628_io_b),
    .io_ci(FullAdder_628_io_ci),
    .io_s(FullAdder_628_io_s),
    .io_co(FullAdder_628_io_co)
  );
  FullAdder FullAdder_629 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_629_io_a),
    .io_b(FullAdder_629_io_b),
    .io_ci(FullAdder_629_io_ci),
    .io_s(FullAdder_629_io_s),
    .io_co(FullAdder_629_io_co)
  );
  HalfAdder HalfAdder_17 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_17_io_a),
    .io_b(HalfAdder_17_io_b),
    .io_s(HalfAdder_17_io_s),
    .io_co(HalfAdder_17_io_co)
  );
  FullAdder FullAdder_630 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_630_io_a),
    .io_b(FullAdder_630_io_b),
    .io_ci(FullAdder_630_io_ci),
    .io_s(FullAdder_630_io_s),
    .io_co(FullAdder_630_io_co)
  );
  FullAdder FullAdder_631 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_631_io_a),
    .io_b(FullAdder_631_io_b),
    .io_ci(FullAdder_631_io_ci),
    .io_s(FullAdder_631_io_s),
    .io_co(FullAdder_631_io_co)
  );
  FullAdder FullAdder_632 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_632_io_a),
    .io_b(FullAdder_632_io_b),
    .io_ci(FullAdder_632_io_ci),
    .io_s(FullAdder_632_io_s),
    .io_co(FullAdder_632_io_co)
  );
  FullAdder FullAdder_633 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_633_io_a),
    .io_b(FullAdder_633_io_b),
    .io_ci(FullAdder_633_io_ci),
    .io_s(FullAdder_633_io_s),
    .io_co(FullAdder_633_io_co)
  );
  FullAdder FullAdder_634 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_634_io_a),
    .io_b(FullAdder_634_io_b),
    .io_ci(FullAdder_634_io_ci),
    .io_s(FullAdder_634_io_s),
    .io_co(FullAdder_634_io_co)
  );
  FullAdder FullAdder_635 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_635_io_a),
    .io_b(FullAdder_635_io_b),
    .io_ci(FullAdder_635_io_ci),
    .io_s(FullAdder_635_io_s),
    .io_co(FullAdder_635_io_co)
  );
  FullAdder FullAdder_636 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_636_io_a),
    .io_b(FullAdder_636_io_b),
    .io_ci(FullAdder_636_io_ci),
    .io_s(FullAdder_636_io_s),
    .io_co(FullAdder_636_io_co)
  );
  FullAdder FullAdder_637 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_637_io_a),
    .io_b(FullAdder_637_io_b),
    .io_ci(FullAdder_637_io_ci),
    .io_s(FullAdder_637_io_s),
    .io_co(FullAdder_637_io_co)
  );
  FullAdder FullAdder_638 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_638_io_a),
    .io_b(FullAdder_638_io_b),
    .io_ci(FullAdder_638_io_ci),
    .io_s(FullAdder_638_io_s),
    .io_co(FullAdder_638_io_co)
  );
  FullAdder FullAdder_639 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_639_io_a),
    .io_b(FullAdder_639_io_b),
    .io_ci(FullAdder_639_io_ci),
    .io_s(FullAdder_639_io_s),
    .io_co(FullAdder_639_io_co)
  );
  FullAdder FullAdder_640 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_640_io_a),
    .io_b(FullAdder_640_io_b),
    .io_ci(FullAdder_640_io_ci),
    .io_s(FullAdder_640_io_s),
    .io_co(FullAdder_640_io_co)
  );
  FullAdder FullAdder_641 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_641_io_a),
    .io_b(FullAdder_641_io_b),
    .io_ci(FullAdder_641_io_ci),
    .io_s(FullAdder_641_io_s),
    .io_co(FullAdder_641_io_co)
  );
  FullAdder FullAdder_642 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_642_io_a),
    .io_b(FullAdder_642_io_b),
    .io_ci(FullAdder_642_io_ci),
    .io_s(FullAdder_642_io_s),
    .io_co(FullAdder_642_io_co)
  );
  FullAdder FullAdder_643 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_643_io_a),
    .io_b(FullAdder_643_io_b),
    .io_ci(FullAdder_643_io_ci),
    .io_s(FullAdder_643_io_s),
    .io_co(FullAdder_643_io_co)
  );
  FullAdder FullAdder_644 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_644_io_a),
    .io_b(FullAdder_644_io_b),
    .io_ci(FullAdder_644_io_ci),
    .io_s(FullAdder_644_io_s),
    .io_co(FullAdder_644_io_co)
  );
  FullAdder FullAdder_645 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_645_io_a),
    .io_b(FullAdder_645_io_b),
    .io_ci(FullAdder_645_io_ci),
    .io_s(FullAdder_645_io_s),
    .io_co(FullAdder_645_io_co)
  );
  FullAdder FullAdder_646 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_646_io_a),
    .io_b(FullAdder_646_io_b),
    .io_ci(FullAdder_646_io_ci),
    .io_s(FullAdder_646_io_s),
    .io_co(FullAdder_646_io_co)
  );
  FullAdder FullAdder_647 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_647_io_a),
    .io_b(FullAdder_647_io_b),
    .io_ci(FullAdder_647_io_ci),
    .io_s(FullAdder_647_io_s),
    .io_co(FullAdder_647_io_co)
  );
  FullAdder FullAdder_648 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_648_io_a),
    .io_b(FullAdder_648_io_b),
    .io_ci(FullAdder_648_io_ci),
    .io_s(FullAdder_648_io_s),
    .io_co(FullAdder_648_io_co)
  );
  FullAdder FullAdder_649 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_649_io_a),
    .io_b(FullAdder_649_io_b),
    .io_ci(FullAdder_649_io_ci),
    .io_s(FullAdder_649_io_s),
    .io_co(FullAdder_649_io_co)
  );
  FullAdder FullAdder_650 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_650_io_a),
    .io_b(FullAdder_650_io_b),
    .io_ci(FullAdder_650_io_ci),
    .io_s(FullAdder_650_io_s),
    .io_co(FullAdder_650_io_co)
  );
  FullAdder FullAdder_651 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_651_io_a),
    .io_b(FullAdder_651_io_b),
    .io_ci(FullAdder_651_io_ci),
    .io_s(FullAdder_651_io_s),
    .io_co(FullAdder_651_io_co)
  );
  FullAdder FullAdder_652 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_652_io_a),
    .io_b(FullAdder_652_io_b),
    .io_ci(FullAdder_652_io_ci),
    .io_s(FullAdder_652_io_s),
    .io_co(FullAdder_652_io_co)
  );
  FullAdder FullAdder_653 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_653_io_a),
    .io_b(FullAdder_653_io_b),
    .io_ci(FullAdder_653_io_ci),
    .io_s(FullAdder_653_io_s),
    .io_co(FullAdder_653_io_co)
  );
  FullAdder FullAdder_654 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_654_io_a),
    .io_b(FullAdder_654_io_b),
    .io_ci(FullAdder_654_io_ci),
    .io_s(FullAdder_654_io_s),
    .io_co(FullAdder_654_io_co)
  );
  FullAdder FullAdder_655 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_655_io_a),
    .io_b(FullAdder_655_io_b),
    .io_ci(FullAdder_655_io_ci),
    .io_s(FullAdder_655_io_s),
    .io_co(FullAdder_655_io_co)
  );
  FullAdder FullAdder_656 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_656_io_a),
    .io_b(FullAdder_656_io_b),
    .io_ci(FullAdder_656_io_ci),
    .io_s(FullAdder_656_io_s),
    .io_co(FullAdder_656_io_co)
  );
  FullAdder FullAdder_657 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_657_io_a),
    .io_b(FullAdder_657_io_b),
    .io_ci(FullAdder_657_io_ci),
    .io_s(FullAdder_657_io_s),
    .io_co(FullAdder_657_io_co)
  );
  FullAdder FullAdder_658 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_658_io_a),
    .io_b(FullAdder_658_io_b),
    .io_ci(FullAdder_658_io_ci),
    .io_s(FullAdder_658_io_s),
    .io_co(FullAdder_658_io_co)
  );
  FullAdder FullAdder_659 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_659_io_a),
    .io_b(FullAdder_659_io_b),
    .io_ci(FullAdder_659_io_ci),
    .io_s(FullAdder_659_io_s),
    .io_co(FullAdder_659_io_co)
  );
  FullAdder FullAdder_660 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_660_io_a),
    .io_b(FullAdder_660_io_b),
    .io_ci(FullAdder_660_io_ci),
    .io_s(FullAdder_660_io_s),
    .io_co(FullAdder_660_io_co)
  );
  FullAdder FullAdder_661 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_661_io_a),
    .io_b(FullAdder_661_io_b),
    .io_ci(FullAdder_661_io_ci),
    .io_s(FullAdder_661_io_s),
    .io_co(FullAdder_661_io_co)
  );
  FullAdder FullAdder_662 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_662_io_a),
    .io_b(FullAdder_662_io_b),
    .io_ci(FullAdder_662_io_ci),
    .io_s(FullAdder_662_io_s),
    .io_co(FullAdder_662_io_co)
  );
  FullAdder FullAdder_663 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_663_io_a),
    .io_b(FullAdder_663_io_b),
    .io_ci(FullAdder_663_io_ci),
    .io_s(FullAdder_663_io_s),
    .io_co(FullAdder_663_io_co)
  );
  FullAdder FullAdder_664 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_664_io_a),
    .io_b(FullAdder_664_io_b),
    .io_ci(FullAdder_664_io_ci),
    .io_s(FullAdder_664_io_s),
    .io_co(FullAdder_664_io_co)
  );
  FullAdder FullAdder_665 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_665_io_a),
    .io_b(FullAdder_665_io_b),
    .io_ci(FullAdder_665_io_ci),
    .io_s(FullAdder_665_io_s),
    .io_co(FullAdder_665_io_co)
  );
  FullAdder FullAdder_666 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_666_io_a),
    .io_b(FullAdder_666_io_b),
    .io_ci(FullAdder_666_io_ci),
    .io_s(FullAdder_666_io_s),
    .io_co(FullAdder_666_io_co)
  );
  FullAdder FullAdder_667 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_667_io_a),
    .io_b(FullAdder_667_io_b),
    .io_ci(FullAdder_667_io_ci),
    .io_s(FullAdder_667_io_s),
    .io_co(FullAdder_667_io_co)
  );
  FullAdder FullAdder_668 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_668_io_a),
    .io_b(FullAdder_668_io_b),
    .io_ci(FullAdder_668_io_ci),
    .io_s(FullAdder_668_io_s),
    .io_co(FullAdder_668_io_co)
  );
  FullAdder FullAdder_669 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_669_io_a),
    .io_b(FullAdder_669_io_b),
    .io_ci(FullAdder_669_io_ci),
    .io_s(FullAdder_669_io_s),
    .io_co(FullAdder_669_io_co)
  );
  FullAdder FullAdder_670 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_670_io_a),
    .io_b(FullAdder_670_io_b),
    .io_ci(FullAdder_670_io_ci),
    .io_s(FullAdder_670_io_s),
    .io_co(FullAdder_670_io_co)
  );
  FullAdder FullAdder_671 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_671_io_a),
    .io_b(FullAdder_671_io_b),
    .io_ci(FullAdder_671_io_ci),
    .io_s(FullAdder_671_io_s),
    .io_co(FullAdder_671_io_co)
  );
  FullAdder FullAdder_672 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_672_io_a),
    .io_b(FullAdder_672_io_b),
    .io_ci(FullAdder_672_io_ci),
    .io_s(FullAdder_672_io_s),
    .io_co(FullAdder_672_io_co)
  );
  FullAdder FullAdder_673 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_673_io_a),
    .io_b(FullAdder_673_io_b),
    .io_ci(FullAdder_673_io_ci),
    .io_s(FullAdder_673_io_s),
    .io_co(FullAdder_673_io_co)
  );
  FullAdder FullAdder_674 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_674_io_a),
    .io_b(FullAdder_674_io_b),
    .io_ci(FullAdder_674_io_ci),
    .io_s(FullAdder_674_io_s),
    .io_co(FullAdder_674_io_co)
  );
  FullAdder FullAdder_675 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_675_io_a),
    .io_b(FullAdder_675_io_b),
    .io_ci(FullAdder_675_io_ci),
    .io_s(FullAdder_675_io_s),
    .io_co(FullAdder_675_io_co)
  );
  FullAdder FullAdder_676 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_676_io_a),
    .io_b(FullAdder_676_io_b),
    .io_ci(FullAdder_676_io_ci),
    .io_s(FullAdder_676_io_s),
    .io_co(FullAdder_676_io_co)
  );
  FullAdder FullAdder_677 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_677_io_a),
    .io_b(FullAdder_677_io_b),
    .io_ci(FullAdder_677_io_ci),
    .io_s(FullAdder_677_io_s),
    .io_co(FullAdder_677_io_co)
  );
  FullAdder FullAdder_678 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_678_io_a),
    .io_b(FullAdder_678_io_b),
    .io_ci(FullAdder_678_io_ci),
    .io_s(FullAdder_678_io_s),
    .io_co(FullAdder_678_io_co)
  );
  FullAdder FullAdder_679 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_679_io_a),
    .io_b(FullAdder_679_io_b),
    .io_ci(FullAdder_679_io_ci),
    .io_s(FullAdder_679_io_s),
    .io_co(FullAdder_679_io_co)
  );
  FullAdder FullAdder_680 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_680_io_a),
    .io_b(FullAdder_680_io_b),
    .io_ci(FullAdder_680_io_ci),
    .io_s(FullAdder_680_io_s),
    .io_co(FullAdder_680_io_co)
  );
  FullAdder FullAdder_681 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_681_io_a),
    .io_b(FullAdder_681_io_b),
    .io_ci(FullAdder_681_io_ci),
    .io_s(FullAdder_681_io_s),
    .io_co(FullAdder_681_io_co)
  );
  FullAdder FullAdder_682 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_682_io_a),
    .io_b(FullAdder_682_io_b),
    .io_ci(FullAdder_682_io_ci),
    .io_s(FullAdder_682_io_s),
    .io_co(FullAdder_682_io_co)
  );
  FullAdder FullAdder_683 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_683_io_a),
    .io_b(FullAdder_683_io_b),
    .io_ci(FullAdder_683_io_ci),
    .io_s(FullAdder_683_io_s),
    .io_co(FullAdder_683_io_co)
  );
  FullAdder FullAdder_684 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_684_io_a),
    .io_b(FullAdder_684_io_b),
    .io_ci(FullAdder_684_io_ci),
    .io_s(FullAdder_684_io_s),
    .io_co(FullAdder_684_io_co)
  );
  FullAdder FullAdder_685 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_685_io_a),
    .io_b(FullAdder_685_io_b),
    .io_ci(FullAdder_685_io_ci),
    .io_s(FullAdder_685_io_s),
    .io_co(FullAdder_685_io_co)
  );
  FullAdder FullAdder_686 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_686_io_a),
    .io_b(FullAdder_686_io_b),
    .io_ci(FullAdder_686_io_ci),
    .io_s(FullAdder_686_io_s),
    .io_co(FullAdder_686_io_co)
  );
  FullAdder FullAdder_687 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_687_io_a),
    .io_b(FullAdder_687_io_b),
    .io_ci(FullAdder_687_io_ci),
    .io_s(FullAdder_687_io_s),
    .io_co(FullAdder_687_io_co)
  );
  FullAdder FullAdder_688 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_688_io_a),
    .io_b(FullAdder_688_io_b),
    .io_ci(FullAdder_688_io_ci),
    .io_s(FullAdder_688_io_s),
    .io_co(FullAdder_688_io_co)
  );
  FullAdder FullAdder_689 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_689_io_a),
    .io_b(FullAdder_689_io_b),
    .io_ci(FullAdder_689_io_ci),
    .io_s(FullAdder_689_io_s),
    .io_co(FullAdder_689_io_co)
  );
  FullAdder FullAdder_690 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_690_io_a),
    .io_b(FullAdder_690_io_b),
    .io_ci(FullAdder_690_io_ci),
    .io_s(FullAdder_690_io_s),
    .io_co(FullAdder_690_io_co)
  );
  FullAdder FullAdder_691 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_691_io_a),
    .io_b(FullAdder_691_io_b),
    .io_ci(FullAdder_691_io_ci),
    .io_s(FullAdder_691_io_s),
    .io_co(FullAdder_691_io_co)
  );
  FullAdder FullAdder_692 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_692_io_a),
    .io_b(FullAdder_692_io_b),
    .io_ci(FullAdder_692_io_ci),
    .io_s(FullAdder_692_io_s),
    .io_co(FullAdder_692_io_co)
  );
  FullAdder FullAdder_693 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_693_io_a),
    .io_b(FullAdder_693_io_b),
    .io_ci(FullAdder_693_io_ci),
    .io_s(FullAdder_693_io_s),
    .io_co(FullAdder_693_io_co)
  );
  FullAdder FullAdder_694 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_694_io_a),
    .io_b(FullAdder_694_io_b),
    .io_ci(FullAdder_694_io_ci),
    .io_s(FullAdder_694_io_s),
    .io_co(FullAdder_694_io_co)
  );
  FullAdder FullAdder_695 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_695_io_a),
    .io_b(FullAdder_695_io_b),
    .io_ci(FullAdder_695_io_ci),
    .io_s(FullAdder_695_io_s),
    .io_co(FullAdder_695_io_co)
  );
  FullAdder FullAdder_696 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_696_io_a),
    .io_b(FullAdder_696_io_b),
    .io_ci(FullAdder_696_io_ci),
    .io_s(FullAdder_696_io_s),
    .io_co(FullAdder_696_io_co)
  );
  FullAdder FullAdder_697 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_697_io_a),
    .io_b(FullAdder_697_io_b),
    .io_ci(FullAdder_697_io_ci),
    .io_s(FullAdder_697_io_s),
    .io_co(FullAdder_697_io_co)
  );
  FullAdder FullAdder_698 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_698_io_a),
    .io_b(FullAdder_698_io_b),
    .io_ci(FullAdder_698_io_ci),
    .io_s(FullAdder_698_io_s),
    .io_co(FullAdder_698_io_co)
  );
  FullAdder FullAdder_699 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_699_io_a),
    .io_b(FullAdder_699_io_b),
    .io_ci(FullAdder_699_io_ci),
    .io_s(FullAdder_699_io_s),
    .io_co(FullAdder_699_io_co)
  );
  FullAdder FullAdder_700 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_700_io_a),
    .io_b(FullAdder_700_io_b),
    .io_ci(FullAdder_700_io_ci),
    .io_s(FullAdder_700_io_s),
    .io_co(FullAdder_700_io_co)
  );
  FullAdder FullAdder_701 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_701_io_a),
    .io_b(FullAdder_701_io_b),
    .io_ci(FullAdder_701_io_ci),
    .io_s(FullAdder_701_io_s),
    .io_co(FullAdder_701_io_co)
  );
  FullAdder FullAdder_702 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_702_io_a),
    .io_b(FullAdder_702_io_b),
    .io_ci(FullAdder_702_io_ci),
    .io_s(FullAdder_702_io_s),
    .io_co(FullAdder_702_io_co)
  );
  FullAdder FullAdder_703 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_703_io_a),
    .io_b(FullAdder_703_io_b),
    .io_ci(FullAdder_703_io_ci),
    .io_s(FullAdder_703_io_s),
    .io_co(FullAdder_703_io_co)
  );
  FullAdder FullAdder_704 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_704_io_a),
    .io_b(FullAdder_704_io_b),
    .io_ci(FullAdder_704_io_ci),
    .io_s(FullAdder_704_io_s),
    .io_co(FullAdder_704_io_co)
  );
  FullAdder FullAdder_705 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_705_io_a),
    .io_b(FullAdder_705_io_b),
    .io_ci(FullAdder_705_io_ci),
    .io_s(FullAdder_705_io_s),
    .io_co(FullAdder_705_io_co)
  );
  FullAdder FullAdder_706 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_706_io_a),
    .io_b(FullAdder_706_io_b),
    .io_ci(FullAdder_706_io_ci),
    .io_s(FullAdder_706_io_s),
    .io_co(FullAdder_706_io_co)
  );
  FullAdder FullAdder_707 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_707_io_a),
    .io_b(FullAdder_707_io_b),
    .io_ci(FullAdder_707_io_ci),
    .io_s(FullAdder_707_io_s),
    .io_co(FullAdder_707_io_co)
  );
  FullAdder FullAdder_708 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_708_io_a),
    .io_b(FullAdder_708_io_b),
    .io_ci(FullAdder_708_io_ci),
    .io_s(FullAdder_708_io_s),
    .io_co(FullAdder_708_io_co)
  );
  FullAdder FullAdder_709 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_709_io_a),
    .io_b(FullAdder_709_io_b),
    .io_ci(FullAdder_709_io_ci),
    .io_s(FullAdder_709_io_s),
    .io_co(FullAdder_709_io_co)
  );
  FullAdder FullAdder_710 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_710_io_a),
    .io_b(FullAdder_710_io_b),
    .io_ci(FullAdder_710_io_ci),
    .io_s(FullAdder_710_io_s),
    .io_co(FullAdder_710_io_co)
  );
  FullAdder FullAdder_711 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_711_io_a),
    .io_b(FullAdder_711_io_b),
    .io_ci(FullAdder_711_io_ci),
    .io_s(FullAdder_711_io_s),
    .io_co(FullAdder_711_io_co)
  );
  FullAdder FullAdder_712 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_712_io_a),
    .io_b(FullAdder_712_io_b),
    .io_ci(FullAdder_712_io_ci),
    .io_s(FullAdder_712_io_s),
    .io_co(FullAdder_712_io_co)
  );
  HalfAdder HalfAdder_18 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_18_io_a),
    .io_b(HalfAdder_18_io_b),
    .io_s(HalfAdder_18_io_s),
    .io_co(HalfAdder_18_io_co)
  );
  FullAdder FullAdder_713 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_713_io_a),
    .io_b(FullAdder_713_io_b),
    .io_ci(FullAdder_713_io_ci),
    .io_s(FullAdder_713_io_s),
    .io_co(FullAdder_713_io_co)
  );
  FullAdder FullAdder_714 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_714_io_a),
    .io_b(FullAdder_714_io_b),
    .io_ci(FullAdder_714_io_ci),
    .io_s(FullAdder_714_io_s),
    .io_co(FullAdder_714_io_co)
  );
  FullAdder FullAdder_715 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_715_io_a),
    .io_b(FullAdder_715_io_b),
    .io_ci(FullAdder_715_io_ci),
    .io_s(FullAdder_715_io_s),
    .io_co(FullAdder_715_io_co)
  );
  FullAdder FullAdder_716 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_716_io_a),
    .io_b(FullAdder_716_io_b),
    .io_ci(FullAdder_716_io_ci),
    .io_s(FullAdder_716_io_s),
    .io_co(FullAdder_716_io_co)
  );
  FullAdder FullAdder_717 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_717_io_a),
    .io_b(FullAdder_717_io_b),
    .io_ci(FullAdder_717_io_ci),
    .io_s(FullAdder_717_io_s),
    .io_co(FullAdder_717_io_co)
  );
  FullAdder FullAdder_718 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_718_io_a),
    .io_b(FullAdder_718_io_b),
    .io_ci(FullAdder_718_io_ci),
    .io_s(FullAdder_718_io_s),
    .io_co(FullAdder_718_io_co)
  );
  FullAdder FullAdder_719 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_719_io_a),
    .io_b(FullAdder_719_io_b),
    .io_ci(FullAdder_719_io_ci),
    .io_s(FullAdder_719_io_s),
    .io_co(FullAdder_719_io_co)
  );
  FullAdder FullAdder_720 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_720_io_a),
    .io_b(FullAdder_720_io_b),
    .io_ci(FullAdder_720_io_ci),
    .io_s(FullAdder_720_io_s),
    .io_co(FullAdder_720_io_co)
  );
  FullAdder FullAdder_721 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_721_io_a),
    .io_b(FullAdder_721_io_b),
    .io_ci(FullAdder_721_io_ci),
    .io_s(FullAdder_721_io_s),
    .io_co(FullAdder_721_io_co)
  );
  FullAdder FullAdder_722 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_722_io_a),
    .io_b(FullAdder_722_io_b),
    .io_ci(FullAdder_722_io_ci),
    .io_s(FullAdder_722_io_s),
    .io_co(FullAdder_722_io_co)
  );
  FullAdder FullAdder_723 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_723_io_a),
    .io_b(FullAdder_723_io_b),
    .io_ci(FullAdder_723_io_ci),
    .io_s(FullAdder_723_io_s),
    .io_co(FullAdder_723_io_co)
  );
  FullAdder FullAdder_724 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_724_io_a),
    .io_b(FullAdder_724_io_b),
    .io_ci(FullAdder_724_io_ci),
    .io_s(FullAdder_724_io_s),
    .io_co(FullAdder_724_io_co)
  );
  FullAdder FullAdder_725 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_725_io_a),
    .io_b(FullAdder_725_io_b),
    .io_ci(FullAdder_725_io_ci),
    .io_s(FullAdder_725_io_s),
    .io_co(FullAdder_725_io_co)
  );
  FullAdder FullAdder_726 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_726_io_a),
    .io_b(FullAdder_726_io_b),
    .io_ci(FullAdder_726_io_ci),
    .io_s(FullAdder_726_io_s),
    .io_co(FullAdder_726_io_co)
  );
  FullAdder FullAdder_727 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_727_io_a),
    .io_b(FullAdder_727_io_b),
    .io_ci(FullAdder_727_io_ci),
    .io_s(FullAdder_727_io_s),
    .io_co(FullAdder_727_io_co)
  );
  FullAdder FullAdder_728 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_728_io_a),
    .io_b(FullAdder_728_io_b),
    .io_ci(FullAdder_728_io_ci),
    .io_s(FullAdder_728_io_s),
    .io_co(FullAdder_728_io_co)
  );
  FullAdder FullAdder_729 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_729_io_a),
    .io_b(FullAdder_729_io_b),
    .io_ci(FullAdder_729_io_ci),
    .io_s(FullAdder_729_io_s),
    .io_co(FullAdder_729_io_co)
  );
  FullAdder FullAdder_730 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_730_io_a),
    .io_b(FullAdder_730_io_b),
    .io_ci(FullAdder_730_io_ci),
    .io_s(FullAdder_730_io_s),
    .io_co(FullAdder_730_io_co)
  );
  FullAdder FullAdder_731 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_731_io_a),
    .io_b(FullAdder_731_io_b),
    .io_ci(FullAdder_731_io_ci),
    .io_s(FullAdder_731_io_s),
    .io_co(FullAdder_731_io_co)
  );
  FullAdder FullAdder_732 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_732_io_a),
    .io_b(FullAdder_732_io_b),
    .io_ci(FullAdder_732_io_ci),
    .io_s(FullAdder_732_io_s),
    .io_co(FullAdder_732_io_co)
  );
  FullAdder FullAdder_733 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_733_io_a),
    .io_b(FullAdder_733_io_b),
    .io_ci(FullAdder_733_io_ci),
    .io_s(FullAdder_733_io_s),
    .io_co(FullAdder_733_io_co)
  );
  FullAdder FullAdder_734 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_734_io_a),
    .io_b(FullAdder_734_io_b),
    .io_ci(FullAdder_734_io_ci),
    .io_s(FullAdder_734_io_s),
    .io_co(FullAdder_734_io_co)
  );
  FullAdder FullAdder_735 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_735_io_a),
    .io_b(FullAdder_735_io_b),
    .io_ci(FullAdder_735_io_ci),
    .io_s(FullAdder_735_io_s),
    .io_co(FullAdder_735_io_co)
  );
  FullAdder FullAdder_736 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_736_io_a),
    .io_b(FullAdder_736_io_b),
    .io_ci(FullAdder_736_io_ci),
    .io_s(FullAdder_736_io_s),
    .io_co(FullAdder_736_io_co)
  );
  FullAdder FullAdder_737 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_737_io_a),
    .io_b(FullAdder_737_io_b),
    .io_ci(FullAdder_737_io_ci),
    .io_s(FullAdder_737_io_s),
    .io_co(FullAdder_737_io_co)
  );
  FullAdder FullAdder_738 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_738_io_a),
    .io_b(FullAdder_738_io_b),
    .io_ci(FullAdder_738_io_ci),
    .io_s(FullAdder_738_io_s),
    .io_co(FullAdder_738_io_co)
  );
  FullAdder FullAdder_739 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_739_io_a),
    .io_b(FullAdder_739_io_b),
    .io_ci(FullAdder_739_io_ci),
    .io_s(FullAdder_739_io_s),
    .io_co(FullAdder_739_io_co)
  );
  FullAdder FullAdder_740 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_740_io_a),
    .io_b(FullAdder_740_io_b),
    .io_ci(FullAdder_740_io_ci),
    .io_s(FullAdder_740_io_s),
    .io_co(FullAdder_740_io_co)
  );
  FullAdder FullAdder_741 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_741_io_a),
    .io_b(FullAdder_741_io_b),
    .io_ci(FullAdder_741_io_ci),
    .io_s(FullAdder_741_io_s),
    .io_co(FullAdder_741_io_co)
  );
  FullAdder FullAdder_742 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_742_io_a),
    .io_b(FullAdder_742_io_b),
    .io_ci(FullAdder_742_io_ci),
    .io_s(FullAdder_742_io_s),
    .io_co(FullAdder_742_io_co)
  );
  FullAdder FullAdder_743 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_743_io_a),
    .io_b(FullAdder_743_io_b),
    .io_ci(FullAdder_743_io_ci),
    .io_s(FullAdder_743_io_s),
    .io_co(FullAdder_743_io_co)
  );
  FullAdder FullAdder_744 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_744_io_a),
    .io_b(FullAdder_744_io_b),
    .io_ci(FullAdder_744_io_ci),
    .io_s(FullAdder_744_io_s),
    .io_co(FullAdder_744_io_co)
  );
  FullAdder FullAdder_745 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_745_io_a),
    .io_b(FullAdder_745_io_b),
    .io_ci(FullAdder_745_io_ci),
    .io_s(FullAdder_745_io_s),
    .io_co(FullAdder_745_io_co)
  );
  FullAdder FullAdder_746 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_746_io_a),
    .io_b(FullAdder_746_io_b),
    .io_ci(FullAdder_746_io_ci),
    .io_s(FullAdder_746_io_s),
    .io_co(FullAdder_746_io_co)
  );
  FullAdder FullAdder_747 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_747_io_a),
    .io_b(FullAdder_747_io_b),
    .io_ci(FullAdder_747_io_ci),
    .io_s(FullAdder_747_io_s),
    .io_co(FullAdder_747_io_co)
  );
  FullAdder FullAdder_748 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_748_io_a),
    .io_b(FullAdder_748_io_b),
    .io_ci(FullAdder_748_io_ci),
    .io_s(FullAdder_748_io_s),
    .io_co(FullAdder_748_io_co)
  );
  FullAdder FullAdder_749 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_749_io_a),
    .io_b(FullAdder_749_io_b),
    .io_ci(FullAdder_749_io_ci),
    .io_s(FullAdder_749_io_s),
    .io_co(FullAdder_749_io_co)
  );
  FullAdder FullAdder_750 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_750_io_a),
    .io_b(FullAdder_750_io_b),
    .io_ci(FullAdder_750_io_ci),
    .io_s(FullAdder_750_io_s),
    .io_co(FullAdder_750_io_co)
  );
  FullAdder FullAdder_751 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_751_io_a),
    .io_b(FullAdder_751_io_b),
    .io_ci(FullAdder_751_io_ci),
    .io_s(FullAdder_751_io_s),
    .io_co(FullAdder_751_io_co)
  );
  FullAdder FullAdder_752 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_752_io_a),
    .io_b(FullAdder_752_io_b),
    .io_ci(FullAdder_752_io_ci),
    .io_s(FullAdder_752_io_s),
    .io_co(FullAdder_752_io_co)
  );
  FullAdder FullAdder_753 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_753_io_a),
    .io_b(FullAdder_753_io_b),
    .io_ci(FullAdder_753_io_ci),
    .io_s(FullAdder_753_io_s),
    .io_co(FullAdder_753_io_co)
  );
  FullAdder FullAdder_754 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_754_io_a),
    .io_b(FullAdder_754_io_b),
    .io_ci(FullAdder_754_io_ci),
    .io_s(FullAdder_754_io_s),
    .io_co(FullAdder_754_io_co)
  );
  FullAdder FullAdder_755 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_755_io_a),
    .io_b(FullAdder_755_io_b),
    .io_ci(FullAdder_755_io_ci),
    .io_s(FullAdder_755_io_s),
    .io_co(FullAdder_755_io_co)
  );
  FullAdder FullAdder_756 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_756_io_a),
    .io_b(FullAdder_756_io_b),
    .io_ci(FullAdder_756_io_ci),
    .io_s(FullAdder_756_io_s),
    .io_co(FullAdder_756_io_co)
  );
  FullAdder FullAdder_757 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_757_io_a),
    .io_b(FullAdder_757_io_b),
    .io_ci(FullAdder_757_io_ci),
    .io_s(FullAdder_757_io_s),
    .io_co(FullAdder_757_io_co)
  );
  FullAdder FullAdder_758 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_758_io_a),
    .io_b(FullAdder_758_io_b),
    .io_ci(FullAdder_758_io_ci),
    .io_s(FullAdder_758_io_s),
    .io_co(FullAdder_758_io_co)
  );
  FullAdder FullAdder_759 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_759_io_a),
    .io_b(FullAdder_759_io_b),
    .io_ci(FullAdder_759_io_ci),
    .io_s(FullAdder_759_io_s),
    .io_co(FullAdder_759_io_co)
  );
  FullAdder FullAdder_760 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_760_io_a),
    .io_b(FullAdder_760_io_b),
    .io_ci(FullAdder_760_io_ci),
    .io_s(FullAdder_760_io_s),
    .io_co(FullAdder_760_io_co)
  );
  FullAdder FullAdder_761 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_761_io_a),
    .io_b(FullAdder_761_io_b),
    .io_ci(FullAdder_761_io_ci),
    .io_s(FullAdder_761_io_s),
    .io_co(FullAdder_761_io_co)
  );
  FullAdder FullAdder_762 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_762_io_a),
    .io_b(FullAdder_762_io_b),
    .io_ci(FullAdder_762_io_ci),
    .io_s(FullAdder_762_io_s),
    .io_co(FullAdder_762_io_co)
  );
  FullAdder FullAdder_763 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_763_io_a),
    .io_b(FullAdder_763_io_b),
    .io_ci(FullAdder_763_io_ci),
    .io_s(FullAdder_763_io_s),
    .io_co(FullAdder_763_io_co)
  );
  FullAdder FullAdder_764 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_764_io_a),
    .io_b(FullAdder_764_io_b),
    .io_ci(FullAdder_764_io_ci),
    .io_s(FullAdder_764_io_s),
    .io_co(FullAdder_764_io_co)
  );
  FullAdder FullAdder_765 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_765_io_a),
    .io_b(FullAdder_765_io_b),
    .io_ci(FullAdder_765_io_ci),
    .io_s(FullAdder_765_io_s),
    .io_co(FullAdder_765_io_co)
  );
  FullAdder FullAdder_766 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_766_io_a),
    .io_b(FullAdder_766_io_b),
    .io_ci(FullAdder_766_io_ci),
    .io_s(FullAdder_766_io_s),
    .io_co(FullAdder_766_io_co)
  );
  FullAdder FullAdder_767 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_767_io_a),
    .io_b(FullAdder_767_io_b),
    .io_ci(FullAdder_767_io_ci),
    .io_s(FullAdder_767_io_s),
    .io_co(FullAdder_767_io_co)
  );
  FullAdder FullAdder_768 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_768_io_a),
    .io_b(FullAdder_768_io_b),
    .io_ci(FullAdder_768_io_ci),
    .io_s(FullAdder_768_io_s),
    .io_co(FullAdder_768_io_co)
  );
  FullAdder FullAdder_769 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_769_io_a),
    .io_b(FullAdder_769_io_b),
    .io_ci(FullAdder_769_io_ci),
    .io_s(FullAdder_769_io_s),
    .io_co(FullAdder_769_io_co)
  );
  FullAdder FullAdder_770 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_770_io_a),
    .io_b(FullAdder_770_io_b),
    .io_ci(FullAdder_770_io_ci),
    .io_s(FullAdder_770_io_s),
    .io_co(FullAdder_770_io_co)
  );
  FullAdder FullAdder_771 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_771_io_a),
    .io_b(FullAdder_771_io_b),
    .io_ci(FullAdder_771_io_ci),
    .io_s(FullAdder_771_io_s),
    .io_co(FullAdder_771_io_co)
  );
  HalfAdder HalfAdder_19 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_19_io_a),
    .io_b(HalfAdder_19_io_b),
    .io_s(HalfAdder_19_io_s),
    .io_co(HalfAdder_19_io_co)
  );
  FullAdder FullAdder_772 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_772_io_a),
    .io_b(FullAdder_772_io_b),
    .io_ci(FullAdder_772_io_ci),
    .io_s(FullAdder_772_io_s),
    .io_co(FullAdder_772_io_co)
  );
  FullAdder FullAdder_773 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_773_io_a),
    .io_b(FullAdder_773_io_b),
    .io_ci(FullAdder_773_io_ci),
    .io_s(FullAdder_773_io_s),
    .io_co(FullAdder_773_io_co)
  );
  FullAdder FullAdder_774 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_774_io_a),
    .io_b(FullAdder_774_io_b),
    .io_ci(FullAdder_774_io_ci),
    .io_s(FullAdder_774_io_s),
    .io_co(FullAdder_774_io_co)
  );
  FullAdder FullAdder_775 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_775_io_a),
    .io_b(FullAdder_775_io_b),
    .io_ci(FullAdder_775_io_ci),
    .io_s(FullAdder_775_io_s),
    .io_co(FullAdder_775_io_co)
  );
  FullAdder FullAdder_776 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_776_io_a),
    .io_b(FullAdder_776_io_b),
    .io_ci(FullAdder_776_io_ci),
    .io_s(FullAdder_776_io_s),
    .io_co(FullAdder_776_io_co)
  );
  FullAdder FullAdder_777 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_777_io_a),
    .io_b(FullAdder_777_io_b),
    .io_ci(FullAdder_777_io_ci),
    .io_s(FullAdder_777_io_s),
    .io_co(FullAdder_777_io_co)
  );
  FullAdder FullAdder_778 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_778_io_a),
    .io_b(FullAdder_778_io_b),
    .io_ci(FullAdder_778_io_ci),
    .io_s(FullAdder_778_io_s),
    .io_co(FullAdder_778_io_co)
  );
  FullAdder FullAdder_779 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_779_io_a),
    .io_b(FullAdder_779_io_b),
    .io_ci(FullAdder_779_io_ci),
    .io_s(FullAdder_779_io_s),
    .io_co(FullAdder_779_io_co)
  );
  FullAdder FullAdder_780 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_780_io_a),
    .io_b(FullAdder_780_io_b),
    .io_ci(FullAdder_780_io_ci),
    .io_s(FullAdder_780_io_s),
    .io_co(FullAdder_780_io_co)
  );
  FullAdder FullAdder_781 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_781_io_a),
    .io_b(FullAdder_781_io_b),
    .io_ci(FullAdder_781_io_ci),
    .io_s(FullAdder_781_io_s),
    .io_co(FullAdder_781_io_co)
  );
  FullAdder FullAdder_782 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_782_io_a),
    .io_b(FullAdder_782_io_b),
    .io_ci(FullAdder_782_io_ci),
    .io_s(FullAdder_782_io_s),
    .io_co(FullAdder_782_io_co)
  );
  FullAdder FullAdder_783 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_783_io_a),
    .io_b(FullAdder_783_io_b),
    .io_ci(FullAdder_783_io_ci),
    .io_s(FullAdder_783_io_s),
    .io_co(FullAdder_783_io_co)
  );
  FullAdder FullAdder_784 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_784_io_a),
    .io_b(FullAdder_784_io_b),
    .io_ci(FullAdder_784_io_ci),
    .io_s(FullAdder_784_io_s),
    .io_co(FullAdder_784_io_co)
  );
  FullAdder FullAdder_785 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_785_io_a),
    .io_b(FullAdder_785_io_b),
    .io_ci(FullAdder_785_io_ci),
    .io_s(FullAdder_785_io_s),
    .io_co(FullAdder_785_io_co)
  );
  FullAdder FullAdder_786 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_786_io_a),
    .io_b(FullAdder_786_io_b),
    .io_ci(FullAdder_786_io_ci),
    .io_s(FullAdder_786_io_s),
    .io_co(FullAdder_786_io_co)
  );
  FullAdder FullAdder_787 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_787_io_a),
    .io_b(FullAdder_787_io_b),
    .io_ci(FullAdder_787_io_ci),
    .io_s(FullAdder_787_io_s),
    .io_co(FullAdder_787_io_co)
  );
  FullAdder FullAdder_788 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_788_io_a),
    .io_b(FullAdder_788_io_b),
    .io_ci(FullAdder_788_io_ci),
    .io_s(FullAdder_788_io_s),
    .io_co(FullAdder_788_io_co)
  );
  FullAdder FullAdder_789 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_789_io_a),
    .io_b(FullAdder_789_io_b),
    .io_ci(FullAdder_789_io_ci),
    .io_s(FullAdder_789_io_s),
    .io_co(FullAdder_789_io_co)
  );
  FullAdder FullAdder_790 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_790_io_a),
    .io_b(FullAdder_790_io_b),
    .io_ci(FullAdder_790_io_ci),
    .io_s(FullAdder_790_io_s),
    .io_co(FullAdder_790_io_co)
  );
  FullAdder FullAdder_791 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_791_io_a),
    .io_b(FullAdder_791_io_b),
    .io_ci(FullAdder_791_io_ci),
    .io_s(FullAdder_791_io_s),
    .io_co(FullAdder_791_io_co)
  );
  FullAdder FullAdder_792 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_792_io_a),
    .io_b(FullAdder_792_io_b),
    .io_ci(FullAdder_792_io_ci),
    .io_s(FullAdder_792_io_s),
    .io_co(FullAdder_792_io_co)
  );
  FullAdder FullAdder_793 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_793_io_a),
    .io_b(FullAdder_793_io_b),
    .io_ci(FullAdder_793_io_ci),
    .io_s(FullAdder_793_io_s),
    .io_co(FullAdder_793_io_co)
  );
  FullAdder FullAdder_794 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_794_io_a),
    .io_b(FullAdder_794_io_b),
    .io_ci(FullAdder_794_io_ci),
    .io_s(FullAdder_794_io_s),
    .io_co(FullAdder_794_io_co)
  );
  FullAdder FullAdder_795 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_795_io_a),
    .io_b(FullAdder_795_io_b),
    .io_ci(FullAdder_795_io_ci),
    .io_s(FullAdder_795_io_s),
    .io_co(FullAdder_795_io_co)
  );
  FullAdder FullAdder_796 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_796_io_a),
    .io_b(FullAdder_796_io_b),
    .io_ci(FullAdder_796_io_ci),
    .io_s(FullAdder_796_io_s),
    .io_co(FullAdder_796_io_co)
  );
  FullAdder FullAdder_797 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_797_io_a),
    .io_b(FullAdder_797_io_b),
    .io_ci(FullAdder_797_io_ci),
    .io_s(FullAdder_797_io_s),
    .io_co(FullAdder_797_io_co)
  );
  FullAdder FullAdder_798 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_798_io_a),
    .io_b(FullAdder_798_io_b),
    .io_ci(FullAdder_798_io_ci),
    .io_s(FullAdder_798_io_s),
    .io_co(FullAdder_798_io_co)
  );
  FullAdder FullAdder_799 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_799_io_a),
    .io_b(FullAdder_799_io_b),
    .io_ci(FullAdder_799_io_ci),
    .io_s(FullAdder_799_io_s),
    .io_co(FullAdder_799_io_co)
  );
  FullAdder FullAdder_800 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_800_io_a),
    .io_b(FullAdder_800_io_b),
    .io_ci(FullAdder_800_io_ci),
    .io_s(FullAdder_800_io_s),
    .io_co(FullAdder_800_io_co)
  );
  FullAdder FullAdder_801 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_801_io_a),
    .io_b(FullAdder_801_io_b),
    .io_ci(FullAdder_801_io_ci),
    .io_s(FullAdder_801_io_s),
    .io_co(FullAdder_801_io_co)
  );
  FullAdder FullAdder_802 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_802_io_a),
    .io_b(FullAdder_802_io_b),
    .io_ci(FullAdder_802_io_ci),
    .io_s(FullAdder_802_io_s),
    .io_co(FullAdder_802_io_co)
  );
  FullAdder FullAdder_803 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_803_io_a),
    .io_b(FullAdder_803_io_b),
    .io_ci(FullAdder_803_io_ci),
    .io_s(FullAdder_803_io_s),
    .io_co(FullAdder_803_io_co)
  );
  FullAdder FullAdder_804 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_804_io_a),
    .io_b(FullAdder_804_io_b),
    .io_ci(FullAdder_804_io_ci),
    .io_s(FullAdder_804_io_s),
    .io_co(FullAdder_804_io_co)
  );
  FullAdder FullAdder_805 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_805_io_a),
    .io_b(FullAdder_805_io_b),
    .io_ci(FullAdder_805_io_ci),
    .io_s(FullAdder_805_io_s),
    .io_co(FullAdder_805_io_co)
  );
  FullAdder FullAdder_806 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_806_io_a),
    .io_b(FullAdder_806_io_b),
    .io_ci(FullAdder_806_io_ci),
    .io_s(FullAdder_806_io_s),
    .io_co(FullAdder_806_io_co)
  );
  FullAdder FullAdder_807 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_807_io_a),
    .io_b(FullAdder_807_io_b),
    .io_ci(FullAdder_807_io_ci),
    .io_s(FullAdder_807_io_s),
    .io_co(FullAdder_807_io_co)
  );
  FullAdder FullAdder_808 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_808_io_a),
    .io_b(FullAdder_808_io_b),
    .io_ci(FullAdder_808_io_ci),
    .io_s(FullAdder_808_io_s),
    .io_co(FullAdder_808_io_co)
  );
  FullAdder FullAdder_809 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_809_io_a),
    .io_b(FullAdder_809_io_b),
    .io_ci(FullAdder_809_io_ci),
    .io_s(FullAdder_809_io_s),
    .io_co(FullAdder_809_io_co)
  );
  FullAdder FullAdder_810 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_810_io_a),
    .io_b(FullAdder_810_io_b),
    .io_ci(FullAdder_810_io_ci),
    .io_s(FullAdder_810_io_s),
    .io_co(FullAdder_810_io_co)
  );
  FullAdder FullAdder_811 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_811_io_a),
    .io_b(FullAdder_811_io_b),
    .io_ci(FullAdder_811_io_ci),
    .io_s(FullAdder_811_io_s),
    .io_co(FullAdder_811_io_co)
  );
  FullAdder FullAdder_812 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_812_io_a),
    .io_b(FullAdder_812_io_b),
    .io_ci(FullAdder_812_io_ci),
    .io_s(FullAdder_812_io_s),
    .io_co(FullAdder_812_io_co)
  );
  FullAdder FullAdder_813 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_813_io_a),
    .io_b(FullAdder_813_io_b),
    .io_ci(FullAdder_813_io_ci),
    .io_s(FullAdder_813_io_s),
    .io_co(FullAdder_813_io_co)
  );
  FullAdder FullAdder_814 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_814_io_a),
    .io_b(FullAdder_814_io_b),
    .io_ci(FullAdder_814_io_ci),
    .io_s(FullAdder_814_io_s),
    .io_co(FullAdder_814_io_co)
  );
  FullAdder FullAdder_815 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_815_io_a),
    .io_b(FullAdder_815_io_b),
    .io_ci(FullAdder_815_io_ci),
    .io_s(FullAdder_815_io_s),
    .io_co(FullAdder_815_io_co)
  );
  FullAdder FullAdder_816 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_816_io_a),
    .io_b(FullAdder_816_io_b),
    .io_ci(FullAdder_816_io_ci),
    .io_s(FullAdder_816_io_s),
    .io_co(FullAdder_816_io_co)
  );
  FullAdder FullAdder_817 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_817_io_a),
    .io_b(FullAdder_817_io_b),
    .io_ci(FullAdder_817_io_ci),
    .io_s(FullAdder_817_io_s),
    .io_co(FullAdder_817_io_co)
  );
  FullAdder FullAdder_818 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_818_io_a),
    .io_b(FullAdder_818_io_b),
    .io_ci(FullAdder_818_io_ci),
    .io_s(FullAdder_818_io_s),
    .io_co(FullAdder_818_io_co)
  );
  FullAdder FullAdder_819 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_819_io_a),
    .io_b(FullAdder_819_io_b),
    .io_ci(FullAdder_819_io_ci),
    .io_s(FullAdder_819_io_s),
    .io_co(FullAdder_819_io_co)
  );
  FullAdder FullAdder_820 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_820_io_a),
    .io_b(FullAdder_820_io_b),
    .io_ci(FullAdder_820_io_ci),
    .io_s(FullAdder_820_io_s),
    .io_co(FullAdder_820_io_co)
  );
  FullAdder FullAdder_821 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_821_io_a),
    .io_b(FullAdder_821_io_b),
    .io_ci(FullAdder_821_io_ci),
    .io_s(FullAdder_821_io_s),
    .io_co(FullAdder_821_io_co)
  );
  FullAdder FullAdder_822 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_822_io_a),
    .io_b(FullAdder_822_io_b),
    .io_ci(FullAdder_822_io_ci),
    .io_s(FullAdder_822_io_s),
    .io_co(FullAdder_822_io_co)
  );
  FullAdder FullAdder_823 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_823_io_a),
    .io_b(FullAdder_823_io_b),
    .io_ci(FullAdder_823_io_ci),
    .io_s(FullAdder_823_io_s),
    .io_co(FullAdder_823_io_co)
  );
  FullAdder FullAdder_824 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_824_io_a),
    .io_b(FullAdder_824_io_b),
    .io_ci(FullAdder_824_io_ci),
    .io_s(FullAdder_824_io_s),
    .io_co(FullAdder_824_io_co)
  );
  FullAdder FullAdder_825 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_825_io_a),
    .io_b(FullAdder_825_io_b),
    .io_ci(FullAdder_825_io_ci),
    .io_s(FullAdder_825_io_s),
    .io_co(FullAdder_825_io_co)
  );
  FullAdder FullAdder_826 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_826_io_a),
    .io_b(FullAdder_826_io_b),
    .io_ci(FullAdder_826_io_ci),
    .io_s(FullAdder_826_io_s),
    .io_co(FullAdder_826_io_co)
  );
  FullAdder FullAdder_827 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_827_io_a),
    .io_b(FullAdder_827_io_b),
    .io_ci(FullAdder_827_io_ci),
    .io_s(FullAdder_827_io_s),
    .io_co(FullAdder_827_io_co)
  );
  FullAdder FullAdder_828 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_828_io_a),
    .io_b(FullAdder_828_io_b),
    .io_ci(FullAdder_828_io_ci),
    .io_s(FullAdder_828_io_s),
    .io_co(FullAdder_828_io_co)
  );
  FullAdder FullAdder_829 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_829_io_a),
    .io_b(FullAdder_829_io_b),
    .io_ci(FullAdder_829_io_ci),
    .io_s(FullAdder_829_io_s),
    .io_co(FullAdder_829_io_co)
  );
  FullAdder FullAdder_830 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_830_io_a),
    .io_b(FullAdder_830_io_b),
    .io_ci(FullAdder_830_io_ci),
    .io_s(FullAdder_830_io_s),
    .io_co(FullAdder_830_io_co)
  );
  FullAdder FullAdder_831 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_831_io_a),
    .io_b(FullAdder_831_io_b),
    .io_ci(FullAdder_831_io_ci),
    .io_s(FullAdder_831_io_s),
    .io_co(FullAdder_831_io_co)
  );
  FullAdder FullAdder_832 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_832_io_a),
    .io_b(FullAdder_832_io_b),
    .io_ci(FullAdder_832_io_ci),
    .io_s(FullAdder_832_io_s),
    .io_co(FullAdder_832_io_co)
  );
  FullAdder FullAdder_833 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_833_io_a),
    .io_b(FullAdder_833_io_b),
    .io_ci(FullAdder_833_io_ci),
    .io_s(FullAdder_833_io_s),
    .io_co(FullAdder_833_io_co)
  );
  FullAdder FullAdder_834 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_834_io_a),
    .io_b(FullAdder_834_io_b),
    .io_ci(FullAdder_834_io_ci),
    .io_s(FullAdder_834_io_s),
    .io_co(FullAdder_834_io_co)
  );
  FullAdder FullAdder_835 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_835_io_a),
    .io_b(FullAdder_835_io_b),
    .io_ci(FullAdder_835_io_ci),
    .io_s(FullAdder_835_io_s),
    .io_co(FullAdder_835_io_co)
  );
  FullAdder FullAdder_836 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_836_io_a),
    .io_b(FullAdder_836_io_b),
    .io_ci(FullAdder_836_io_ci),
    .io_s(FullAdder_836_io_s),
    .io_co(FullAdder_836_io_co)
  );
  FullAdder FullAdder_837 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_837_io_a),
    .io_b(FullAdder_837_io_b),
    .io_ci(FullAdder_837_io_ci),
    .io_s(FullAdder_837_io_s),
    .io_co(FullAdder_837_io_co)
  );
  FullAdder FullAdder_838 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_838_io_a),
    .io_b(FullAdder_838_io_b),
    .io_ci(FullAdder_838_io_ci),
    .io_s(FullAdder_838_io_s),
    .io_co(FullAdder_838_io_co)
  );
  FullAdder FullAdder_839 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_839_io_a),
    .io_b(FullAdder_839_io_b),
    .io_ci(FullAdder_839_io_ci),
    .io_s(FullAdder_839_io_s),
    .io_co(FullAdder_839_io_co)
  );
  FullAdder FullAdder_840 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_840_io_a),
    .io_b(FullAdder_840_io_b),
    .io_ci(FullAdder_840_io_ci),
    .io_s(FullAdder_840_io_s),
    .io_co(FullAdder_840_io_co)
  );
  FullAdder FullAdder_841 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_841_io_a),
    .io_b(FullAdder_841_io_b),
    .io_ci(FullAdder_841_io_ci),
    .io_s(FullAdder_841_io_s),
    .io_co(FullAdder_841_io_co)
  );
  FullAdder FullAdder_842 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_842_io_a),
    .io_b(FullAdder_842_io_b),
    .io_ci(FullAdder_842_io_ci),
    .io_s(FullAdder_842_io_s),
    .io_co(FullAdder_842_io_co)
  );
  FullAdder FullAdder_843 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_843_io_a),
    .io_b(FullAdder_843_io_b),
    .io_ci(FullAdder_843_io_ci),
    .io_s(FullAdder_843_io_s),
    .io_co(FullAdder_843_io_co)
  );
  FullAdder FullAdder_844 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_844_io_a),
    .io_b(FullAdder_844_io_b),
    .io_ci(FullAdder_844_io_ci),
    .io_s(FullAdder_844_io_s),
    .io_co(FullAdder_844_io_co)
  );
  FullAdder FullAdder_845 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_845_io_a),
    .io_b(FullAdder_845_io_b),
    .io_ci(FullAdder_845_io_ci),
    .io_s(FullAdder_845_io_s),
    .io_co(FullAdder_845_io_co)
  );
  FullAdder FullAdder_846 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_846_io_a),
    .io_b(FullAdder_846_io_b),
    .io_ci(FullAdder_846_io_ci),
    .io_s(FullAdder_846_io_s),
    .io_co(FullAdder_846_io_co)
  );
  FullAdder FullAdder_847 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_847_io_a),
    .io_b(FullAdder_847_io_b),
    .io_ci(FullAdder_847_io_ci),
    .io_s(FullAdder_847_io_s),
    .io_co(FullAdder_847_io_co)
  );
  FullAdder FullAdder_848 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_848_io_a),
    .io_b(FullAdder_848_io_b),
    .io_ci(FullAdder_848_io_ci),
    .io_s(FullAdder_848_io_s),
    .io_co(FullAdder_848_io_co)
  );
  FullAdder FullAdder_849 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_849_io_a),
    .io_b(FullAdder_849_io_b),
    .io_ci(FullAdder_849_io_ci),
    .io_s(FullAdder_849_io_s),
    .io_co(FullAdder_849_io_co)
  );
  FullAdder FullAdder_850 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_850_io_a),
    .io_b(FullAdder_850_io_b),
    .io_ci(FullAdder_850_io_ci),
    .io_s(FullAdder_850_io_s),
    .io_co(FullAdder_850_io_co)
  );
  FullAdder FullAdder_851 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_851_io_a),
    .io_b(FullAdder_851_io_b),
    .io_ci(FullAdder_851_io_ci),
    .io_s(FullAdder_851_io_s),
    .io_co(FullAdder_851_io_co)
  );
  FullAdder FullAdder_852 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_852_io_a),
    .io_b(FullAdder_852_io_b),
    .io_ci(FullAdder_852_io_ci),
    .io_s(FullAdder_852_io_s),
    .io_co(FullAdder_852_io_co)
  );
  FullAdder FullAdder_853 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_853_io_a),
    .io_b(FullAdder_853_io_b),
    .io_ci(FullAdder_853_io_ci),
    .io_s(FullAdder_853_io_s),
    .io_co(FullAdder_853_io_co)
  );
  FullAdder FullAdder_854 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_854_io_a),
    .io_b(FullAdder_854_io_b),
    .io_ci(FullAdder_854_io_ci),
    .io_s(FullAdder_854_io_s),
    .io_co(FullAdder_854_io_co)
  );
  FullAdder FullAdder_855 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_855_io_a),
    .io_b(FullAdder_855_io_b),
    .io_ci(FullAdder_855_io_ci),
    .io_s(FullAdder_855_io_s),
    .io_co(FullAdder_855_io_co)
  );
  FullAdder FullAdder_856 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_856_io_a),
    .io_b(FullAdder_856_io_b),
    .io_ci(FullAdder_856_io_ci),
    .io_s(FullAdder_856_io_s),
    .io_co(FullAdder_856_io_co)
  );
  FullAdder FullAdder_857 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_857_io_a),
    .io_b(FullAdder_857_io_b),
    .io_ci(FullAdder_857_io_ci),
    .io_s(FullAdder_857_io_s),
    .io_co(FullAdder_857_io_co)
  );
  FullAdder FullAdder_858 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_858_io_a),
    .io_b(FullAdder_858_io_b),
    .io_ci(FullAdder_858_io_ci),
    .io_s(FullAdder_858_io_s),
    .io_co(FullAdder_858_io_co)
  );
  FullAdder FullAdder_859 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_859_io_a),
    .io_b(FullAdder_859_io_b),
    .io_ci(FullAdder_859_io_ci),
    .io_s(FullAdder_859_io_s),
    .io_co(FullAdder_859_io_co)
  );
  FullAdder FullAdder_860 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_860_io_a),
    .io_b(FullAdder_860_io_b),
    .io_ci(FullAdder_860_io_ci),
    .io_s(FullAdder_860_io_s),
    .io_co(FullAdder_860_io_co)
  );
  FullAdder FullAdder_861 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_861_io_a),
    .io_b(FullAdder_861_io_b),
    .io_ci(FullAdder_861_io_ci),
    .io_s(FullAdder_861_io_s),
    .io_co(FullAdder_861_io_co)
  );
  FullAdder FullAdder_862 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_862_io_a),
    .io_b(FullAdder_862_io_b),
    .io_ci(FullAdder_862_io_ci),
    .io_s(FullAdder_862_io_s),
    .io_co(FullAdder_862_io_co)
  );
  FullAdder FullAdder_863 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_863_io_a),
    .io_b(FullAdder_863_io_b),
    .io_ci(FullAdder_863_io_ci),
    .io_s(FullAdder_863_io_s),
    .io_co(FullAdder_863_io_co)
  );
  FullAdder FullAdder_864 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_864_io_a),
    .io_b(FullAdder_864_io_b),
    .io_ci(FullAdder_864_io_ci),
    .io_s(FullAdder_864_io_s),
    .io_co(FullAdder_864_io_co)
  );
  FullAdder FullAdder_865 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_865_io_a),
    .io_b(FullAdder_865_io_b),
    .io_ci(FullAdder_865_io_ci),
    .io_s(FullAdder_865_io_s),
    .io_co(FullAdder_865_io_co)
  );
  FullAdder FullAdder_866 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_866_io_a),
    .io_b(FullAdder_866_io_b),
    .io_ci(FullAdder_866_io_ci),
    .io_s(FullAdder_866_io_s),
    .io_co(FullAdder_866_io_co)
  );
  FullAdder FullAdder_867 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_867_io_a),
    .io_b(FullAdder_867_io_b),
    .io_ci(FullAdder_867_io_ci),
    .io_s(FullAdder_867_io_s),
    .io_co(FullAdder_867_io_co)
  );
  FullAdder FullAdder_868 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_868_io_a),
    .io_b(FullAdder_868_io_b),
    .io_ci(FullAdder_868_io_ci),
    .io_s(FullAdder_868_io_s),
    .io_co(FullAdder_868_io_co)
  );
  FullAdder FullAdder_869 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_869_io_a),
    .io_b(FullAdder_869_io_b),
    .io_ci(FullAdder_869_io_ci),
    .io_s(FullAdder_869_io_s),
    .io_co(FullAdder_869_io_co)
  );
  FullAdder FullAdder_870 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_870_io_a),
    .io_b(FullAdder_870_io_b),
    .io_ci(FullAdder_870_io_ci),
    .io_s(FullAdder_870_io_s),
    .io_co(FullAdder_870_io_co)
  );
  FullAdder FullAdder_871 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_871_io_a),
    .io_b(FullAdder_871_io_b),
    .io_ci(FullAdder_871_io_ci),
    .io_s(FullAdder_871_io_s),
    .io_co(FullAdder_871_io_co)
  );
  FullAdder FullAdder_872 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_872_io_a),
    .io_b(FullAdder_872_io_b),
    .io_ci(FullAdder_872_io_ci),
    .io_s(FullAdder_872_io_s),
    .io_co(FullAdder_872_io_co)
  );
  FullAdder FullAdder_873 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_873_io_a),
    .io_b(FullAdder_873_io_b),
    .io_ci(FullAdder_873_io_ci),
    .io_s(FullAdder_873_io_s),
    .io_co(FullAdder_873_io_co)
  );
  FullAdder FullAdder_874 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_874_io_a),
    .io_b(FullAdder_874_io_b),
    .io_ci(FullAdder_874_io_ci),
    .io_s(FullAdder_874_io_s),
    .io_co(FullAdder_874_io_co)
  );
  FullAdder FullAdder_875 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_875_io_a),
    .io_b(FullAdder_875_io_b),
    .io_ci(FullAdder_875_io_ci),
    .io_s(FullAdder_875_io_s),
    .io_co(FullAdder_875_io_co)
  );
  FullAdder FullAdder_876 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_876_io_a),
    .io_b(FullAdder_876_io_b),
    .io_ci(FullAdder_876_io_ci),
    .io_s(FullAdder_876_io_s),
    .io_co(FullAdder_876_io_co)
  );
  FullAdder FullAdder_877 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_877_io_a),
    .io_b(FullAdder_877_io_b),
    .io_ci(FullAdder_877_io_ci),
    .io_s(FullAdder_877_io_s),
    .io_co(FullAdder_877_io_co)
  );
  FullAdder FullAdder_878 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_878_io_a),
    .io_b(FullAdder_878_io_b),
    .io_ci(FullAdder_878_io_ci),
    .io_s(FullAdder_878_io_s),
    .io_co(FullAdder_878_io_co)
  );
  FullAdder FullAdder_879 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_879_io_a),
    .io_b(FullAdder_879_io_b),
    .io_ci(FullAdder_879_io_ci),
    .io_s(FullAdder_879_io_s),
    .io_co(FullAdder_879_io_co)
  );
  FullAdder FullAdder_880 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_880_io_a),
    .io_b(FullAdder_880_io_b),
    .io_ci(FullAdder_880_io_ci),
    .io_s(FullAdder_880_io_s),
    .io_co(FullAdder_880_io_co)
  );
  HalfAdder HalfAdder_20 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_20_io_a),
    .io_b(HalfAdder_20_io_b),
    .io_s(HalfAdder_20_io_s),
    .io_co(HalfAdder_20_io_co)
  );
  FullAdder FullAdder_881 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_881_io_a),
    .io_b(FullAdder_881_io_b),
    .io_ci(FullAdder_881_io_ci),
    .io_s(FullAdder_881_io_s),
    .io_co(FullAdder_881_io_co)
  );
  FullAdder FullAdder_882 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_882_io_a),
    .io_b(FullAdder_882_io_b),
    .io_ci(FullAdder_882_io_ci),
    .io_s(FullAdder_882_io_s),
    .io_co(FullAdder_882_io_co)
  );
  FullAdder FullAdder_883 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_883_io_a),
    .io_b(FullAdder_883_io_b),
    .io_ci(FullAdder_883_io_ci),
    .io_s(FullAdder_883_io_s),
    .io_co(FullAdder_883_io_co)
  );
  FullAdder FullAdder_884 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_884_io_a),
    .io_b(FullAdder_884_io_b),
    .io_ci(FullAdder_884_io_ci),
    .io_s(FullAdder_884_io_s),
    .io_co(FullAdder_884_io_co)
  );
  FullAdder FullAdder_885 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_885_io_a),
    .io_b(FullAdder_885_io_b),
    .io_ci(FullAdder_885_io_ci),
    .io_s(FullAdder_885_io_s),
    .io_co(FullAdder_885_io_co)
  );
  FullAdder FullAdder_886 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_886_io_a),
    .io_b(FullAdder_886_io_b),
    .io_ci(FullAdder_886_io_ci),
    .io_s(FullAdder_886_io_s),
    .io_co(FullAdder_886_io_co)
  );
  FullAdder FullAdder_887 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_887_io_a),
    .io_b(FullAdder_887_io_b),
    .io_ci(FullAdder_887_io_ci),
    .io_s(FullAdder_887_io_s),
    .io_co(FullAdder_887_io_co)
  );
  FullAdder FullAdder_888 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_888_io_a),
    .io_b(FullAdder_888_io_b),
    .io_ci(FullAdder_888_io_ci),
    .io_s(FullAdder_888_io_s),
    .io_co(FullAdder_888_io_co)
  );
  FullAdder FullAdder_889 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_889_io_a),
    .io_b(FullAdder_889_io_b),
    .io_ci(FullAdder_889_io_ci),
    .io_s(FullAdder_889_io_s),
    .io_co(FullAdder_889_io_co)
  );
  FullAdder FullAdder_890 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_890_io_a),
    .io_b(FullAdder_890_io_b),
    .io_ci(FullAdder_890_io_ci),
    .io_s(FullAdder_890_io_s),
    .io_co(FullAdder_890_io_co)
  );
  FullAdder FullAdder_891 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_891_io_a),
    .io_b(FullAdder_891_io_b),
    .io_ci(FullAdder_891_io_ci),
    .io_s(FullAdder_891_io_s),
    .io_co(FullAdder_891_io_co)
  );
  FullAdder FullAdder_892 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_892_io_a),
    .io_b(FullAdder_892_io_b),
    .io_ci(FullAdder_892_io_ci),
    .io_s(FullAdder_892_io_s),
    .io_co(FullAdder_892_io_co)
  );
  FullAdder FullAdder_893 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_893_io_a),
    .io_b(FullAdder_893_io_b),
    .io_ci(FullAdder_893_io_ci),
    .io_s(FullAdder_893_io_s),
    .io_co(FullAdder_893_io_co)
  );
  FullAdder FullAdder_894 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_894_io_a),
    .io_b(FullAdder_894_io_b),
    .io_ci(FullAdder_894_io_ci),
    .io_s(FullAdder_894_io_s),
    .io_co(FullAdder_894_io_co)
  );
  FullAdder FullAdder_895 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_895_io_a),
    .io_b(FullAdder_895_io_b),
    .io_ci(FullAdder_895_io_ci),
    .io_s(FullAdder_895_io_s),
    .io_co(FullAdder_895_io_co)
  );
  FullAdder FullAdder_896 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_896_io_a),
    .io_b(FullAdder_896_io_b),
    .io_ci(FullAdder_896_io_ci),
    .io_s(FullAdder_896_io_s),
    .io_co(FullAdder_896_io_co)
  );
  FullAdder FullAdder_897 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_897_io_a),
    .io_b(FullAdder_897_io_b),
    .io_ci(FullAdder_897_io_ci),
    .io_s(FullAdder_897_io_s),
    .io_co(FullAdder_897_io_co)
  );
  FullAdder FullAdder_898 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_898_io_a),
    .io_b(FullAdder_898_io_b),
    .io_ci(FullAdder_898_io_ci),
    .io_s(FullAdder_898_io_s),
    .io_co(FullAdder_898_io_co)
  );
  FullAdder FullAdder_899 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_899_io_a),
    .io_b(FullAdder_899_io_b),
    .io_ci(FullAdder_899_io_ci),
    .io_s(FullAdder_899_io_s),
    .io_co(FullAdder_899_io_co)
  );
  FullAdder FullAdder_900 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_900_io_a),
    .io_b(FullAdder_900_io_b),
    .io_ci(FullAdder_900_io_ci),
    .io_s(FullAdder_900_io_s),
    .io_co(FullAdder_900_io_co)
  );
  FullAdder FullAdder_901 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_901_io_a),
    .io_b(FullAdder_901_io_b),
    .io_ci(FullAdder_901_io_ci),
    .io_s(FullAdder_901_io_s),
    .io_co(FullAdder_901_io_co)
  );
  FullAdder FullAdder_902 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_902_io_a),
    .io_b(FullAdder_902_io_b),
    .io_ci(FullAdder_902_io_ci),
    .io_s(FullAdder_902_io_s),
    .io_co(FullAdder_902_io_co)
  );
  FullAdder FullAdder_903 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_903_io_a),
    .io_b(FullAdder_903_io_b),
    .io_ci(FullAdder_903_io_ci),
    .io_s(FullAdder_903_io_s),
    .io_co(FullAdder_903_io_co)
  );
  FullAdder FullAdder_904 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_904_io_a),
    .io_b(FullAdder_904_io_b),
    .io_ci(FullAdder_904_io_ci),
    .io_s(FullAdder_904_io_s),
    .io_co(FullAdder_904_io_co)
  );
  FullAdder FullAdder_905 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_905_io_a),
    .io_b(FullAdder_905_io_b),
    .io_ci(FullAdder_905_io_ci),
    .io_s(FullAdder_905_io_s),
    .io_co(FullAdder_905_io_co)
  );
  FullAdder FullAdder_906 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_906_io_a),
    .io_b(FullAdder_906_io_b),
    .io_ci(FullAdder_906_io_ci),
    .io_s(FullAdder_906_io_s),
    .io_co(FullAdder_906_io_co)
  );
  FullAdder FullAdder_907 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_907_io_a),
    .io_b(FullAdder_907_io_b),
    .io_ci(FullAdder_907_io_ci),
    .io_s(FullAdder_907_io_s),
    .io_co(FullAdder_907_io_co)
  );
  FullAdder FullAdder_908 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_908_io_a),
    .io_b(FullAdder_908_io_b),
    .io_ci(FullAdder_908_io_ci),
    .io_s(FullAdder_908_io_s),
    .io_co(FullAdder_908_io_co)
  );
  FullAdder FullAdder_909 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_909_io_a),
    .io_b(FullAdder_909_io_b),
    .io_ci(FullAdder_909_io_ci),
    .io_s(FullAdder_909_io_s),
    .io_co(FullAdder_909_io_co)
  );
  FullAdder FullAdder_910 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_910_io_a),
    .io_b(FullAdder_910_io_b),
    .io_ci(FullAdder_910_io_ci),
    .io_s(FullAdder_910_io_s),
    .io_co(FullAdder_910_io_co)
  );
  FullAdder FullAdder_911 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_911_io_a),
    .io_b(FullAdder_911_io_b),
    .io_ci(FullAdder_911_io_ci),
    .io_s(FullAdder_911_io_s),
    .io_co(FullAdder_911_io_co)
  );
  FullAdder FullAdder_912 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_912_io_a),
    .io_b(FullAdder_912_io_b),
    .io_ci(FullAdder_912_io_ci),
    .io_s(FullAdder_912_io_s),
    .io_co(FullAdder_912_io_co)
  );
  FullAdder FullAdder_913 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_913_io_a),
    .io_b(FullAdder_913_io_b),
    .io_ci(FullAdder_913_io_ci),
    .io_s(FullAdder_913_io_s),
    .io_co(FullAdder_913_io_co)
  );
  FullAdder FullAdder_914 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_914_io_a),
    .io_b(FullAdder_914_io_b),
    .io_ci(FullAdder_914_io_ci),
    .io_s(FullAdder_914_io_s),
    .io_co(FullAdder_914_io_co)
  );
  FullAdder FullAdder_915 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_915_io_a),
    .io_b(FullAdder_915_io_b),
    .io_ci(FullAdder_915_io_ci),
    .io_s(FullAdder_915_io_s),
    .io_co(FullAdder_915_io_co)
  );
  FullAdder FullAdder_916 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_916_io_a),
    .io_b(FullAdder_916_io_b),
    .io_ci(FullAdder_916_io_ci),
    .io_s(FullAdder_916_io_s),
    .io_co(FullAdder_916_io_co)
  );
  FullAdder FullAdder_917 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_917_io_a),
    .io_b(FullAdder_917_io_b),
    .io_ci(FullAdder_917_io_ci),
    .io_s(FullAdder_917_io_s),
    .io_co(FullAdder_917_io_co)
  );
  FullAdder FullAdder_918 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_918_io_a),
    .io_b(FullAdder_918_io_b),
    .io_ci(FullAdder_918_io_ci),
    .io_s(FullAdder_918_io_s),
    .io_co(FullAdder_918_io_co)
  );
  FullAdder FullAdder_919 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_919_io_a),
    .io_b(FullAdder_919_io_b),
    .io_ci(FullAdder_919_io_ci),
    .io_s(FullAdder_919_io_s),
    .io_co(FullAdder_919_io_co)
  );
  FullAdder FullAdder_920 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_920_io_a),
    .io_b(FullAdder_920_io_b),
    .io_ci(FullAdder_920_io_ci),
    .io_s(FullAdder_920_io_s),
    .io_co(FullAdder_920_io_co)
  );
  FullAdder FullAdder_921 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_921_io_a),
    .io_b(FullAdder_921_io_b),
    .io_ci(FullAdder_921_io_ci),
    .io_s(FullAdder_921_io_s),
    .io_co(FullAdder_921_io_co)
  );
  FullAdder FullAdder_922 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_922_io_a),
    .io_b(FullAdder_922_io_b),
    .io_ci(FullAdder_922_io_ci),
    .io_s(FullAdder_922_io_s),
    .io_co(FullAdder_922_io_co)
  );
  FullAdder FullAdder_923 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_923_io_a),
    .io_b(FullAdder_923_io_b),
    .io_ci(FullAdder_923_io_ci),
    .io_s(FullAdder_923_io_s),
    .io_co(FullAdder_923_io_co)
  );
  FullAdder FullAdder_924 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_924_io_a),
    .io_b(FullAdder_924_io_b),
    .io_ci(FullAdder_924_io_ci),
    .io_s(FullAdder_924_io_s),
    .io_co(FullAdder_924_io_co)
  );
  FullAdder FullAdder_925 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_925_io_a),
    .io_b(FullAdder_925_io_b),
    .io_ci(FullAdder_925_io_ci),
    .io_s(FullAdder_925_io_s),
    .io_co(FullAdder_925_io_co)
  );
  FullAdder FullAdder_926 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_926_io_a),
    .io_b(FullAdder_926_io_b),
    .io_ci(FullAdder_926_io_ci),
    .io_s(FullAdder_926_io_s),
    .io_co(FullAdder_926_io_co)
  );
  FullAdder FullAdder_927 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_927_io_a),
    .io_b(FullAdder_927_io_b),
    .io_ci(FullAdder_927_io_ci),
    .io_s(FullAdder_927_io_s),
    .io_co(FullAdder_927_io_co)
  );
  FullAdder FullAdder_928 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_928_io_a),
    .io_b(FullAdder_928_io_b),
    .io_ci(FullAdder_928_io_ci),
    .io_s(FullAdder_928_io_s),
    .io_co(FullAdder_928_io_co)
  );
  FullAdder FullAdder_929 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_929_io_a),
    .io_b(FullAdder_929_io_b),
    .io_ci(FullAdder_929_io_ci),
    .io_s(FullAdder_929_io_s),
    .io_co(FullAdder_929_io_co)
  );
  FullAdder FullAdder_930 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_930_io_a),
    .io_b(FullAdder_930_io_b),
    .io_ci(FullAdder_930_io_ci),
    .io_s(FullAdder_930_io_s),
    .io_co(FullAdder_930_io_co)
  );
  FullAdder FullAdder_931 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_931_io_a),
    .io_b(FullAdder_931_io_b),
    .io_ci(FullAdder_931_io_ci),
    .io_s(FullAdder_931_io_s),
    .io_co(FullAdder_931_io_co)
  );
  FullAdder FullAdder_932 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_932_io_a),
    .io_b(FullAdder_932_io_b),
    .io_ci(FullAdder_932_io_ci),
    .io_s(FullAdder_932_io_s),
    .io_co(FullAdder_932_io_co)
  );
  FullAdder FullAdder_933 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_933_io_a),
    .io_b(FullAdder_933_io_b),
    .io_ci(FullAdder_933_io_ci),
    .io_s(FullAdder_933_io_s),
    .io_co(FullAdder_933_io_co)
  );
  FullAdder FullAdder_934 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_934_io_a),
    .io_b(FullAdder_934_io_b),
    .io_ci(FullAdder_934_io_ci),
    .io_s(FullAdder_934_io_s),
    .io_co(FullAdder_934_io_co)
  );
  FullAdder FullAdder_935 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_935_io_a),
    .io_b(FullAdder_935_io_b),
    .io_ci(FullAdder_935_io_ci),
    .io_s(FullAdder_935_io_s),
    .io_co(FullAdder_935_io_co)
  );
  FullAdder FullAdder_936 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_936_io_a),
    .io_b(FullAdder_936_io_b),
    .io_ci(FullAdder_936_io_ci),
    .io_s(FullAdder_936_io_s),
    .io_co(FullAdder_936_io_co)
  );
  FullAdder FullAdder_937 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_937_io_a),
    .io_b(FullAdder_937_io_b),
    .io_ci(FullAdder_937_io_ci),
    .io_s(FullAdder_937_io_s),
    .io_co(FullAdder_937_io_co)
  );
  FullAdder FullAdder_938 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_938_io_a),
    .io_b(FullAdder_938_io_b),
    .io_ci(FullAdder_938_io_ci),
    .io_s(FullAdder_938_io_s),
    .io_co(FullAdder_938_io_co)
  );
  FullAdder FullAdder_939 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_939_io_a),
    .io_b(FullAdder_939_io_b),
    .io_ci(FullAdder_939_io_ci),
    .io_s(FullAdder_939_io_s),
    .io_co(FullAdder_939_io_co)
  );
  FullAdder FullAdder_940 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_940_io_a),
    .io_b(FullAdder_940_io_b),
    .io_ci(FullAdder_940_io_ci),
    .io_s(FullAdder_940_io_s),
    .io_co(FullAdder_940_io_co)
  );
  FullAdder FullAdder_941 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_941_io_a),
    .io_b(FullAdder_941_io_b),
    .io_ci(FullAdder_941_io_ci),
    .io_s(FullAdder_941_io_s),
    .io_co(FullAdder_941_io_co)
  );
  FullAdder FullAdder_942 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_942_io_a),
    .io_b(FullAdder_942_io_b),
    .io_ci(FullAdder_942_io_ci),
    .io_s(FullAdder_942_io_s),
    .io_co(FullAdder_942_io_co)
  );
  FullAdder FullAdder_943 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_943_io_a),
    .io_b(FullAdder_943_io_b),
    .io_ci(FullAdder_943_io_ci),
    .io_s(FullAdder_943_io_s),
    .io_co(FullAdder_943_io_co)
  );
  FullAdder FullAdder_944 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_944_io_a),
    .io_b(FullAdder_944_io_b),
    .io_ci(FullAdder_944_io_ci),
    .io_s(FullAdder_944_io_s),
    .io_co(FullAdder_944_io_co)
  );
  FullAdder FullAdder_945 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_945_io_a),
    .io_b(FullAdder_945_io_b),
    .io_ci(FullAdder_945_io_ci),
    .io_s(FullAdder_945_io_s),
    .io_co(FullAdder_945_io_co)
  );
  FullAdder FullAdder_946 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_946_io_a),
    .io_b(FullAdder_946_io_b),
    .io_ci(FullAdder_946_io_ci),
    .io_s(FullAdder_946_io_s),
    .io_co(FullAdder_946_io_co)
  );
  FullAdder FullAdder_947 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_947_io_a),
    .io_b(FullAdder_947_io_b),
    .io_ci(FullAdder_947_io_ci),
    .io_s(FullAdder_947_io_s),
    .io_co(FullAdder_947_io_co)
  );
  FullAdder FullAdder_948 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_948_io_a),
    .io_b(FullAdder_948_io_b),
    .io_ci(FullAdder_948_io_ci),
    .io_s(FullAdder_948_io_s),
    .io_co(FullAdder_948_io_co)
  );
  FullAdder FullAdder_949 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_949_io_a),
    .io_b(FullAdder_949_io_b),
    .io_ci(FullAdder_949_io_ci),
    .io_s(FullAdder_949_io_s),
    .io_co(FullAdder_949_io_co)
  );
  FullAdder FullAdder_950 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_950_io_a),
    .io_b(FullAdder_950_io_b),
    .io_ci(FullAdder_950_io_ci),
    .io_s(FullAdder_950_io_s),
    .io_co(FullAdder_950_io_co)
  );
  FullAdder FullAdder_951 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_951_io_a),
    .io_b(FullAdder_951_io_b),
    .io_ci(FullAdder_951_io_ci),
    .io_s(FullAdder_951_io_s),
    .io_co(FullAdder_951_io_co)
  );
  FullAdder FullAdder_952 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_952_io_a),
    .io_b(FullAdder_952_io_b),
    .io_ci(FullAdder_952_io_ci),
    .io_s(FullAdder_952_io_s),
    .io_co(FullAdder_952_io_co)
  );
  FullAdder FullAdder_953 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_953_io_a),
    .io_b(FullAdder_953_io_b),
    .io_ci(FullAdder_953_io_ci),
    .io_s(FullAdder_953_io_s),
    .io_co(FullAdder_953_io_co)
  );
  FullAdder FullAdder_954 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_954_io_a),
    .io_b(FullAdder_954_io_b),
    .io_ci(FullAdder_954_io_ci),
    .io_s(FullAdder_954_io_s),
    .io_co(FullAdder_954_io_co)
  );
  FullAdder FullAdder_955 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_955_io_a),
    .io_b(FullAdder_955_io_b),
    .io_ci(FullAdder_955_io_ci),
    .io_s(FullAdder_955_io_s),
    .io_co(FullAdder_955_io_co)
  );
  FullAdder FullAdder_956 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_956_io_a),
    .io_b(FullAdder_956_io_b),
    .io_ci(FullAdder_956_io_ci),
    .io_s(FullAdder_956_io_s),
    .io_co(FullAdder_956_io_co)
  );
  FullAdder FullAdder_957 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_957_io_a),
    .io_b(FullAdder_957_io_b),
    .io_ci(FullAdder_957_io_ci),
    .io_s(FullAdder_957_io_s),
    .io_co(FullAdder_957_io_co)
  );
  FullAdder FullAdder_958 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_958_io_a),
    .io_b(FullAdder_958_io_b),
    .io_ci(FullAdder_958_io_ci),
    .io_s(FullAdder_958_io_s),
    .io_co(FullAdder_958_io_co)
  );
  FullAdder FullAdder_959 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_959_io_a),
    .io_b(FullAdder_959_io_b),
    .io_ci(FullAdder_959_io_ci),
    .io_s(FullAdder_959_io_s),
    .io_co(FullAdder_959_io_co)
  );
  FullAdder FullAdder_960 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_960_io_a),
    .io_b(FullAdder_960_io_b),
    .io_ci(FullAdder_960_io_ci),
    .io_s(FullAdder_960_io_s),
    .io_co(FullAdder_960_io_co)
  );
  FullAdder FullAdder_961 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_961_io_a),
    .io_b(FullAdder_961_io_b),
    .io_ci(FullAdder_961_io_ci),
    .io_s(FullAdder_961_io_s),
    .io_co(FullAdder_961_io_co)
  );
  FullAdder FullAdder_962 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_962_io_a),
    .io_b(FullAdder_962_io_b),
    .io_ci(FullAdder_962_io_ci),
    .io_s(FullAdder_962_io_s),
    .io_co(FullAdder_962_io_co)
  );
  FullAdder FullAdder_963 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_963_io_a),
    .io_b(FullAdder_963_io_b),
    .io_ci(FullAdder_963_io_ci),
    .io_s(FullAdder_963_io_s),
    .io_co(FullAdder_963_io_co)
  );
  FullAdder FullAdder_964 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_964_io_a),
    .io_b(FullAdder_964_io_b),
    .io_ci(FullAdder_964_io_ci),
    .io_s(FullAdder_964_io_s),
    .io_co(FullAdder_964_io_co)
  );
  FullAdder FullAdder_965 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_965_io_a),
    .io_b(FullAdder_965_io_b),
    .io_ci(FullAdder_965_io_ci),
    .io_s(FullAdder_965_io_s),
    .io_co(FullAdder_965_io_co)
  );
  FullAdder FullAdder_966 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_966_io_a),
    .io_b(FullAdder_966_io_b),
    .io_ci(FullAdder_966_io_ci),
    .io_s(FullAdder_966_io_s),
    .io_co(FullAdder_966_io_co)
  );
  FullAdder FullAdder_967 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_967_io_a),
    .io_b(FullAdder_967_io_b),
    .io_ci(FullAdder_967_io_ci),
    .io_s(FullAdder_967_io_s),
    .io_co(FullAdder_967_io_co)
  );
  FullAdder FullAdder_968 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_968_io_a),
    .io_b(FullAdder_968_io_b),
    .io_ci(FullAdder_968_io_ci),
    .io_s(FullAdder_968_io_s),
    .io_co(FullAdder_968_io_co)
  );
  FullAdder FullAdder_969 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_969_io_a),
    .io_b(FullAdder_969_io_b),
    .io_ci(FullAdder_969_io_ci),
    .io_s(FullAdder_969_io_s),
    .io_co(FullAdder_969_io_co)
  );
  FullAdder FullAdder_970 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_970_io_a),
    .io_b(FullAdder_970_io_b),
    .io_ci(FullAdder_970_io_ci),
    .io_s(FullAdder_970_io_s),
    .io_co(FullAdder_970_io_co)
  );
  FullAdder FullAdder_971 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_971_io_a),
    .io_b(FullAdder_971_io_b),
    .io_ci(FullAdder_971_io_ci),
    .io_s(FullAdder_971_io_s),
    .io_co(FullAdder_971_io_co)
  );
  FullAdder FullAdder_972 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_972_io_a),
    .io_b(FullAdder_972_io_b),
    .io_ci(FullAdder_972_io_ci),
    .io_s(FullAdder_972_io_s),
    .io_co(FullAdder_972_io_co)
  );
  FullAdder FullAdder_973 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_973_io_a),
    .io_b(FullAdder_973_io_b),
    .io_ci(FullAdder_973_io_ci),
    .io_s(FullAdder_973_io_s),
    .io_co(FullAdder_973_io_co)
  );
  FullAdder FullAdder_974 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_974_io_a),
    .io_b(FullAdder_974_io_b),
    .io_ci(FullAdder_974_io_ci),
    .io_s(FullAdder_974_io_s),
    .io_co(FullAdder_974_io_co)
  );
  FullAdder FullAdder_975 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_975_io_a),
    .io_b(FullAdder_975_io_b),
    .io_ci(FullAdder_975_io_ci),
    .io_s(FullAdder_975_io_s),
    .io_co(FullAdder_975_io_co)
  );
  FullAdder FullAdder_976 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_976_io_a),
    .io_b(FullAdder_976_io_b),
    .io_ci(FullAdder_976_io_ci),
    .io_s(FullAdder_976_io_s),
    .io_co(FullAdder_976_io_co)
  );
  FullAdder FullAdder_977 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_977_io_a),
    .io_b(FullAdder_977_io_b),
    .io_ci(FullAdder_977_io_ci),
    .io_s(FullAdder_977_io_s),
    .io_co(FullAdder_977_io_co)
  );
  HalfAdder HalfAdder_21 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_21_io_a),
    .io_b(HalfAdder_21_io_b),
    .io_s(HalfAdder_21_io_s),
    .io_co(HalfAdder_21_io_co)
  );
  FullAdder FullAdder_978 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_978_io_a),
    .io_b(FullAdder_978_io_b),
    .io_ci(FullAdder_978_io_ci),
    .io_s(FullAdder_978_io_s),
    .io_co(FullAdder_978_io_co)
  );
  FullAdder FullAdder_979 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_979_io_a),
    .io_b(FullAdder_979_io_b),
    .io_ci(FullAdder_979_io_ci),
    .io_s(FullAdder_979_io_s),
    .io_co(FullAdder_979_io_co)
  );
  FullAdder FullAdder_980 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_980_io_a),
    .io_b(FullAdder_980_io_b),
    .io_ci(FullAdder_980_io_ci),
    .io_s(FullAdder_980_io_s),
    .io_co(FullAdder_980_io_co)
  );
  FullAdder FullAdder_981 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_981_io_a),
    .io_b(FullAdder_981_io_b),
    .io_ci(FullAdder_981_io_ci),
    .io_s(FullAdder_981_io_s),
    .io_co(FullAdder_981_io_co)
  );
  FullAdder FullAdder_982 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_982_io_a),
    .io_b(FullAdder_982_io_b),
    .io_ci(FullAdder_982_io_ci),
    .io_s(FullAdder_982_io_s),
    .io_co(FullAdder_982_io_co)
  );
  FullAdder FullAdder_983 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_983_io_a),
    .io_b(FullAdder_983_io_b),
    .io_ci(FullAdder_983_io_ci),
    .io_s(FullAdder_983_io_s),
    .io_co(FullAdder_983_io_co)
  );
  FullAdder FullAdder_984 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_984_io_a),
    .io_b(FullAdder_984_io_b),
    .io_ci(FullAdder_984_io_ci),
    .io_s(FullAdder_984_io_s),
    .io_co(FullAdder_984_io_co)
  );
  FullAdder FullAdder_985 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_985_io_a),
    .io_b(FullAdder_985_io_b),
    .io_ci(FullAdder_985_io_ci),
    .io_s(FullAdder_985_io_s),
    .io_co(FullAdder_985_io_co)
  );
  FullAdder FullAdder_986 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_986_io_a),
    .io_b(FullAdder_986_io_b),
    .io_ci(FullAdder_986_io_ci),
    .io_s(FullAdder_986_io_s),
    .io_co(FullAdder_986_io_co)
  );
  FullAdder FullAdder_987 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_987_io_a),
    .io_b(FullAdder_987_io_b),
    .io_ci(FullAdder_987_io_ci),
    .io_s(FullAdder_987_io_s),
    .io_co(FullAdder_987_io_co)
  );
  FullAdder FullAdder_988 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_988_io_a),
    .io_b(FullAdder_988_io_b),
    .io_ci(FullAdder_988_io_ci),
    .io_s(FullAdder_988_io_s),
    .io_co(FullAdder_988_io_co)
  );
  FullAdder FullAdder_989 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_989_io_a),
    .io_b(FullAdder_989_io_b),
    .io_ci(FullAdder_989_io_ci),
    .io_s(FullAdder_989_io_s),
    .io_co(FullAdder_989_io_co)
  );
  FullAdder FullAdder_990 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_990_io_a),
    .io_b(FullAdder_990_io_b),
    .io_ci(FullAdder_990_io_ci),
    .io_s(FullAdder_990_io_s),
    .io_co(FullAdder_990_io_co)
  );
  FullAdder FullAdder_991 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_991_io_a),
    .io_b(FullAdder_991_io_b),
    .io_ci(FullAdder_991_io_ci),
    .io_s(FullAdder_991_io_s),
    .io_co(FullAdder_991_io_co)
  );
  FullAdder FullAdder_992 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_992_io_a),
    .io_b(FullAdder_992_io_b),
    .io_ci(FullAdder_992_io_ci),
    .io_s(FullAdder_992_io_s),
    .io_co(FullAdder_992_io_co)
  );
  FullAdder FullAdder_993 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_993_io_a),
    .io_b(FullAdder_993_io_b),
    .io_ci(FullAdder_993_io_ci),
    .io_s(FullAdder_993_io_s),
    .io_co(FullAdder_993_io_co)
  );
  FullAdder FullAdder_994 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_994_io_a),
    .io_b(FullAdder_994_io_b),
    .io_ci(FullAdder_994_io_ci),
    .io_s(FullAdder_994_io_s),
    .io_co(FullAdder_994_io_co)
  );
  FullAdder FullAdder_995 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_995_io_a),
    .io_b(FullAdder_995_io_b),
    .io_ci(FullAdder_995_io_ci),
    .io_s(FullAdder_995_io_s),
    .io_co(FullAdder_995_io_co)
  );
  FullAdder FullAdder_996 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_996_io_a),
    .io_b(FullAdder_996_io_b),
    .io_ci(FullAdder_996_io_ci),
    .io_s(FullAdder_996_io_s),
    .io_co(FullAdder_996_io_co)
  );
  FullAdder FullAdder_997 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_997_io_a),
    .io_b(FullAdder_997_io_b),
    .io_ci(FullAdder_997_io_ci),
    .io_s(FullAdder_997_io_s),
    .io_co(FullAdder_997_io_co)
  );
  FullAdder FullAdder_998 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_998_io_a),
    .io_b(FullAdder_998_io_b),
    .io_ci(FullAdder_998_io_ci),
    .io_s(FullAdder_998_io_s),
    .io_co(FullAdder_998_io_co)
  );
  FullAdder FullAdder_999 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_999_io_a),
    .io_b(FullAdder_999_io_b),
    .io_ci(FullAdder_999_io_ci),
    .io_s(FullAdder_999_io_s),
    .io_co(FullAdder_999_io_co)
  );
  FullAdder FullAdder_1000 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1000_io_a),
    .io_b(FullAdder_1000_io_b),
    .io_ci(FullAdder_1000_io_ci),
    .io_s(FullAdder_1000_io_s),
    .io_co(FullAdder_1000_io_co)
  );
  FullAdder FullAdder_1001 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1001_io_a),
    .io_b(FullAdder_1001_io_b),
    .io_ci(FullAdder_1001_io_ci),
    .io_s(FullAdder_1001_io_s),
    .io_co(FullAdder_1001_io_co)
  );
  FullAdder FullAdder_1002 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1002_io_a),
    .io_b(FullAdder_1002_io_b),
    .io_ci(FullAdder_1002_io_ci),
    .io_s(FullAdder_1002_io_s),
    .io_co(FullAdder_1002_io_co)
  );
  FullAdder FullAdder_1003 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1003_io_a),
    .io_b(FullAdder_1003_io_b),
    .io_ci(FullAdder_1003_io_ci),
    .io_s(FullAdder_1003_io_s),
    .io_co(FullAdder_1003_io_co)
  );
  FullAdder FullAdder_1004 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1004_io_a),
    .io_b(FullAdder_1004_io_b),
    .io_ci(FullAdder_1004_io_ci),
    .io_s(FullAdder_1004_io_s),
    .io_co(FullAdder_1004_io_co)
  );
  FullAdder FullAdder_1005 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1005_io_a),
    .io_b(FullAdder_1005_io_b),
    .io_ci(FullAdder_1005_io_ci),
    .io_s(FullAdder_1005_io_s),
    .io_co(FullAdder_1005_io_co)
  );
  FullAdder FullAdder_1006 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1006_io_a),
    .io_b(FullAdder_1006_io_b),
    .io_ci(FullAdder_1006_io_ci),
    .io_s(FullAdder_1006_io_s),
    .io_co(FullAdder_1006_io_co)
  );
  FullAdder FullAdder_1007 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1007_io_a),
    .io_b(FullAdder_1007_io_b),
    .io_ci(FullAdder_1007_io_ci),
    .io_s(FullAdder_1007_io_s),
    .io_co(FullAdder_1007_io_co)
  );
  FullAdder FullAdder_1008 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1008_io_a),
    .io_b(FullAdder_1008_io_b),
    .io_ci(FullAdder_1008_io_ci),
    .io_s(FullAdder_1008_io_s),
    .io_co(FullAdder_1008_io_co)
  );
  FullAdder FullAdder_1009 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1009_io_a),
    .io_b(FullAdder_1009_io_b),
    .io_ci(FullAdder_1009_io_ci),
    .io_s(FullAdder_1009_io_s),
    .io_co(FullAdder_1009_io_co)
  );
  FullAdder FullAdder_1010 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1010_io_a),
    .io_b(FullAdder_1010_io_b),
    .io_ci(FullAdder_1010_io_ci),
    .io_s(FullAdder_1010_io_s),
    .io_co(FullAdder_1010_io_co)
  );
  FullAdder FullAdder_1011 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1011_io_a),
    .io_b(FullAdder_1011_io_b),
    .io_ci(FullAdder_1011_io_ci),
    .io_s(FullAdder_1011_io_s),
    .io_co(FullAdder_1011_io_co)
  );
  FullAdder FullAdder_1012 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1012_io_a),
    .io_b(FullAdder_1012_io_b),
    .io_ci(FullAdder_1012_io_ci),
    .io_s(FullAdder_1012_io_s),
    .io_co(FullAdder_1012_io_co)
  );
  FullAdder FullAdder_1013 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1013_io_a),
    .io_b(FullAdder_1013_io_b),
    .io_ci(FullAdder_1013_io_ci),
    .io_s(FullAdder_1013_io_s),
    .io_co(FullAdder_1013_io_co)
  );
  FullAdder FullAdder_1014 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1014_io_a),
    .io_b(FullAdder_1014_io_b),
    .io_ci(FullAdder_1014_io_ci),
    .io_s(FullAdder_1014_io_s),
    .io_co(FullAdder_1014_io_co)
  );
  FullAdder FullAdder_1015 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1015_io_a),
    .io_b(FullAdder_1015_io_b),
    .io_ci(FullAdder_1015_io_ci),
    .io_s(FullAdder_1015_io_s),
    .io_co(FullAdder_1015_io_co)
  );
  FullAdder FullAdder_1016 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1016_io_a),
    .io_b(FullAdder_1016_io_b),
    .io_ci(FullAdder_1016_io_ci),
    .io_s(FullAdder_1016_io_s),
    .io_co(FullAdder_1016_io_co)
  );
  FullAdder FullAdder_1017 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1017_io_a),
    .io_b(FullAdder_1017_io_b),
    .io_ci(FullAdder_1017_io_ci),
    .io_s(FullAdder_1017_io_s),
    .io_co(FullAdder_1017_io_co)
  );
  FullAdder FullAdder_1018 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1018_io_a),
    .io_b(FullAdder_1018_io_b),
    .io_ci(FullAdder_1018_io_ci),
    .io_s(FullAdder_1018_io_s),
    .io_co(FullAdder_1018_io_co)
  );
  FullAdder FullAdder_1019 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1019_io_a),
    .io_b(FullAdder_1019_io_b),
    .io_ci(FullAdder_1019_io_ci),
    .io_s(FullAdder_1019_io_s),
    .io_co(FullAdder_1019_io_co)
  );
  FullAdder FullAdder_1020 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1020_io_a),
    .io_b(FullAdder_1020_io_b),
    .io_ci(FullAdder_1020_io_ci),
    .io_s(FullAdder_1020_io_s),
    .io_co(FullAdder_1020_io_co)
  );
  FullAdder FullAdder_1021 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1021_io_a),
    .io_b(FullAdder_1021_io_b),
    .io_ci(FullAdder_1021_io_ci),
    .io_s(FullAdder_1021_io_s),
    .io_co(FullAdder_1021_io_co)
  );
  FullAdder FullAdder_1022 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1022_io_a),
    .io_b(FullAdder_1022_io_b),
    .io_ci(FullAdder_1022_io_ci),
    .io_s(FullAdder_1022_io_s),
    .io_co(FullAdder_1022_io_co)
  );
  FullAdder FullAdder_1023 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1023_io_a),
    .io_b(FullAdder_1023_io_b),
    .io_ci(FullAdder_1023_io_ci),
    .io_s(FullAdder_1023_io_s),
    .io_co(FullAdder_1023_io_co)
  );
  FullAdder FullAdder_1024 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1024_io_a),
    .io_b(FullAdder_1024_io_b),
    .io_ci(FullAdder_1024_io_ci),
    .io_s(FullAdder_1024_io_s),
    .io_co(FullAdder_1024_io_co)
  );
  FullAdder FullAdder_1025 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1025_io_a),
    .io_b(FullAdder_1025_io_b),
    .io_ci(FullAdder_1025_io_ci),
    .io_s(FullAdder_1025_io_s),
    .io_co(FullAdder_1025_io_co)
  );
  FullAdder FullAdder_1026 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1026_io_a),
    .io_b(FullAdder_1026_io_b),
    .io_ci(FullAdder_1026_io_ci),
    .io_s(FullAdder_1026_io_s),
    .io_co(FullAdder_1026_io_co)
  );
  FullAdder FullAdder_1027 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1027_io_a),
    .io_b(FullAdder_1027_io_b),
    .io_ci(FullAdder_1027_io_ci),
    .io_s(FullAdder_1027_io_s),
    .io_co(FullAdder_1027_io_co)
  );
  FullAdder FullAdder_1028 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1028_io_a),
    .io_b(FullAdder_1028_io_b),
    .io_ci(FullAdder_1028_io_ci),
    .io_s(FullAdder_1028_io_s),
    .io_co(FullAdder_1028_io_co)
  );
  FullAdder FullAdder_1029 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1029_io_a),
    .io_b(FullAdder_1029_io_b),
    .io_ci(FullAdder_1029_io_ci),
    .io_s(FullAdder_1029_io_s),
    .io_co(FullAdder_1029_io_co)
  );
  FullAdder FullAdder_1030 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1030_io_a),
    .io_b(FullAdder_1030_io_b),
    .io_ci(FullAdder_1030_io_ci),
    .io_s(FullAdder_1030_io_s),
    .io_co(FullAdder_1030_io_co)
  );
  FullAdder FullAdder_1031 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1031_io_a),
    .io_b(FullAdder_1031_io_b),
    .io_ci(FullAdder_1031_io_ci),
    .io_s(FullAdder_1031_io_s),
    .io_co(FullAdder_1031_io_co)
  );
  FullAdder FullAdder_1032 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1032_io_a),
    .io_b(FullAdder_1032_io_b),
    .io_ci(FullAdder_1032_io_ci),
    .io_s(FullAdder_1032_io_s),
    .io_co(FullAdder_1032_io_co)
  );
  FullAdder FullAdder_1033 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1033_io_a),
    .io_b(FullAdder_1033_io_b),
    .io_ci(FullAdder_1033_io_ci),
    .io_s(FullAdder_1033_io_s),
    .io_co(FullAdder_1033_io_co)
  );
  FullAdder FullAdder_1034 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1034_io_a),
    .io_b(FullAdder_1034_io_b),
    .io_ci(FullAdder_1034_io_ci),
    .io_s(FullAdder_1034_io_s),
    .io_co(FullAdder_1034_io_co)
  );
  FullAdder FullAdder_1035 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1035_io_a),
    .io_b(FullAdder_1035_io_b),
    .io_ci(FullAdder_1035_io_ci),
    .io_s(FullAdder_1035_io_s),
    .io_co(FullAdder_1035_io_co)
  );
  FullAdder FullAdder_1036 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1036_io_a),
    .io_b(FullAdder_1036_io_b),
    .io_ci(FullAdder_1036_io_ci),
    .io_s(FullAdder_1036_io_s),
    .io_co(FullAdder_1036_io_co)
  );
  FullAdder FullAdder_1037 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1037_io_a),
    .io_b(FullAdder_1037_io_b),
    .io_ci(FullAdder_1037_io_ci),
    .io_s(FullAdder_1037_io_s),
    .io_co(FullAdder_1037_io_co)
  );
  FullAdder FullAdder_1038 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1038_io_a),
    .io_b(FullAdder_1038_io_b),
    .io_ci(FullAdder_1038_io_ci),
    .io_s(FullAdder_1038_io_s),
    .io_co(FullAdder_1038_io_co)
  );
  FullAdder FullAdder_1039 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1039_io_a),
    .io_b(FullAdder_1039_io_b),
    .io_ci(FullAdder_1039_io_ci),
    .io_s(FullAdder_1039_io_s),
    .io_co(FullAdder_1039_io_co)
  );
  FullAdder FullAdder_1040 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1040_io_a),
    .io_b(FullAdder_1040_io_b),
    .io_ci(FullAdder_1040_io_ci),
    .io_s(FullAdder_1040_io_s),
    .io_co(FullAdder_1040_io_co)
  );
  FullAdder FullAdder_1041 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1041_io_a),
    .io_b(FullAdder_1041_io_b),
    .io_ci(FullAdder_1041_io_ci),
    .io_s(FullAdder_1041_io_s),
    .io_co(FullAdder_1041_io_co)
  );
  FullAdder FullAdder_1042 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1042_io_a),
    .io_b(FullAdder_1042_io_b),
    .io_ci(FullAdder_1042_io_ci),
    .io_s(FullAdder_1042_io_s),
    .io_co(FullAdder_1042_io_co)
  );
  FullAdder FullAdder_1043 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1043_io_a),
    .io_b(FullAdder_1043_io_b),
    .io_ci(FullAdder_1043_io_ci),
    .io_s(FullAdder_1043_io_s),
    .io_co(FullAdder_1043_io_co)
  );
  FullAdder FullAdder_1044 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1044_io_a),
    .io_b(FullAdder_1044_io_b),
    .io_ci(FullAdder_1044_io_ci),
    .io_s(FullAdder_1044_io_s),
    .io_co(FullAdder_1044_io_co)
  );
  FullAdder FullAdder_1045 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1045_io_a),
    .io_b(FullAdder_1045_io_b),
    .io_ci(FullAdder_1045_io_ci),
    .io_s(FullAdder_1045_io_s),
    .io_co(FullAdder_1045_io_co)
  );
  FullAdder FullAdder_1046 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1046_io_a),
    .io_b(FullAdder_1046_io_b),
    .io_ci(FullAdder_1046_io_ci),
    .io_s(FullAdder_1046_io_s),
    .io_co(FullAdder_1046_io_co)
  );
  FullAdder FullAdder_1047 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1047_io_a),
    .io_b(FullAdder_1047_io_b),
    .io_ci(FullAdder_1047_io_ci),
    .io_s(FullAdder_1047_io_s),
    .io_co(FullAdder_1047_io_co)
  );
  FullAdder FullAdder_1048 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1048_io_a),
    .io_b(FullAdder_1048_io_b),
    .io_ci(FullAdder_1048_io_ci),
    .io_s(FullAdder_1048_io_s),
    .io_co(FullAdder_1048_io_co)
  );
  FullAdder FullAdder_1049 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1049_io_a),
    .io_b(FullAdder_1049_io_b),
    .io_ci(FullAdder_1049_io_ci),
    .io_s(FullAdder_1049_io_s),
    .io_co(FullAdder_1049_io_co)
  );
  FullAdder FullAdder_1050 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1050_io_a),
    .io_b(FullAdder_1050_io_b),
    .io_ci(FullAdder_1050_io_ci),
    .io_s(FullAdder_1050_io_s),
    .io_co(FullAdder_1050_io_co)
  );
  FullAdder FullAdder_1051 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1051_io_a),
    .io_b(FullAdder_1051_io_b),
    .io_ci(FullAdder_1051_io_ci),
    .io_s(FullAdder_1051_io_s),
    .io_co(FullAdder_1051_io_co)
  );
  FullAdder FullAdder_1052 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1052_io_a),
    .io_b(FullAdder_1052_io_b),
    .io_ci(FullAdder_1052_io_ci),
    .io_s(FullAdder_1052_io_s),
    .io_co(FullAdder_1052_io_co)
  );
  FullAdder FullAdder_1053 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1053_io_a),
    .io_b(FullAdder_1053_io_b),
    .io_ci(FullAdder_1053_io_ci),
    .io_s(FullAdder_1053_io_s),
    .io_co(FullAdder_1053_io_co)
  );
  FullAdder FullAdder_1054 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1054_io_a),
    .io_b(FullAdder_1054_io_b),
    .io_ci(FullAdder_1054_io_ci),
    .io_s(FullAdder_1054_io_s),
    .io_co(FullAdder_1054_io_co)
  );
  FullAdder FullAdder_1055 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1055_io_a),
    .io_b(FullAdder_1055_io_b),
    .io_ci(FullAdder_1055_io_ci),
    .io_s(FullAdder_1055_io_s),
    .io_co(FullAdder_1055_io_co)
  );
  FullAdder FullAdder_1056 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1056_io_a),
    .io_b(FullAdder_1056_io_b),
    .io_ci(FullAdder_1056_io_ci),
    .io_s(FullAdder_1056_io_s),
    .io_co(FullAdder_1056_io_co)
  );
  FullAdder FullAdder_1057 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1057_io_a),
    .io_b(FullAdder_1057_io_b),
    .io_ci(FullAdder_1057_io_ci),
    .io_s(FullAdder_1057_io_s),
    .io_co(FullAdder_1057_io_co)
  );
  FullAdder FullAdder_1058 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1058_io_a),
    .io_b(FullAdder_1058_io_b),
    .io_ci(FullAdder_1058_io_ci),
    .io_s(FullAdder_1058_io_s),
    .io_co(FullAdder_1058_io_co)
  );
  FullAdder FullAdder_1059 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1059_io_a),
    .io_b(FullAdder_1059_io_b),
    .io_ci(FullAdder_1059_io_ci),
    .io_s(FullAdder_1059_io_s),
    .io_co(FullAdder_1059_io_co)
  );
  FullAdder FullAdder_1060 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1060_io_a),
    .io_b(FullAdder_1060_io_b),
    .io_ci(FullAdder_1060_io_ci),
    .io_s(FullAdder_1060_io_s),
    .io_co(FullAdder_1060_io_co)
  );
  FullAdder FullAdder_1061 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1061_io_a),
    .io_b(FullAdder_1061_io_b),
    .io_ci(FullAdder_1061_io_ci),
    .io_s(FullAdder_1061_io_s),
    .io_co(FullAdder_1061_io_co)
  );
  FullAdder FullAdder_1062 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1062_io_a),
    .io_b(FullAdder_1062_io_b),
    .io_ci(FullAdder_1062_io_ci),
    .io_s(FullAdder_1062_io_s),
    .io_co(FullAdder_1062_io_co)
  );
  FullAdder FullAdder_1063 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1063_io_a),
    .io_b(FullAdder_1063_io_b),
    .io_ci(FullAdder_1063_io_ci),
    .io_s(FullAdder_1063_io_s),
    .io_co(FullAdder_1063_io_co)
  );
  FullAdder FullAdder_1064 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1064_io_a),
    .io_b(FullAdder_1064_io_b),
    .io_ci(FullAdder_1064_io_ci),
    .io_s(FullAdder_1064_io_s),
    .io_co(FullAdder_1064_io_co)
  );
  FullAdder FullAdder_1065 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1065_io_a),
    .io_b(FullAdder_1065_io_b),
    .io_ci(FullAdder_1065_io_ci),
    .io_s(FullAdder_1065_io_s),
    .io_co(FullAdder_1065_io_co)
  );
  FullAdder FullAdder_1066 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1066_io_a),
    .io_b(FullAdder_1066_io_b),
    .io_ci(FullAdder_1066_io_ci),
    .io_s(FullAdder_1066_io_s),
    .io_co(FullAdder_1066_io_co)
  );
  FullAdder FullAdder_1067 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1067_io_a),
    .io_b(FullAdder_1067_io_b),
    .io_ci(FullAdder_1067_io_ci),
    .io_s(FullAdder_1067_io_s),
    .io_co(FullAdder_1067_io_co)
  );
  FullAdder FullAdder_1068 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1068_io_a),
    .io_b(FullAdder_1068_io_b),
    .io_ci(FullAdder_1068_io_ci),
    .io_s(FullAdder_1068_io_s),
    .io_co(FullAdder_1068_io_co)
  );
  FullAdder FullAdder_1069 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1069_io_a),
    .io_b(FullAdder_1069_io_b),
    .io_ci(FullAdder_1069_io_ci),
    .io_s(FullAdder_1069_io_s),
    .io_co(FullAdder_1069_io_co)
  );
  FullAdder FullAdder_1070 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1070_io_a),
    .io_b(FullAdder_1070_io_b),
    .io_ci(FullAdder_1070_io_ci),
    .io_s(FullAdder_1070_io_s),
    .io_co(FullAdder_1070_io_co)
  );
  FullAdder FullAdder_1071 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1071_io_a),
    .io_b(FullAdder_1071_io_b),
    .io_ci(FullAdder_1071_io_ci),
    .io_s(FullAdder_1071_io_s),
    .io_co(FullAdder_1071_io_co)
  );
  FullAdder FullAdder_1072 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1072_io_a),
    .io_b(FullAdder_1072_io_b),
    .io_ci(FullAdder_1072_io_ci),
    .io_s(FullAdder_1072_io_s),
    .io_co(FullAdder_1072_io_co)
  );
  FullAdder FullAdder_1073 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1073_io_a),
    .io_b(FullAdder_1073_io_b),
    .io_ci(FullAdder_1073_io_ci),
    .io_s(FullAdder_1073_io_s),
    .io_co(FullAdder_1073_io_co)
  );
  FullAdder FullAdder_1074 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1074_io_a),
    .io_b(FullAdder_1074_io_b),
    .io_ci(FullAdder_1074_io_ci),
    .io_s(FullAdder_1074_io_s),
    .io_co(FullAdder_1074_io_co)
  );
  FullAdder FullAdder_1075 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1075_io_a),
    .io_b(FullAdder_1075_io_b),
    .io_ci(FullAdder_1075_io_ci),
    .io_s(FullAdder_1075_io_s),
    .io_co(FullAdder_1075_io_co)
  );
  FullAdder FullAdder_1076 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1076_io_a),
    .io_b(FullAdder_1076_io_b),
    .io_ci(FullAdder_1076_io_ci),
    .io_s(FullAdder_1076_io_s),
    .io_co(FullAdder_1076_io_co)
  );
  FullAdder FullAdder_1077 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1077_io_a),
    .io_b(FullAdder_1077_io_b),
    .io_ci(FullAdder_1077_io_ci),
    .io_s(FullAdder_1077_io_s),
    .io_co(FullAdder_1077_io_co)
  );
  FullAdder FullAdder_1078 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1078_io_a),
    .io_b(FullAdder_1078_io_b),
    .io_ci(FullAdder_1078_io_ci),
    .io_s(FullAdder_1078_io_s),
    .io_co(FullAdder_1078_io_co)
  );
  FullAdder FullAdder_1079 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1079_io_a),
    .io_b(FullAdder_1079_io_b),
    .io_ci(FullAdder_1079_io_ci),
    .io_s(FullAdder_1079_io_s),
    .io_co(FullAdder_1079_io_co)
  );
  FullAdder FullAdder_1080 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1080_io_a),
    .io_b(FullAdder_1080_io_b),
    .io_ci(FullAdder_1080_io_ci),
    .io_s(FullAdder_1080_io_s),
    .io_co(FullAdder_1080_io_co)
  );
  FullAdder FullAdder_1081 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1081_io_a),
    .io_b(FullAdder_1081_io_b),
    .io_ci(FullAdder_1081_io_ci),
    .io_s(FullAdder_1081_io_s),
    .io_co(FullAdder_1081_io_co)
  );
  FullAdder FullAdder_1082 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1082_io_a),
    .io_b(FullAdder_1082_io_b),
    .io_ci(FullAdder_1082_io_ci),
    .io_s(FullAdder_1082_io_s),
    .io_co(FullAdder_1082_io_co)
  );
  FullAdder FullAdder_1083 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1083_io_a),
    .io_b(FullAdder_1083_io_b),
    .io_ci(FullAdder_1083_io_ci),
    .io_s(FullAdder_1083_io_s),
    .io_co(FullAdder_1083_io_co)
  );
  FullAdder FullAdder_1084 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1084_io_a),
    .io_b(FullAdder_1084_io_b),
    .io_ci(FullAdder_1084_io_ci),
    .io_s(FullAdder_1084_io_s),
    .io_co(FullAdder_1084_io_co)
  );
  FullAdder FullAdder_1085 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1085_io_a),
    .io_b(FullAdder_1085_io_b),
    .io_ci(FullAdder_1085_io_ci),
    .io_s(FullAdder_1085_io_s),
    .io_co(FullAdder_1085_io_co)
  );
  FullAdder FullAdder_1086 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1086_io_a),
    .io_b(FullAdder_1086_io_b),
    .io_ci(FullAdder_1086_io_ci),
    .io_s(FullAdder_1086_io_s),
    .io_co(FullAdder_1086_io_co)
  );
  FullAdder FullAdder_1087 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1087_io_a),
    .io_b(FullAdder_1087_io_b),
    .io_ci(FullAdder_1087_io_ci),
    .io_s(FullAdder_1087_io_s),
    .io_co(FullAdder_1087_io_co)
  );
  FullAdder FullAdder_1088 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1088_io_a),
    .io_b(FullAdder_1088_io_b),
    .io_ci(FullAdder_1088_io_ci),
    .io_s(FullAdder_1088_io_s),
    .io_co(FullAdder_1088_io_co)
  );
  FullAdder FullAdder_1089 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1089_io_a),
    .io_b(FullAdder_1089_io_b),
    .io_ci(FullAdder_1089_io_ci),
    .io_s(FullAdder_1089_io_s),
    .io_co(FullAdder_1089_io_co)
  );
  FullAdder FullAdder_1090 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1090_io_a),
    .io_b(FullAdder_1090_io_b),
    .io_ci(FullAdder_1090_io_ci),
    .io_s(FullAdder_1090_io_s),
    .io_co(FullAdder_1090_io_co)
  );
  FullAdder FullAdder_1091 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1091_io_a),
    .io_b(FullAdder_1091_io_b),
    .io_ci(FullAdder_1091_io_ci),
    .io_s(FullAdder_1091_io_s),
    .io_co(FullAdder_1091_io_co)
  );
  FullAdder FullAdder_1092 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1092_io_a),
    .io_b(FullAdder_1092_io_b),
    .io_ci(FullAdder_1092_io_ci),
    .io_s(FullAdder_1092_io_s),
    .io_co(FullAdder_1092_io_co)
  );
  FullAdder FullAdder_1093 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1093_io_a),
    .io_b(FullAdder_1093_io_b),
    .io_ci(FullAdder_1093_io_ci),
    .io_s(FullAdder_1093_io_s),
    .io_co(FullAdder_1093_io_co)
  );
  FullAdder FullAdder_1094 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1094_io_a),
    .io_b(FullAdder_1094_io_b),
    .io_ci(FullAdder_1094_io_ci),
    .io_s(FullAdder_1094_io_s),
    .io_co(FullAdder_1094_io_co)
  );
  FullAdder FullAdder_1095 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1095_io_a),
    .io_b(FullAdder_1095_io_b),
    .io_ci(FullAdder_1095_io_ci),
    .io_s(FullAdder_1095_io_s),
    .io_co(FullAdder_1095_io_co)
  );
  FullAdder FullAdder_1096 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1096_io_a),
    .io_b(FullAdder_1096_io_b),
    .io_ci(FullAdder_1096_io_ci),
    .io_s(FullAdder_1096_io_s),
    .io_co(FullAdder_1096_io_co)
  );
  FullAdder FullAdder_1097 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1097_io_a),
    .io_b(FullAdder_1097_io_b),
    .io_ci(FullAdder_1097_io_ci),
    .io_s(FullAdder_1097_io_s),
    .io_co(FullAdder_1097_io_co)
  );
  FullAdder FullAdder_1098 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1098_io_a),
    .io_b(FullAdder_1098_io_b),
    .io_ci(FullAdder_1098_io_ci),
    .io_s(FullAdder_1098_io_s),
    .io_co(FullAdder_1098_io_co)
  );
  FullAdder FullAdder_1099 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1099_io_a),
    .io_b(FullAdder_1099_io_b),
    .io_ci(FullAdder_1099_io_ci),
    .io_s(FullAdder_1099_io_s),
    .io_co(FullAdder_1099_io_co)
  );
  FullAdder FullAdder_1100 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1100_io_a),
    .io_b(FullAdder_1100_io_b),
    .io_ci(FullAdder_1100_io_ci),
    .io_s(FullAdder_1100_io_s),
    .io_co(FullAdder_1100_io_co)
  );
  HalfAdder HalfAdder_22 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_22_io_a),
    .io_b(HalfAdder_22_io_b),
    .io_s(HalfAdder_22_io_s),
    .io_co(HalfAdder_22_io_co)
  );
  FullAdder FullAdder_1101 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1101_io_a),
    .io_b(FullAdder_1101_io_b),
    .io_ci(FullAdder_1101_io_ci),
    .io_s(FullAdder_1101_io_s),
    .io_co(FullAdder_1101_io_co)
  );
  FullAdder FullAdder_1102 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1102_io_a),
    .io_b(FullAdder_1102_io_b),
    .io_ci(FullAdder_1102_io_ci),
    .io_s(FullAdder_1102_io_s),
    .io_co(FullAdder_1102_io_co)
  );
  FullAdder FullAdder_1103 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1103_io_a),
    .io_b(FullAdder_1103_io_b),
    .io_ci(FullAdder_1103_io_ci),
    .io_s(FullAdder_1103_io_s),
    .io_co(FullAdder_1103_io_co)
  );
  FullAdder FullAdder_1104 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1104_io_a),
    .io_b(FullAdder_1104_io_b),
    .io_ci(FullAdder_1104_io_ci),
    .io_s(FullAdder_1104_io_s),
    .io_co(FullAdder_1104_io_co)
  );
  FullAdder FullAdder_1105 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1105_io_a),
    .io_b(FullAdder_1105_io_b),
    .io_ci(FullAdder_1105_io_ci),
    .io_s(FullAdder_1105_io_s),
    .io_co(FullAdder_1105_io_co)
  );
  FullAdder FullAdder_1106 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1106_io_a),
    .io_b(FullAdder_1106_io_b),
    .io_ci(FullAdder_1106_io_ci),
    .io_s(FullAdder_1106_io_s),
    .io_co(FullAdder_1106_io_co)
  );
  FullAdder FullAdder_1107 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1107_io_a),
    .io_b(FullAdder_1107_io_b),
    .io_ci(FullAdder_1107_io_ci),
    .io_s(FullAdder_1107_io_s),
    .io_co(FullAdder_1107_io_co)
  );
  FullAdder FullAdder_1108 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1108_io_a),
    .io_b(FullAdder_1108_io_b),
    .io_ci(FullAdder_1108_io_ci),
    .io_s(FullAdder_1108_io_s),
    .io_co(FullAdder_1108_io_co)
  );
  FullAdder FullAdder_1109 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1109_io_a),
    .io_b(FullAdder_1109_io_b),
    .io_ci(FullAdder_1109_io_ci),
    .io_s(FullAdder_1109_io_s),
    .io_co(FullAdder_1109_io_co)
  );
  FullAdder FullAdder_1110 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1110_io_a),
    .io_b(FullAdder_1110_io_b),
    .io_ci(FullAdder_1110_io_ci),
    .io_s(FullAdder_1110_io_s),
    .io_co(FullAdder_1110_io_co)
  );
  FullAdder FullAdder_1111 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1111_io_a),
    .io_b(FullAdder_1111_io_b),
    .io_ci(FullAdder_1111_io_ci),
    .io_s(FullAdder_1111_io_s),
    .io_co(FullAdder_1111_io_co)
  );
  FullAdder FullAdder_1112 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1112_io_a),
    .io_b(FullAdder_1112_io_b),
    .io_ci(FullAdder_1112_io_ci),
    .io_s(FullAdder_1112_io_s),
    .io_co(FullAdder_1112_io_co)
  );
  FullAdder FullAdder_1113 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1113_io_a),
    .io_b(FullAdder_1113_io_b),
    .io_ci(FullAdder_1113_io_ci),
    .io_s(FullAdder_1113_io_s),
    .io_co(FullAdder_1113_io_co)
  );
  FullAdder FullAdder_1114 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1114_io_a),
    .io_b(FullAdder_1114_io_b),
    .io_ci(FullAdder_1114_io_ci),
    .io_s(FullAdder_1114_io_s),
    .io_co(FullAdder_1114_io_co)
  );
  FullAdder FullAdder_1115 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1115_io_a),
    .io_b(FullAdder_1115_io_b),
    .io_ci(FullAdder_1115_io_ci),
    .io_s(FullAdder_1115_io_s),
    .io_co(FullAdder_1115_io_co)
  );
  FullAdder FullAdder_1116 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1116_io_a),
    .io_b(FullAdder_1116_io_b),
    .io_ci(FullAdder_1116_io_ci),
    .io_s(FullAdder_1116_io_s),
    .io_co(FullAdder_1116_io_co)
  );
  FullAdder FullAdder_1117 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1117_io_a),
    .io_b(FullAdder_1117_io_b),
    .io_ci(FullAdder_1117_io_ci),
    .io_s(FullAdder_1117_io_s),
    .io_co(FullAdder_1117_io_co)
  );
  FullAdder FullAdder_1118 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1118_io_a),
    .io_b(FullAdder_1118_io_b),
    .io_ci(FullAdder_1118_io_ci),
    .io_s(FullAdder_1118_io_s),
    .io_co(FullAdder_1118_io_co)
  );
  FullAdder FullAdder_1119 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1119_io_a),
    .io_b(FullAdder_1119_io_b),
    .io_ci(FullAdder_1119_io_ci),
    .io_s(FullAdder_1119_io_s),
    .io_co(FullAdder_1119_io_co)
  );
  FullAdder FullAdder_1120 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1120_io_a),
    .io_b(FullAdder_1120_io_b),
    .io_ci(FullAdder_1120_io_ci),
    .io_s(FullAdder_1120_io_s),
    .io_co(FullAdder_1120_io_co)
  );
  FullAdder FullAdder_1121 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1121_io_a),
    .io_b(FullAdder_1121_io_b),
    .io_ci(FullAdder_1121_io_ci),
    .io_s(FullAdder_1121_io_s),
    .io_co(FullAdder_1121_io_co)
  );
  FullAdder FullAdder_1122 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1122_io_a),
    .io_b(FullAdder_1122_io_b),
    .io_ci(FullAdder_1122_io_ci),
    .io_s(FullAdder_1122_io_s),
    .io_co(FullAdder_1122_io_co)
  );
  FullAdder FullAdder_1123 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1123_io_a),
    .io_b(FullAdder_1123_io_b),
    .io_ci(FullAdder_1123_io_ci),
    .io_s(FullAdder_1123_io_s),
    .io_co(FullAdder_1123_io_co)
  );
  FullAdder FullAdder_1124 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1124_io_a),
    .io_b(FullAdder_1124_io_b),
    .io_ci(FullAdder_1124_io_ci),
    .io_s(FullAdder_1124_io_s),
    .io_co(FullAdder_1124_io_co)
  );
  FullAdder FullAdder_1125 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1125_io_a),
    .io_b(FullAdder_1125_io_b),
    .io_ci(FullAdder_1125_io_ci),
    .io_s(FullAdder_1125_io_s),
    .io_co(FullAdder_1125_io_co)
  );
  FullAdder FullAdder_1126 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1126_io_a),
    .io_b(FullAdder_1126_io_b),
    .io_ci(FullAdder_1126_io_ci),
    .io_s(FullAdder_1126_io_s),
    .io_co(FullAdder_1126_io_co)
  );
  FullAdder FullAdder_1127 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1127_io_a),
    .io_b(FullAdder_1127_io_b),
    .io_ci(FullAdder_1127_io_ci),
    .io_s(FullAdder_1127_io_s),
    .io_co(FullAdder_1127_io_co)
  );
  FullAdder FullAdder_1128 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1128_io_a),
    .io_b(FullAdder_1128_io_b),
    .io_ci(FullAdder_1128_io_ci),
    .io_s(FullAdder_1128_io_s),
    .io_co(FullAdder_1128_io_co)
  );
  FullAdder FullAdder_1129 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1129_io_a),
    .io_b(FullAdder_1129_io_b),
    .io_ci(FullAdder_1129_io_ci),
    .io_s(FullAdder_1129_io_s),
    .io_co(FullAdder_1129_io_co)
  );
  FullAdder FullAdder_1130 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1130_io_a),
    .io_b(FullAdder_1130_io_b),
    .io_ci(FullAdder_1130_io_ci),
    .io_s(FullAdder_1130_io_s),
    .io_co(FullAdder_1130_io_co)
  );
  FullAdder FullAdder_1131 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1131_io_a),
    .io_b(FullAdder_1131_io_b),
    .io_ci(FullAdder_1131_io_ci),
    .io_s(FullAdder_1131_io_s),
    .io_co(FullAdder_1131_io_co)
  );
  FullAdder FullAdder_1132 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1132_io_a),
    .io_b(FullAdder_1132_io_b),
    .io_ci(FullAdder_1132_io_ci),
    .io_s(FullAdder_1132_io_s),
    .io_co(FullAdder_1132_io_co)
  );
  FullAdder FullAdder_1133 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1133_io_a),
    .io_b(FullAdder_1133_io_b),
    .io_ci(FullAdder_1133_io_ci),
    .io_s(FullAdder_1133_io_s),
    .io_co(FullAdder_1133_io_co)
  );
  FullAdder FullAdder_1134 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1134_io_a),
    .io_b(FullAdder_1134_io_b),
    .io_ci(FullAdder_1134_io_ci),
    .io_s(FullAdder_1134_io_s),
    .io_co(FullAdder_1134_io_co)
  );
  FullAdder FullAdder_1135 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1135_io_a),
    .io_b(FullAdder_1135_io_b),
    .io_ci(FullAdder_1135_io_ci),
    .io_s(FullAdder_1135_io_s),
    .io_co(FullAdder_1135_io_co)
  );
  HalfAdder HalfAdder_23 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_23_io_a),
    .io_b(HalfAdder_23_io_b),
    .io_s(HalfAdder_23_io_s),
    .io_co(HalfAdder_23_io_co)
  );
  FullAdder FullAdder_1136 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1136_io_a),
    .io_b(FullAdder_1136_io_b),
    .io_ci(FullAdder_1136_io_ci),
    .io_s(FullAdder_1136_io_s),
    .io_co(FullAdder_1136_io_co)
  );
  FullAdder FullAdder_1137 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1137_io_a),
    .io_b(FullAdder_1137_io_b),
    .io_ci(FullAdder_1137_io_ci),
    .io_s(FullAdder_1137_io_s),
    .io_co(FullAdder_1137_io_co)
  );
  FullAdder FullAdder_1138 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1138_io_a),
    .io_b(FullAdder_1138_io_b),
    .io_ci(FullAdder_1138_io_ci),
    .io_s(FullAdder_1138_io_s),
    .io_co(FullAdder_1138_io_co)
  );
  FullAdder FullAdder_1139 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1139_io_a),
    .io_b(FullAdder_1139_io_b),
    .io_ci(FullAdder_1139_io_ci),
    .io_s(FullAdder_1139_io_s),
    .io_co(FullAdder_1139_io_co)
  );
  FullAdder FullAdder_1140 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1140_io_a),
    .io_b(FullAdder_1140_io_b),
    .io_ci(FullAdder_1140_io_ci),
    .io_s(FullAdder_1140_io_s),
    .io_co(FullAdder_1140_io_co)
  );
  FullAdder FullAdder_1141 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1141_io_a),
    .io_b(FullAdder_1141_io_b),
    .io_ci(FullAdder_1141_io_ci),
    .io_s(FullAdder_1141_io_s),
    .io_co(FullAdder_1141_io_co)
  );
  FullAdder FullAdder_1142 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1142_io_a),
    .io_b(FullAdder_1142_io_b),
    .io_ci(FullAdder_1142_io_ci),
    .io_s(FullAdder_1142_io_s),
    .io_co(FullAdder_1142_io_co)
  );
  FullAdder FullAdder_1143 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1143_io_a),
    .io_b(FullAdder_1143_io_b),
    .io_ci(FullAdder_1143_io_ci),
    .io_s(FullAdder_1143_io_s),
    .io_co(FullAdder_1143_io_co)
  );
  FullAdder FullAdder_1144 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1144_io_a),
    .io_b(FullAdder_1144_io_b),
    .io_ci(FullAdder_1144_io_ci),
    .io_s(FullAdder_1144_io_s),
    .io_co(FullAdder_1144_io_co)
  );
  FullAdder FullAdder_1145 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1145_io_a),
    .io_b(FullAdder_1145_io_b),
    .io_ci(FullAdder_1145_io_ci),
    .io_s(FullAdder_1145_io_s),
    .io_co(FullAdder_1145_io_co)
  );
  FullAdder FullAdder_1146 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1146_io_a),
    .io_b(FullAdder_1146_io_b),
    .io_ci(FullAdder_1146_io_ci),
    .io_s(FullAdder_1146_io_s),
    .io_co(FullAdder_1146_io_co)
  );
  FullAdder FullAdder_1147 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1147_io_a),
    .io_b(FullAdder_1147_io_b),
    .io_ci(FullAdder_1147_io_ci),
    .io_s(FullAdder_1147_io_s),
    .io_co(FullAdder_1147_io_co)
  );
  FullAdder FullAdder_1148 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1148_io_a),
    .io_b(FullAdder_1148_io_b),
    .io_ci(FullAdder_1148_io_ci),
    .io_s(FullAdder_1148_io_s),
    .io_co(FullAdder_1148_io_co)
  );
  FullAdder FullAdder_1149 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1149_io_a),
    .io_b(FullAdder_1149_io_b),
    .io_ci(FullAdder_1149_io_ci),
    .io_s(FullAdder_1149_io_s),
    .io_co(FullAdder_1149_io_co)
  );
  FullAdder FullAdder_1150 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1150_io_a),
    .io_b(FullAdder_1150_io_b),
    .io_ci(FullAdder_1150_io_ci),
    .io_s(FullAdder_1150_io_s),
    .io_co(FullAdder_1150_io_co)
  );
  FullAdder FullAdder_1151 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1151_io_a),
    .io_b(FullAdder_1151_io_b),
    .io_ci(FullAdder_1151_io_ci),
    .io_s(FullAdder_1151_io_s),
    .io_co(FullAdder_1151_io_co)
  );
  FullAdder FullAdder_1152 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1152_io_a),
    .io_b(FullAdder_1152_io_b),
    .io_ci(FullAdder_1152_io_ci),
    .io_s(FullAdder_1152_io_s),
    .io_co(FullAdder_1152_io_co)
  );
  FullAdder FullAdder_1153 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1153_io_a),
    .io_b(FullAdder_1153_io_b),
    .io_ci(FullAdder_1153_io_ci),
    .io_s(FullAdder_1153_io_s),
    .io_co(FullAdder_1153_io_co)
  );
  FullAdder FullAdder_1154 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1154_io_a),
    .io_b(FullAdder_1154_io_b),
    .io_ci(FullAdder_1154_io_ci),
    .io_s(FullAdder_1154_io_s),
    .io_co(FullAdder_1154_io_co)
  );
  FullAdder FullAdder_1155 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1155_io_a),
    .io_b(FullAdder_1155_io_b),
    .io_ci(FullAdder_1155_io_ci),
    .io_s(FullAdder_1155_io_s),
    .io_co(FullAdder_1155_io_co)
  );
  FullAdder FullAdder_1156 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1156_io_a),
    .io_b(FullAdder_1156_io_b),
    .io_ci(FullAdder_1156_io_ci),
    .io_s(FullAdder_1156_io_s),
    .io_co(FullAdder_1156_io_co)
  );
  FullAdder FullAdder_1157 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1157_io_a),
    .io_b(FullAdder_1157_io_b),
    .io_ci(FullAdder_1157_io_ci),
    .io_s(FullAdder_1157_io_s),
    .io_co(FullAdder_1157_io_co)
  );
  FullAdder FullAdder_1158 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1158_io_a),
    .io_b(FullAdder_1158_io_b),
    .io_ci(FullAdder_1158_io_ci),
    .io_s(FullAdder_1158_io_s),
    .io_co(FullAdder_1158_io_co)
  );
  FullAdder FullAdder_1159 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1159_io_a),
    .io_b(FullAdder_1159_io_b),
    .io_ci(FullAdder_1159_io_ci),
    .io_s(FullAdder_1159_io_s),
    .io_co(FullAdder_1159_io_co)
  );
  FullAdder FullAdder_1160 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1160_io_a),
    .io_b(FullAdder_1160_io_b),
    .io_ci(FullAdder_1160_io_ci),
    .io_s(FullAdder_1160_io_s),
    .io_co(FullAdder_1160_io_co)
  );
  FullAdder FullAdder_1161 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1161_io_a),
    .io_b(FullAdder_1161_io_b),
    .io_ci(FullAdder_1161_io_ci),
    .io_s(FullAdder_1161_io_s),
    .io_co(FullAdder_1161_io_co)
  );
  FullAdder FullAdder_1162 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1162_io_a),
    .io_b(FullAdder_1162_io_b),
    .io_ci(FullAdder_1162_io_ci),
    .io_s(FullAdder_1162_io_s),
    .io_co(FullAdder_1162_io_co)
  );
  FullAdder FullAdder_1163 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1163_io_a),
    .io_b(FullAdder_1163_io_b),
    .io_ci(FullAdder_1163_io_ci),
    .io_s(FullAdder_1163_io_s),
    .io_co(FullAdder_1163_io_co)
  );
  FullAdder FullAdder_1164 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1164_io_a),
    .io_b(FullAdder_1164_io_b),
    .io_ci(FullAdder_1164_io_ci),
    .io_s(FullAdder_1164_io_s),
    .io_co(FullAdder_1164_io_co)
  );
  FullAdder FullAdder_1165 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1165_io_a),
    .io_b(FullAdder_1165_io_b),
    .io_ci(FullAdder_1165_io_ci),
    .io_s(FullAdder_1165_io_s),
    .io_co(FullAdder_1165_io_co)
  );
  FullAdder FullAdder_1166 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1166_io_a),
    .io_b(FullAdder_1166_io_b),
    .io_ci(FullAdder_1166_io_ci),
    .io_s(FullAdder_1166_io_s),
    .io_co(FullAdder_1166_io_co)
  );
  FullAdder FullAdder_1167 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1167_io_a),
    .io_b(FullAdder_1167_io_b),
    .io_ci(FullAdder_1167_io_ci),
    .io_s(FullAdder_1167_io_s),
    .io_co(FullAdder_1167_io_co)
  );
  HalfAdder HalfAdder_24 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_24_io_a),
    .io_b(HalfAdder_24_io_b),
    .io_s(HalfAdder_24_io_s),
    .io_co(HalfAdder_24_io_co)
  );
  FullAdder FullAdder_1168 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1168_io_a),
    .io_b(FullAdder_1168_io_b),
    .io_ci(FullAdder_1168_io_ci),
    .io_s(FullAdder_1168_io_s),
    .io_co(FullAdder_1168_io_co)
  );
  FullAdder FullAdder_1169 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1169_io_a),
    .io_b(FullAdder_1169_io_b),
    .io_ci(FullAdder_1169_io_ci),
    .io_s(FullAdder_1169_io_s),
    .io_co(FullAdder_1169_io_co)
  );
  FullAdder FullAdder_1170 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1170_io_a),
    .io_b(FullAdder_1170_io_b),
    .io_ci(FullAdder_1170_io_ci),
    .io_s(FullAdder_1170_io_s),
    .io_co(FullAdder_1170_io_co)
  );
  FullAdder FullAdder_1171 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1171_io_a),
    .io_b(FullAdder_1171_io_b),
    .io_ci(FullAdder_1171_io_ci),
    .io_s(FullAdder_1171_io_s),
    .io_co(FullAdder_1171_io_co)
  );
  FullAdder FullAdder_1172 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1172_io_a),
    .io_b(FullAdder_1172_io_b),
    .io_ci(FullAdder_1172_io_ci),
    .io_s(FullAdder_1172_io_s),
    .io_co(FullAdder_1172_io_co)
  );
  FullAdder FullAdder_1173 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1173_io_a),
    .io_b(FullAdder_1173_io_b),
    .io_ci(FullAdder_1173_io_ci),
    .io_s(FullAdder_1173_io_s),
    .io_co(FullAdder_1173_io_co)
  );
  FullAdder FullAdder_1174 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1174_io_a),
    .io_b(FullAdder_1174_io_b),
    .io_ci(FullAdder_1174_io_ci),
    .io_s(FullAdder_1174_io_s),
    .io_co(FullAdder_1174_io_co)
  );
  FullAdder FullAdder_1175 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1175_io_a),
    .io_b(FullAdder_1175_io_b),
    .io_ci(FullAdder_1175_io_ci),
    .io_s(FullAdder_1175_io_s),
    .io_co(FullAdder_1175_io_co)
  );
  FullAdder FullAdder_1176 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1176_io_a),
    .io_b(FullAdder_1176_io_b),
    .io_ci(FullAdder_1176_io_ci),
    .io_s(FullAdder_1176_io_s),
    .io_co(FullAdder_1176_io_co)
  );
  FullAdder FullAdder_1177 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1177_io_a),
    .io_b(FullAdder_1177_io_b),
    .io_ci(FullAdder_1177_io_ci),
    .io_s(FullAdder_1177_io_s),
    .io_co(FullAdder_1177_io_co)
  );
  FullAdder FullAdder_1178 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1178_io_a),
    .io_b(FullAdder_1178_io_b),
    .io_ci(FullAdder_1178_io_ci),
    .io_s(FullAdder_1178_io_s),
    .io_co(FullAdder_1178_io_co)
  );
  FullAdder FullAdder_1179 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1179_io_a),
    .io_b(FullAdder_1179_io_b),
    .io_ci(FullAdder_1179_io_ci),
    .io_s(FullAdder_1179_io_s),
    .io_co(FullAdder_1179_io_co)
  );
  FullAdder FullAdder_1180 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1180_io_a),
    .io_b(FullAdder_1180_io_b),
    .io_ci(FullAdder_1180_io_ci),
    .io_s(FullAdder_1180_io_s),
    .io_co(FullAdder_1180_io_co)
  );
  FullAdder FullAdder_1181 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1181_io_a),
    .io_b(FullAdder_1181_io_b),
    .io_ci(FullAdder_1181_io_ci),
    .io_s(FullAdder_1181_io_s),
    .io_co(FullAdder_1181_io_co)
  );
  FullAdder FullAdder_1182 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1182_io_a),
    .io_b(FullAdder_1182_io_b),
    .io_ci(FullAdder_1182_io_ci),
    .io_s(FullAdder_1182_io_s),
    .io_co(FullAdder_1182_io_co)
  );
  FullAdder FullAdder_1183 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1183_io_a),
    .io_b(FullAdder_1183_io_b),
    .io_ci(FullAdder_1183_io_ci),
    .io_s(FullAdder_1183_io_s),
    .io_co(FullAdder_1183_io_co)
  );
  FullAdder FullAdder_1184 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1184_io_a),
    .io_b(FullAdder_1184_io_b),
    .io_ci(FullAdder_1184_io_ci),
    .io_s(FullAdder_1184_io_s),
    .io_co(FullAdder_1184_io_co)
  );
  FullAdder FullAdder_1185 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1185_io_a),
    .io_b(FullAdder_1185_io_b),
    .io_ci(FullAdder_1185_io_ci),
    .io_s(FullAdder_1185_io_s),
    .io_co(FullAdder_1185_io_co)
  );
  FullAdder FullAdder_1186 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1186_io_a),
    .io_b(FullAdder_1186_io_b),
    .io_ci(FullAdder_1186_io_ci),
    .io_s(FullAdder_1186_io_s),
    .io_co(FullAdder_1186_io_co)
  );
  FullAdder FullAdder_1187 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1187_io_a),
    .io_b(FullAdder_1187_io_b),
    .io_ci(FullAdder_1187_io_ci),
    .io_s(FullAdder_1187_io_s),
    .io_co(FullAdder_1187_io_co)
  );
  FullAdder FullAdder_1188 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1188_io_a),
    .io_b(FullAdder_1188_io_b),
    .io_ci(FullAdder_1188_io_ci),
    .io_s(FullAdder_1188_io_s),
    .io_co(FullAdder_1188_io_co)
  );
  FullAdder FullAdder_1189 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1189_io_a),
    .io_b(FullAdder_1189_io_b),
    .io_ci(FullAdder_1189_io_ci),
    .io_s(FullAdder_1189_io_s),
    .io_co(FullAdder_1189_io_co)
  );
  FullAdder FullAdder_1190 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1190_io_a),
    .io_b(FullAdder_1190_io_b),
    .io_ci(FullAdder_1190_io_ci),
    .io_s(FullAdder_1190_io_s),
    .io_co(FullAdder_1190_io_co)
  );
  FullAdder FullAdder_1191 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1191_io_a),
    .io_b(FullAdder_1191_io_b),
    .io_ci(FullAdder_1191_io_ci),
    .io_s(FullAdder_1191_io_s),
    .io_co(FullAdder_1191_io_co)
  );
  FullAdder FullAdder_1192 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1192_io_a),
    .io_b(FullAdder_1192_io_b),
    .io_ci(FullAdder_1192_io_ci),
    .io_s(FullAdder_1192_io_s),
    .io_co(FullAdder_1192_io_co)
  );
  FullAdder FullAdder_1193 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1193_io_a),
    .io_b(FullAdder_1193_io_b),
    .io_ci(FullAdder_1193_io_ci),
    .io_s(FullAdder_1193_io_s),
    .io_co(FullAdder_1193_io_co)
  );
  FullAdder FullAdder_1194 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1194_io_a),
    .io_b(FullAdder_1194_io_b),
    .io_ci(FullAdder_1194_io_ci),
    .io_s(FullAdder_1194_io_s),
    .io_co(FullAdder_1194_io_co)
  );
  FullAdder FullAdder_1195 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1195_io_a),
    .io_b(FullAdder_1195_io_b),
    .io_ci(FullAdder_1195_io_ci),
    .io_s(FullAdder_1195_io_s),
    .io_co(FullAdder_1195_io_co)
  );
  FullAdder FullAdder_1196 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1196_io_a),
    .io_b(FullAdder_1196_io_b),
    .io_ci(FullAdder_1196_io_ci),
    .io_s(FullAdder_1196_io_s),
    .io_co(FullAdder_1196_io_co)
  );
  HalfAdder HalfAdder_25 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_25_io_a),
    .io_b(HalfAdder_25_io_b),
    .io_s(HalfAdder_25_io_s),
    .io_co(HalfAdder_25_io_co)
  );
  FullAdder FullAdder_1197 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1197_io_a),
    .io_b(FullAdder_1197_io_b),
    .io_ci(FullAdder_1197_io_ci),
    .io_s(FullAdder_1197_io_s),
    .io_co(FullAdder_1197_io_co)
  );
  FullAdder FullAdder_1198 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1198_io_a),
    .io_b(FullAdder_1198_io_b),
    .io_ci(FullAdder_1198_io_ci),
    .io_s(FullAdder_1198_io_s),
    .io_co(FullAdder_1198_io_co)
  );
  FullAdder FullAdder_1199 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1199_io_a),
    .io_b(FullAdder_1199_io_b),
    .io_ci(FullAdder_1199_io_ci),
    .io_s(FullAdder_1199_io_s),
    .io_co(FullAdder_1199_io_co)
  );
  FullAdder FullAdder_1200 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1200_io_a),
    .io_b(FullAdder_1200_io_b),
    .io_ci(FullAdder_1200_io_ci),
    .io_s(FullAdder_1200_io_s),
    .io_co(FullAdder_1200_io_co)
  );
  FullAdder FullAdder_1201 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1201_io_a),
    .io_b(FullAdder_1201_io_b),
    .io_ci(FullAdder_1201_io_ci),
    .io_s(FullAdder_1201_io_s),
    .io_co(FullAdder_1201_io_co)
  );
  FullAdder FullAdder_1202 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1202_io_a),
    .io_b(FullAdder_1202_io_b),
    .io_ci(FullAdder_1202_io_ci),
    .io_s(FullAdder_1202_io_s),
    .io_co(FullAdder_1202_io_co)
  );
  FullAdder FullAdder_1203 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1203_io_a),
    .io_b(FullAdder_1203_io_b),
    .io_ci(FullAdder_1203_io_ci),
    .io_s(FullAdder_1203_io_s),
    .io_co(FullAdder_1203_io_co)
  );
  FullAdder FullAdder_1204 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1204_io_a),
    .io_b(FullAdder_1204_io_b),
    .io_ci(FullAdder_1204_io_ci),
    .io_s(FullAdder_1204_io_s),
    .io_co(FullAdder_1204_io_co)
  );
  FullAdder FullAdder_1205 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1205_io_a),
    .io_b(FullAdder_1205_io_b),
    .io_ci(FullAdder_1205_io_ci),
    .io_s(FullAdder_1205_io_s),
    .io_co(FullAdder_1205_io_co)
  );
  FullAdder FullAdder_1206 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1206_io_a),
    .io_b(FullAdder_1206_io_b),
    .io_ci(FullAdder_1206_io_ci),
    .io_s(FullAdder_1206_io_s),
    .io_co(FullAdder_1206_io_co)
  );
  FullAdder FullAdder_1207 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1207_io_a),
    .io_b(FullAdder_1207_io_b),
    .io_ci(FullAdder_1207_io_ci),
    .io_s(FullAdder_1207_io_s),
    .io_co(FullAdder_1207_io_co)
  );
  FullAdder FullAdder_1208 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1208_io_a),
    .io_b(FullAdder_1208_io_b),
    .io_ci(FullAdder_1208_io_ci),
    .io_s(FullAdder_1208_io_s),
    .io_co(FullAdder_1208_io_co)
  );
  FullAdder FullAdder_1209 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1209_io_a),
    .io_b(FullAdder_1209_io_b),
    .io_ci(FullAdder_1209_io_ci),
    .io_s(FullAdder_1209_io_s),
    .io_co(FullAdder_1209_io_co)
  );
  FullAdder FullAdder_1210 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1210_io_a),
    .io_b(FullAdder_1210_io_b),
    .io_ci(FullAdder_1210_io_ci),
    .io_s(FullAdder_1210_io_s),
    .io_co(FullAdder_1210_io_co)
  );
  FullAdder FullAdder_1211 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1211_io_a),
    .io_b(FullAdder_1211_io_b),
    .io_ci(FullAdder_1211_io_ci),
    .io_s(FullAdder_1211_io_s),
    .io_co(FullAdder_1211_io_co)
  );
  FullAdder FullAdder_1212 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1212_io_a),
    .io_b(FullAdder_1212_io_b),
    .io_ci(FullAdder_1212_io_ci),
    .io_s(FullAdder_1212_io_s),
    .io_co(FullAdder_1212_io_co)
  );
  FullAdder FullAdder_1213 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1213_io_a),
    .io_b(FullAdder_1213_io_b),
    .io_ci(FullAdder_1213_io_ci),
    .io_s(FullAdder_1213_io_s),
    .io_co(FullAdder_1213_io_co)
  );
  FullAdder FullAdder_1214 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1214_io_a),
    .io_b(FullAdder_1214_io_b),
    .io_ci(FullAdder_1214_io_ci),
    .io_s(FullAdder_1214_io_s),
    .io_co(FullAdder_1214_io_co)
  );
  FullAdder FullAdder_1215 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1215_io_a),
    .io_b(FullAdder_1215_io_b),
    .io_ci(FullAdder_1215_io_ci),
    .io_s(FullAdder_1215_io_s),
    .io_co(FullAdder_1215_io_co)
  );
  FullAdder FullAdder_1216 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1216_io_a),
    .io_b(FullAdder_1216_io_b),
    .io_ci(FullAdder_1216_io_ci),
    .io_s(FullAdder_1216_io_s),
    .io_co(FullAdder_1216_io_co)
  );
  FullAdder FullAdder_1217 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1217_io_a),
    .io_b(FullAdder_1217_io_b),
    .io_ci(FullAdder_1217_io_ci),
    .io_s(FullAdder_1217_io_s),
    .io_co(FullAdder_1217_io_co)
  );
  FullAdder FullAdder_1218 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1218_io_a),
    .io_b(FullAdder_1218_io_b),
    .io_ci(FullAdder_1218_io_ci),
    .io_s(FullAdder_1218_io_s),
    .io_co(FullAdder_1218_io_co)
  );
  FullAdder FullAdder_1219 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1219_io_a),
    .io_b(FullAdder_1219_io_b),
    .io_ci(FullAdder_1219_io_ci),
    .io_s(FullAdder_1219_io_s),
    .io_co(FullAdder_1219_io_co)
  );
  FullAdder FullAdder_1220 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1220_io_a),
    .io_b(FullAdder_1220_io_b),
    .io_ci(FullAdder_1220_io_ci),
    .io_s(FullAdder_1220_io_s),
    .io_co(FullAdder_1220_io_co)
  );
  FullAdder FullAdder_1221 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1221_io_a),
    .io_b(FullAdder_1221_io_b),
    .io_ci(FullAdder_1221_io_ci),
    .io_s(FullAdder_1221_io_s),
    .io_co(FullAdder_1221_io_co)
  );
  FullAdder FullAdder_1222 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1222_io_a),
    .io_b(FullAdder_1222_io_b),
    .io_ci(FullAdder_1222_io_ci),
    .io_s(FullAdder_1222_io_s),
    .io_co(FullAdder_1222_io_co)
  );
  FullAdder FullAdder_1223 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1223_io_a),
    .io_b(FullAdder_1223_io_b),
    .io_ci(FullAdder_1223_io_ci),
    .io_s(FullAdder_1223_io_s),
    .io_co(FullAdder_1223_io_co)
  );
  FullAdder FullAdder_1224 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1224_io_a),
    .io_b(FullAdder_1224_io_b),
    .io_ci(FullAdder_1224_io_ci),
    .io_s(FullAdder_1224_io_s),
    .io_co(FullAdder_1224_io_co)
  );
  FullAdder FullAdder_1225 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1225_io_a),
    .io_b(FullAdder_1225_io_b),
    .io_ci(FullAdder_1225_io_ci),
    .io_s(FullAdder_1225_io_s),
    .io_co(FullAdder_1225_io_co)
  );
  FullAdder FullAdder_1226 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1226_io_a),
    .io_b(FullAdder_1226_io_b),
    .io_ci(FullAdder_1226_io_ci),
    .io_s(FullAdder_1226_io_s),
    .io_co(FullAdder_1226_io_co)
  );
  FullAdder FullAdder_1227 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1227_io_a),
    .io_b(FullAdder_1227_io_b),
    .io_ci(FullAdder_1227_io_ci),
    .io_s(FullAdder_1227_io_s),
    .io_co(FullAdder_1227_io_co)
  );
  FullAdder FullAdder_1228 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1228_io_a),
    .io_b(FullAdder_1228_io_b),
    .io_ci(FullAdder_1228_io_ci),
    .io_s(FullAdder_1228_io_s),
    .io_co(FullAdder_1228_io_co)
  );
  FullAdder FullAdder_1229 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1229_io_a),
    .io_b(FullAdder_1229_io_b),
    .io_ci(FullAdder_1229_io_ci),
    .io_s(FullAdder_1229_io_s),
    .io_co(FullAdder_1229_io_co)
  );
  FullAdder FullAdder_1230 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1230_io_a),
    .io_b(FullAdder_1230_io_b),
    .io_ci(FullAdder_1230_io_ci),
    .io_s(FullAdder_1230_io_s),
    .io_co(FullAdder_1230_io_co)
  );
  FullAdder FullAdder_1231 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1231_io_a),
    .io_b(FullAdder_1231_io_b),
    .io_ci(FullAdder_1231_io_ci),
    .io_s(FullAdder_1231_io_s),
    .io_co(FullAdder_1231_io_co)
  );
  FullAdder FullAdder_1232 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1232_io_a),
    .io_b(FullAdder_1232_io_b),
    .io_ci(FullAdder_1232_io_ci),
    .io_s(FullAdder_1232_io_s),
    .io_co(FullAdder_1232_io_co)
  );
  FullAdder FullAdder_1233 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1233_io_a),
    .io_b(FullAdder_1233_io_b),
    .io_ci(FullAdder_1233_io_ci),
    .io_s(FullAdder_1233_io_s),
    .io_co(FullAdder_1233_io_co)
  );
  FullAdder FullAdder_1234 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1234_io_a),
    .io_b(FullAdder_1234_io_b),
    .io_ci(FullAdder_1234_io_ci),
    .io_s(FullAdder_1234_io_s),
    .io_co(FullAdder_1234_io_co)
  );
  FullAdder FullAdder_1235 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1235_io_a),
    .io_b(FullAdder_1235_io_b),
    .io_ci(FullAdder_1235_io_ci),
    .io_s(FullAdder_1235_io_s),
    .io_co(FullAdder_1235_io_co)
  );
  FullAdder FullAdder_1236 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1236_io_a),
    .io_b(FullAdder_1236_io_b),
    .io_ci(FullAdder_1236_io_ci),
    .io_s(FullAdder_1236_io_s),
    .io_co(FullAdder_1236_io_co)
  );
  FullAdder FullAdder_1237 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1237_io_a),
    .io_b(FullAdder_1237_io_b),
    .io_ci(FullAdder_1237_io_ci),
    .io_s(FullAdder_1237_io_s),
    .io_co(FullAdder_1237_io_co)
  );
  FullAdder FullAdder_1238 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1238_io_a),
    .io_b(FullAdder_1238_io_b),
    .io_ci(FullAdder_1238_io_ci),
    .io_s(FullAdder_1238_io_s),
    .io_co(FullAdder_1238_io_co)
  );
  FullAdder FullAdder_1239 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1239_io_a),
    .io_b(FullAdder_1239_io_b),
    .io_ci(FullAdder_1239_io_ci),
    .io_s(FullAdder_1239_io_s),
    .io_co(FullAdder_1239_io_co)
  );
  FullAdder FullAdder_1240 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1240_io_a),
    .io_b(FullAdder_1240_io_b),
    .io_ci(FullAdder_1240_io_ci),
    .io_s(FullAdder_1240_io_s),
    .io_co(FullAdder_1240_io_co)
  );
  FullAdder FullAdder_1241 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1241_io_a),
    .io_b(FullAdder_1241_io_b),
    .io_ci(FullAdder_1241_io_ci),
    .io_s(FullAdder_1241_io_s),
    .io_co(FullAdder_1241_io_co)
  );
  FullAdder FullAdder_1242 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1242_io_a),
    .io_b(FullAdder_1242_io_b),
    .io_ci(FullAdder_1242_io_ci),
    .io_s(FullAdder_1242_io_s),
    .io_co(FullAdder_1242_io_co)
  );
  FullAdder FullAdder_1243 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1243_io_a),
    .io_b(FullAdder_1243_io_b),
    .io_ci(FullAdder_1243_io_ci),
    .io_s(FullAdder_1243_io_s),
    .io_co(FullAdder_1243_io_co)
  );
  FullAdder FullAdder_1244 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1244_io_a),
    .io_b(FullAdder_1244_io_b),
    .io_ci(FullAdder_1244_io_ci),
    .io_s(FullAdder_1244_io_s),
    .io_co(FullAdder_1244_io_co)
  );
  FullAdder FullAdder_1245 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1245_io_a),
    .io_b(FullAdder_1245_io_b),
    .io_ci(FullAdder_1245_io_ci),
    .io_s(FullAdder_1245_io_s),
    .io_co(FullAdder_1245_io_co)
  );
  HalfAdder HalfAdder_26 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_26_io_a),
    .io_b(HalfAdder_26_io_b),
    .io_s(HalfAdder_26_io_s),
    .io_co(HalfAdder_26_io_co)
  );
  FullAdder FullAdder_1246 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1246_io_a),
    .io_b(FullAdder_1246_io_b),
    .io_ci(FullAdder_1246_io_ci),
    .io_s(FullAdder_1246_io_s),
    .io_co(FullAdder_1246_io_co)
  );
  FullAdder FullAdder_1247 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1247_io_a),
    .io_b(FullAdder_1247_io_b),
    .io_ci(FullAdder_1247_io_ci),
    .io_s(FullAdder_1247_io_s),
    .io_co(FullAdder_1247_io_co)
  );
  FullAdder FullAdder_1248 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1248_io_a),
    .io_b(FullAdder_1248_io_b),
    .io_ci(FullAdder_1248_io_ci),
    .io_s(FullAdder_1248_io_s),
    .io_co(FullAdder_1248_io_co)
  );
  FullAdder FullAdder_1249 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1249_io_a),
    .io_b(FullAdder_1249_io_b),
    .io_ci(FullAdder_1249_io_ci),
    .io_s(FullAdder_1249_io_s),
    .io_co(FullAdder_1249_io_co)
  );
  FullAdder FullAdder_1250 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1250_io_a),
    .io_b(FullAdder_1250_io_b),
    .io_ci(FullAdder_1250_io_ci),
    .io_s(FullAdder_1250_io_s),
    .io_co(FullAdder_1250_io_co)
  );
  FullAdder FullAdder_1251 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1251_io_a),
    .io_b(FullAdder_1251_io_b),
    .io_ci(FullAdder_1251_io_ci),
    .io_s(FullAdder_1251_io_s),
    .io_co(FullAdder_1251_io_co)
  );
  FullAdder FullAdder_1252 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1252_io_a),
    .io_b(FullAdder_1252_io_b),
    .io_ci(FullAdder_1252_io_ci),
    .io_s(FullAdder_1252_io_s),
    .io_co(FullAdder_1252_io_co)
  );
  FullAdder FullAdder_1253 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1253_io_a),
    .io_b(FullAdder_1253_io_b),
    .io_ci(FullAdder_1253_io_ci),
    .io_s(FullAdder_1253_io_s),
    .io_co(FullAdder_1253_io_co)
  );
  FullAdder FullAdder_1254 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1254_io_a),
    .io_b(FullAdder_1254_io_b),
    .io_ci(FullAdder_1254_io_ci),
    .io_s(FullAdder_1254_io_s),
    .io_co(FullAdder_1254_io_co)
  );
  FullAdder FullAdder_1255 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1255_io_a),
    .io_b(FullAdder_1255_io_b),
    .io_ci(FullAdder_1255_io_ci),
    .io_s(FullAdder_1255_io_s),
    .io_co(FullAdder_1255_io_co)
  );
  FullAdder FullAdder_1256 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1256_io_a),
    .io_b(FullAdder_1256_io_b),
    .io_ci(FullAdder_1256_io_ci),
    .io_s(FullAdder_1256_io_s),
    .io_co(FullAdder_1256_io_co)
  );
  FullAdder FullAdder_1257 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1257_io_a),
    .io_b(FullAdder_1257_io_b),
    .io_ci(FullAdder_1257_io_ci),
    .io_s(FullAdder_1257_io_s),
    .io_co(FullAdder_1257_io_co)
  );
  FullAdder FullAdder_1258 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1258_io_a),
    .io_b(FullAdder_1258_io_b),
    .io_ci(FullAdder_1258_io_ci),
    .io_s(FullAdder_1258_io_s),
    .io_co(FullAdder_1258_io_co)
  );
  FullAdder FullAdder_1259 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1259_io_a),
    .io_b(FullAdder_1259_io_b),
    .io_ci(FullAdder_1259_io_ci),
    .io_s(FullAdder_1259_io_s),
    .io_co(FullAdder_1259_io_co)
  );
  FullAdder FullAdder_1260 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1260_io_a),
    .io_b(FullAdder_1260_io_b),
    .io_ci(FullAdder_1260_io_ci),
    .io_s(FullAdder_1260_io_s),
    .io_co(FullAdder_1260_io_co)
  );
  FullAdder FullAdder_1261 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1261_io_a),
    .io_b(FullAdder_1261_io_b),
    .io_ci(FullAdder_1261_io_ci),
    .io_s(FullAdder_1261_io_s),
    .io_co(FullAdder_1261_io_co)
  );
  FullAdder FullAdder_1262 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1262_io_a),
    .io_b(FullAdder_1262_io_b),
    .io_ci(FullAdder_1262_io_ci),
    .io_s(FullAdder_1262_io_s),
    .io_co(FullAdder_1262_io_co)
  );
  FullAdder FullAdder_1263 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1263_io_a),
    .io_b(FullAdder_1263_io_b),
    .io_ci(FullAdder_1263_io_ci),
    .io_s(FullAdder_1263_io_s),
    .io_co(FullAdder_1263_io_co)
  );
  FullAdder FullAdder_1264 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1264_io_a),
    .io_b(FullAdder_1264_io_b),
    .io_ci(FullAdder_1264_io_ci),
    .io_s(FullAdder_1264_io_s),
    .io_co(FullAdder_1264_io_co)
  );
  FullAdder FullAdder_1265 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1265_io_a),
    .io_b(FullAdder_1265_io_b),
    .io_ci(FullAdder_1265_io_ci),
    .io_s(FullAdder_1265_io_s),
    .io_co(FullAdder_1265_io_co)
  );
  HalfAdder HalfAdder_27 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_27_io_a),
    .io_b(HalfAdder_27_io_b),
    .io_s(HalfAdder_27_io_s),
    .io_co(HalfAdder_27_io_co)
  );
  FullAdder FullAdder_1266 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1266_io_a),
    .io_b(FullAdder_1266_io_b),
    .io_ci(FullAdder_1266_io_ci),
    .io_s(FullAdder_1266_io_s),
    .io_co(FullAdder_1266_io_co)
  );
  FullAdder FullAdder_1267 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1267_io_a),
    .io_b(FullAdder_1267_io_b),
    .io_ci(FullAdder_1267_io_ci),
    .io_s(FullAdder_1267_io_s),
    .io_co(FullAdder_1267_io_co)
  );
  FullAdder FullAdder_1268 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1268_io_a),
    .io_b(FullAdder_1268_io_b),
    .io_ci(FullAdder_1268_io_ci),
    .io_s(FullAdder_1268_io_s),
    .io_co(FullAdder_1268_io_co)
  );
  FullAdder FullAdder_1269 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1269_io_a),
    .io_b(FullAdder_1269_io_b),
    .io_ci(FullAdder_1269_io_ci),
    .io_s(FullAdder_1269_io_s),
    .io_co(FullAdder_1269_io_co)
  );
  FullAdder FullAdder_1270 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1270_io_a),
    .io_b(FullAdder_1270_io_b),
    .io_ci(FullAdder_1270_io_ci),
    .io_s(FullAdder_1270_io_s),
    .io_co(FullAdder_1270_io_co)
  );
  FullAdder FullAdder_1271 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1271_io_a),
    .io_b(FullAdder_1271_io_b),
    .io_ci(FullAdder_1271_io_ci),
    .io_s(FullAdder_1271_io_s),
    .io_co(FullAdder_1271_io_co)
  );
  FullAdder FullAdder_1272 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1272_io_a),
    .io_b(FullAdder_1272_io_b),
    .io_ci(FullAdder_1272_io_ci),
    .io_s(FullAdder_1272_io_s),
    .io_co(FullAdder_1272_io_co)
  );
  FullAdder FullAdder_1273 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1273_io_a),
    .io_b(FullAdder_1273_io_b),
    .io_ci(FullAdder_1273_io_ci),
    .io_s(FullAdder_1273_io_s),
    .io_co(FullAdder_1273_io_co)
  );
  FullAdder FullAdder_1274 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1274_io_a),
    .io_b(FullAdder_1274_io_b),
    .io_ci(FullAdder_1274_io_ci),
    .io_s(FullAdder_1274_io_s),
    .io_co(FullAdder_1274_io_co)
  );
  FullAdder FullAdder_1275 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1275_io_a),
    .io_b(FullAdder_1275_io_b),
    .io_ci(FullAdder_1275_io_ci),
    .io_s(FullAdder_1275_io_s),
    .io_co(FullAdder_1275_io_co)
  );
  FullAdder FullAdder_1276 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1276_io_a),
    .io_b(FullAdder_1276_io_b),
    .io_ci(FullAdder_1276_io_ci),
    .io_s(FullAdder_1276_io_s),
    .io_co(FullAdder_1276_io_co)
  );
  FullAdder FullAdder_1277 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1277_io_a),
    .io_b(FullAdder_1277_io_b),
    .io_ci(FullAdder_1277_io_ci),
    .io_s(FullAdder_1277_io_s),
    .io_co(FullAdder_1277_io_co)
  );
  FullAdder FullAdder_1278 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1278_io_a),
    .io_b(FullAdder_1278_io_b),
    .io_ci(FullAdder_1278_io_ci),
    .io_s(FullAdder_1278_io_s),
    .io_co(FullAdder_1278_io_co)
  );
  FullAdder FullAdder_1279 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1279_io_a),
    .io_b(FullAdder_1279_io_b),
    .io_ci(FullAdder_1279_io_ci),
    .io_s(FullAdder_1279_io_s),
    .io_co(FullAdder_1279_io_co)
  );
  FullAdder FullAdder_1280 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1280_io_a),
    .io_b(FullAdder_1280_io_b),
    .io_ci(FullAdder_1280_io_ci),
    .io_s(FullAdder_1280_io_s),
    .io_co(FullAdder_1280_io_co)
  );
  FullAdder FullAdder_1281 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1281_io_a),
    .io_b(FullAdder_1281_io_b),
    .io_ci(FullAdder_1281_io_ci),
    .io_s(FullAdder_1281_io_s),
    .io_co(FullAdder_1281_io_co)
  );
  FullAdder FullAdder_1282 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1282_io_a),
    .io_b(FullAdder_1282_io_b),
    .io_ci(FullAdder_1282_io_ci),
    .io_s(FullAdder_1282_io_s),
    .io_co(FullAdder_1282_io_co)
  );
  HalfAdder HalfAdder_28 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_28_io_a),
    .io_b(HalfAdder_28_io_b),
    .io_s(HalfAdder_28_io_s),
    .io_co(HalfAdder_28_io_co)
  );
  FullAdder FullAdder_1283 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1283_io_a),
    .io_b(FullAdder_1283_io_b),
    .io_ci(FullAdder_1283_io_ci),
    .io_s(FullAdder_1283_io_s),
    .io_co(FullAdder_1283_io_co)
  );
  FullAdder FullAdder_1284 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1284_io_a),
    .io_b(FullAdder_1284_io_b),
    .io_ci(FullAdder_1284_io_ci),
    .io_s(FullAdder_1284_io_s),
    .io_co(FullAdder_1284_io_co)
  );
  FullAdder FullAdder_1285 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1285_io_a),
    .io_b(FullAdder_1285_io_b),
    .io_ci(FullAdder_1285_io_ci),
    .io_s(FullAdder_1285_io_s),
    .io_co(FullAdder_1285_io_co)
  );
  FullAdder FullAdder_1286 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1286_io_a),
    .io_b(FullAdder_1286_io_b),
    .io_ci(FullAdder_1286_io_ci),
    .io_s(FullAdder_1286_io_s),
    .io_co(FullAdder_1286_io_co)
  );
  FullAdder FullAdder_1287 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1287_io_a),
    .io_b(FullAdder_1287_io_b),
    .io_ci(FullAdder_1287_io_ci),
    .io_s(FullAdder_1287_io_s),
    .io_co(FullAdder_1287_io_co)
  );
  FullAdder FullAdder_1288 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1288_io_a),
    .io_b(FullAdder_1288_io_b),
    .io_ci(FullAdder_1288_io_ci),
    .io_s(FullAdder_1288_io_s),
    .io_co(FullAdder_1288_io_co)
  );
  FullAdder FullAdder_1289 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1289_io_a),
    .io_b(FullAdder_1289_io_b),
    .io_ci(FullAdder_1289_io_ci),
    .io_s(FullAdder_1289_io_s),
    .io_co(FullAdder_1289_io_co)
  );
  FullAdder FullAdder_1290 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1290_io_a),
    .io_b(FullAdder_1290_io_b),
    .io_ci(FullAdder_1290_io_ci),
    .io_s(FullAdder_1290_io_s),
    .io_co(FullAdder_1290_io_co)
  );
  FullAdder FullAdder_1291 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1291_io_a),
    .io_b(FullAdder_1291_io_b),
    .io_ci(FullAdder_1291_io_ci),
    .io_s(FullAdder_1291_io_s),
    .io_co(FullAdder_1291_io_co)
  );
  FullAdder FullAdder_1292 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1292_io_a),
    .io_b(FullAdder_1292_io_b),
    .io_ci(FullAdder_1292_io_ci),
    .io_s(FullAdder_1292_io_s),
    .io_co(FullAdder_1292_io_co)
  );
  FullAdder FullAdder_1293 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1293_io_a),
    .io_b(FullAdder_1293_io_b),
    .io_ci(FullAdder_1293_io_ci),
    .io_s(FullAdder_1293_io_s),
    .io_co(FullAdder_1293_io_co)
  );
  FullAdder FullAdder_1294 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1294_io_a),
    .io_b(FullAdder_1294_io_b),
    .io_ci(FullAdder_1294_io_ci),
    .io_s(FullAdder_1294_io_s),
    .io_co(FullAdder_1294_io_co)
  );
  FullAdder FullAdder_1295 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1295_io_a),
    .io_b(FullAdder_1295_io_b),
    .io_ci(FullAdder_1295_io_ci),
    .io_s(FullAdder_1295_io_s),
    .io_co(FullAdder_1295_io_co)
  );
  FullAdder FullAdder_1296 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1296_io_a),
    .io_b(FullAdder_1296_io_b),
    .io_ci(FullAdder_1296_io_ci),
    .io_s(FullAdder_1296_io_s),
    .io_co(FullAdder_1296_io_co)
  );
  HalfAdder HalfAdder_29 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_29_io_a),
    .io_b(HalfAdder_29_io_b),
    .io_s(HalfAdder_29_io_s),
    .io_co(HalfAdder_29_io_co)
  );
  FullAdder FullAdder_1297 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1297_io_a),
    .io_b(FullAdder_1297_io_b),
    .io_ci(FullAdder_1297_io_ci),
    .io_s(FullAdder_1297_io_s),
    .io_co(FullAdder_1297_io_co)
  );
  FullAdder FullAdder_1298 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1298_io_a),
    .io_b(FullAdder_1298_io_b),
    .io_ci(FullAdder_1298_io_ci),
    .io_s(FullAdder_1298_io_s),
    .io_co(FullAdder_1298_io_co)
  );
  FullAdder FullAdder_1299 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1299_io_a),
    .io_b(FullAdder_1299_io_b),
    .io_ci(FullAdder_1299_io_ci),
    .io_s(FullAdder_1299_io_s),
    .io_co(FullAdder_1299_io_co)
  );
  FullAdder FullAdder_1300 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1300_io_a),
    .io_b(FullAdder_1300_io_b),
    .io_ci(FullAdder_1300_io_ci),
    .io_s(FullAdder_1300_io_s),
    .io_co(FullAdder_1300_io_co)
  );
  FullAdder FullAdder_1301 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1301_io_a),
    .io_b(FullAdder_1301_io_b),
    .io_ci(FullAdder_1301_io_ci),
    .io_s(FullAdder_1301_io_s),
    .io_co(FullAdder_1301_io_co)
  );
  FullAdder FullAdder_1302 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1302_io_a),
    .io_b(FullAdder_1302_io_b),
    .io_ci(FullAdder_1302_io_ci),
    .io_s(FullAdder_1302_io_s),
    .io_co(FullAdder_1302_io_co)
  );
  FullAdder FullAdder_1303 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1303_io_a),
    .io_b(FullAdder_1303_io_b),
    .io_ci(FullAdder_1303_io_ci),
    .io_s(FullAdder_1303_io_s),
    .io_co(FullAdder_1303_io_co)
  );
  FullAdder FullAdder_1304 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1304_io_a),
    .io_b(FullAdder_1304_io_b),
    .io_ci(FullAdder_1304_io_ci),
    .io_s(FullAdder_1304_io_s),
    .io_co(FullAdder_1304_io_co)
  );
  FullAdder FullAdder_1305 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1305_io_a),
    .io_b(FullAdder_1305_io_b),
    .io_ci(FullAdder_1305_io_ci),
    .io_s(FullAdder_1305_io_s),
    .io_co(FullAdder_1305_io_co)
  );
  FullAdder FullAdder_1306 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1306_io_a),
    .io_b(FullAdder_1306_io_b),
    .io_ci(FullAdder_1306_io_ci),
    .io_s(FullAdder_1306_io_s),
    .io_co(FullAdder_1306_io_co)
  );
  FullAdder FullAdder_1307 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1307_io_a),
    .io_b(FullAdder_1307_io_b),
    .io_ci(FullAdder_1307_io_ci),
    .io_s(FullAdder_1307_io_s),
    .io_co(FullAdder_1307_io_co)
  );
  HalfAdder HalfAdder_30 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_30_io_a),
    .io_b(HalfAdder_30_io_b),
    .io_s(HalfAdder_30_io_s),
    .io_co(HalfAdder_30_io_co)
  );
  FullAdder FullAdder_1308 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1308_io_a),
    .io_b(FullAdder_1308_io_b),
    .io_ci(FullAdder_1308_io_ci),
    .io_s(FullAdder_1308_io_s),
    .io_co(FullAdder_1308_io_co)
  );
  FullAdder FullAdder_1309 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1309_io_a),
    .io_b(FullAdder_1309_io_b),
    .io_ci(FullAdder_1309_io_ci),
    .io_s(FullAdder_1309_io_s),
    .io_co(FullAdder_1309_io_co)
  );
  FullAdder FullAdder_1310 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1310_io_a),
    .io_b(FullAdder_1310_io_b),
    .io_ci(FullAdder_1310_io_ci),
    .io_s(FullAdder_1310_io_s),
    .io_co(FullAdder_1310_io_co)
  );
  FullAdder FullAdder_1311 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1311_io_a),
    .io_b(FullAdder_1311_io_b),
    .io_ci(FullAdder_1311_io_ci),
    .io_s(FullAdder_1311_io_s),
    .io_co(FullAdder_1311_io_co)
  );
  FullAdder FullAdder_1312 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1312_io_a),
    .io_b(FullAdder_1312_io_b),
    .io_ci(FullAdder_1312_io_ci),
    .io_s(FullAdder_1312_io_s),
    .io_co(FullAdder_1312_io_co)
  );
  FullAdder FullAdder_1313 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1313_io_a),
    .io_b(FullAdder_1313_io_b),
    .io_ci(FullAdder_1313_io_ci),
    .io_s(FullAdder_1313_io_s),
    .io_co(FullAdder_1313_io_co)
  );
  FullAdder FullAdder_1314 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1314_io_a),
    .io_b(FullAdder_1314_io_b),
    .io_ci(FullAdder_1314_io_ci),
    .io_s(FullAdder_1314_io_s),
    .io_co(FullAdder_1314_io_co)
  );
  FullAdder FullAdder_1315 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1315_io_a),
    .io_b(FullAdder_1315_io_b),
    .io_ci(FullAdder_1315_io_ci),
    .io_s(FullAdder_1315_io_s),
    .io_co(FullAdder_1315_io_co)
  );
  HalfAdder HalfAdder_31 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_31_io_a),
    .io_b(HalfAdder_31_io_b),
    .io_s(HalfAdder_31_io_s),
    .io_co(HalfAdder_31_io_co)
  );
  FullAdder FullAdder_1316 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1316_io_a),
    .io_b(FullAdder_1316_io_b),
    .io_ci(FullAdder_1316_io_ci),
    .io_s(FullAdder_1316_io_s),
    .io_co(FullAdder_1316_io_co)
  );
  FullAdder FullAdder_1317 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1317_io_a),
    .io_b(FullAdder_1317_io_b),
    .io_ci(FullAdder_1317_io_ci),
    .io_s(FullAdder_1317_io_s),
    .io_co(FullAdder_1317_io_co)
  );
  FullAdder FullAdder_1318 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1318_io_a),
    .io_b(FullAdder_1318_io_b),
    .io_ci(FullAdder_1318_io_ci),
    .io_s(FullAdder_1318_io_s),
    .io_co(FullAdder_1318_io_co)
  );
  FullAdder FullAdder_1319 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1319_io_a),
    .io_b(FullAdder_1319_io_b),
    .io_ci(FullAdder_1319_io_ci),
    .io_s(FullAdder_1319_io_s),
    .io_co(FullAdder_1319_io_co)
  );
  FullAdder FullAdder_1320 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1320_io_a),
    .io_b(FullAdder_1320_io_b),
    .io_ci(FullAdder_1320_io_ci),
    .io_s(FullAdder_1320_io_s),
    .io_co(FullAdder_1320_io_co)
  );
  HalfAdder HalfAdder_32 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_32_io_a),
    .io_b(HalfAdder_32_io_b),
    .io_s(HalfAdder_32_io_s),
    .io_co(HalfAdder_32_io_co)
  );
  FullAdder FullAdder_1321 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1321_io_a),
    .io_b(FullAdder_1321_io_b),
    .io_ci(FullAdder_1321_io_ci),
    .io_s(FullAdder_1321_io_s),
    .io_co(FullAdder_1321_io_co)
  );
  HalfAdder HalfAdder_33 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_33_io_a),
    .io_b(HalfAdder_33_io_b),
    .io_s(HalfAdder_33_io_s),
    .io_co(HalfAdder_33_io_co)
  );
  HalfAdder HalfAdder_34 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_34_io_a),
    .io_b(HalfAdder_34_io_b),
    .io_s(HalfAdder_34_io_s),
    .io_co(HalfAdder_34_io_co)
  );
  HalfAdder HalfAdder_35 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_35_io_a),
    .io_b(HalfAdder_35_io_b),
    .io_s(HalfAdder_35_io_s),
    .io_co(HalfAdder_35_io_co)
  );
  HalfAdder HalfAdder_36 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_36_io_a),
    .io_b(HalfAdder_36_io_b),
    .io_s(HalfAdder_36_io_s),
    .io_co(HalfAdder_36_io_co)
  );
  FullAdder FullAdder_1322 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1322_io_a),
    .io_b(FullAdder_1322_io_b),
    .io_ci(FullAdder_1322_io_ci),
    .io_s(FullAdder_1322_io_s),
    .io_co(FullAdder_1322_io_co)
  );
  FullAdder FullAdder_1323 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1323_io_a),
    .io_b(FullAdder_1323_io_b),
    .io_ci(FullAdder_1323_io_ci),
    .io_s(FullAdder_1323_io_s),
    .io_co(FullAdder_1323_io_co)
  );
  FullAdder FullAdder_1324 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1324_io_a),
    .io_b(FullAdder_1324_io_b),
    .io_ci(FullAdder_1324_io_ci),
    .io_s(FullAdder_1324_io_s),
    .io_co(FullAdder_1324_io_co)
  );
  FullAdder FullAdder_1325 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1325_io_a),
    .io_b(FullAdder_1325_io_b),
    .io_ci(FullAdder_1325_io_ci),
    .io_s(FullAdder_1325_io_s),
    .io_co(FullAdder_1325_io_co)
  );
  FullAdder FullAdder_1326 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1326_io_a),
    .io_b(FullAdder_1326_io_b),
    .io_ci(FullAdder_1326_io_ci),
    .io_s(FullAdder_1326_io_s),
    .io_co(FullAdder_1326_io_co)
  );
  FullAdder FullAdder_1327 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1327_io_a),
    .io_b(FullAdder_1327_io_b),
    .io_ci(FullAdder_1327_io_ci),
    .io_s(FullAdder_1327_io_s),
    .io_co(FullAdder_1327_io_co)
  );
  FullAdder FullAdder_1328 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1328_io_a),
    .io_b(FullAdder_1328_io_b),
    .io_ci(FullAdder_1328_io_ci),
    .io_s(FullAdder_1328_io_s),
    .io_co(FullAdder_1328_io_co)
  );
  FullAdder FullAdder_1329 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1329_io_a),
    .io_b(FullAdder_1329_io_b),
    .io_ci(FullAdder_1329_io_ci),
    .io_s(FullAdder_1329_io_s),
    .io_co(FullAdder_1329_io_co)
  );
  FullAdder FullAdder_1330 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1330_io_a),
    .io_b(FullAdder_1330_io_b),
    .io_ci(FullAdder_1330_io_ci),
    .io_s(FullAdder_1330_io_s),
    .io_co(FullAdder_1330_io_co)
  );
  FullAdder FullAdder_1331 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1331_io_a),
    .io_b(FullAdder_1331_io_b),
    .io_ci(FullAdder_1331_io_ci),
    .io_s(FullAdder_1331_io_s),
    .io_co(FullAdder_1331_io_co)
  );
  FullAdder FullAdder_1332 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1332_io_a),
    .io_b(FullAdder_1332_io_b),
    .io_ci(FullAdder_1332_io_ci),
    .io_s(FullAdder_1332_io_s),
    .io_co(FullAdder_1332_io_co)
  );
  FullAdder FullAdder_1333 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1333_io_a),
    .io_b(FullAdder_1333_io_b),
    .io_ci(FullAdder_1333_io_ci),
    .io_s(FullAdder_1333_io_s),
    .io_co(FullAdder_1333_io_co)
  );
  FullAdder FullAdder_1334 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1334_io_a),
    .io_b(FullAdder_1334_io_b),
    .io_ci(FullAdder_1334_io_ci),
    .io_s(FullAdder_1334_io_s),
    .io_co(FullAdder_1334_io_co)
  );
  HalfAdder HalfAdder_37 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_37_io_a),
    .io_b(HalfAdder_37_io_b),
    .io_s(HalfAdder_37_io_s),
    .io_co(HalfAdder_37_io_co)
  );
  FullAdder FullAdder_1335 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1335_io_a),
    .io_b(FullAdder_1335_io_b),
    .io_ci(FullAdder_1335_io_ci),
    .io_s(FullAdder_1335_io_s),
    .io_co(FullAdder_1335_io_co)
  );
  FullAdder FullAdder_1336 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1336_io_a),
    .io_b(FullAdder_1336_io_b),
    .io_ci(FullAdder_1336_io_ci),
    .io_s(FullAdder_1336_io_s),
    .io_co(FullAdder_1336_io_co)
  );
  HalfAdder HalfAdder_38 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_38_io_a),
    .io_b(HalfAdder_38_io_b),
    .io_s(HalfAdder_38_io_s),
    .io_co(HalfAdder_38_io_co)
  );
  FullAdder FullAdder_1337 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1337_io_a),
    .io_b(FullAdder_1337_io_b),
    .io_ci(FullAdder_1337_io_ci),
    .io_s(FullAdder_1337_io_s),
    .io_co(FullAdder_1337_io_co)
  );
  FullAdder FullAdder_1338 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1338_io_a),
    .io_b(FullAdder_1338_io_b),
    .io_ci(FullAdder_1338_io_ci),
    .io_s(FullAdder_1338_io_s),
    .io_co(FullAdder_1338_io_co)
  );
  FullAdder FullAdder_1339 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1339_io_a),
    .io_b(FullAdder_1339_io_b),
    .io_ci(FullAdder_1339_io_ci),
    .io_s(FullAdder_1339_io_s),
    .io_co(FullAdder_1339_io_co)
  );
  FullAdder FullAdder_1340 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1340_io_a),
    .io_b(FullAdder_1340_io_b),
    .io_ci(FullAdder_1340_io_ci),
    .io_s(FullAdder_1340_io_s),
    .io_co(FullAdder_1340_io_co)
  );
  FullAdder FullAdder_1341 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1341_io_a),
    .io_b(FullAdder_1341_io_b),
    .io_ci(FullAdder_1341_io_ci),
    .io_s(FullAdder_1341_io_s),
    .io_co(FullAdder_1341_io_co)
  );
  FullAdder FullAdder_1342 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1342_io_a),
    .io_b(FullAdder_1342_io_b),
    .io_ci(FullAdder_1342_io_ci),
    .io_s(FullAdder_1342_io_s),
    .io_co(FullAdder_1342_io_co)
  );
  FullAdder FullAdder_1343 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1343_io_a),
    .io_b(FullAdder_1343_io_b),
    .io_ci(FullAdder_1343_io_ci),
    .io_s(FullAdder_1343_io_s),
    .io_co(FullAdder_1343_io_co)
  );
  FullAdder FullAdder_1344 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1344_io_a),
    .io_b(FullAdder_1344_io_b),
    .io_ci(FullAdder_1344_io_ci),
    .io_s(FullAdder_1344_io_s),
    .io_co(FullAdder_1344_io_co)
  );
  FullAdder FullAdder_1345 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1345_io_a),
    .io_b(FullAdder_1345_io_b),
    .io_ci(FullAdder_1345_io_ci),
    .io_s(FullAdder_1345_io_s),
    .io_co(FullAdder_1345_io_co)
  );
  FullAdder FullAdder_1346 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1346_io_a),
    .io_b(FullAdder_1346_io_b),
    .io_ci(FullAdder_1346_io_ci),
    .io_s(FullAdder_1346_io_s),
    .io_co(FullAdder_1346_io_co)
  );
  FullAdder FullAdder_1347 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1347_io_a),
    .io_b(FullAdder_1347_io_b),
    .io_ci(FullAdder_1347_io_ci),
    .io_s(FullAdder_1347_io_s),
    .io_co(FullAdder_1347_io_co)
  );
  FullAdder FullAdder_1348 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1348_io_a),
    .io_b(FullAdder_1348_io_b),
    .io_ci(FullAdder_1348_io_ci),
    .io_s(FullAdder_1348_io_s),
    .io_co(FullAdder_1348_io_co)
  );
  FullAdder FullAdder_1349 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1349_io_a),
    .io_b(FullAdder_1349_io_b),
    .io_ci(FullAdder_1349_io_ci),
    .io_s(FullAdder_1349_io_s),
    .io_co(FullAdder_1349_io_co)
  );
  FullAdder FullAdder_1350 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1350_io_a),
    .io_b(FullAdder_1350_io_b),
    .io_ci(FullAdder_1350_io_ci),
    .io_s(FullAdder_1350_io_s),
    .io_co(FullAdder_1350_io_co)
  );
  FullAdder FullAdder_1351 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1351_io_a),
    .io_b(FullAdder_1351_io_b),
    .io_ci(FullAdder_1351_io_ci),
    .io_s(FullAdder_1351_io_s),
    .io_co(FullAdder_1351_io_co)
  );
  FullAdder FullAdder_1352 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1352_io_a),
    .io_b(FullAdder_1352_io_b),
    .io_ci(FullAdder_1352_io_ci),
    .io_s(FullAdder_1352_io_s),
    .io_co(FullAdder_1352_io_co)
  );
  FullAdder FullAdder_1353 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1353_io_a),
    .io_b(FullAdder_1353_io_b),
    .io_ci(FullAdder_1353_io_ci),
    .io_s(FullAdder_1353_io_s),
    .io_co(FullAdder_1353_io_co)
  );
  FullAdder FullAdder_1354 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1354_io_a),
    .io_b(FullAdder_1354_io_b),
    .io_ci(FullAdder_1354_io_ci),
    .io_s(FullAdder_1354_io_s),
    .io_co(FullAdder_1354_io_co)
  );
  FullAdder FullAdder_1355 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1355_io_a),
    .io_b(FullAdder_1355_io_b),
    .io_ci(FullAdder_1355_io_ci),
    .io_s(FullAdder_1355_io_s),
    .io_co(FullAdder_1355_io_co)
  );
  FullAdder FullAdder_1356 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1356_io_a),
    .io_b(FullAdder_1356_io_b),
    .io_ci(FullAdder_1356_io_ci),
    .io_s(FullAdder_1356_io_s),
    .io_co(FullAdder_1356_io_co)
  );
  FullAdder FullAdder_1357 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1357_io_a),
    .io_b(FullAdder_1357_io_b),
    .io_ci(FullAdder_1357_io_ci),
    .io_s(FullAdder_1357_io_s),
    .io_co(FullAdder_1357_io_co)
  );
  FullAdder FullAdder_1358 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1358_io_a),
    .io_b(FullAdder_1358_io_b),
    .io_ci(FullAdder_1358_io_ci),
    .io_s(FullAdder_1358_io_s),
    .io_co(FullAdder_1358_io_co)
  );
  FullAdder FullAdder_1359 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1359_io_a),
    .io_b(FullAdder_1359_io_b),
    .io_ci(FullAdder_1359_io_ci),
    .io_s(FullAdder_1359_io_s),
    .io_co(FullAdder_1359_io_co)
  );
  FullAdder FullAdder_1360 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1360_io_a),
    .io_b(FullAdder_1360_io_b),
    .io_ci(FullAdder_1360_io_ci),
    .io_s(FullAdder_1360_io_s),
    .io_co(FullAdder_1360_io_co)
  );
  FullAdder FullAdder_1361 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1361_io_a),
    .io_b(FullAdder_1361_io_b),
    .io_ci(FullAdder_1361_io_ci),
    .io_s(FullAdder_1361_io_s),
    .io_co(FullAdder_1361_io_co)
  );
  HalfAdder HalfAdder_39 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_39_io_a),
    .io_b(HalfAdder_39_io_b),
    .io_s(HalfAdder_39_io_s),
    .io_co(HalfAdder_39_io_co)
  );
  FullAdder FullAdder_1362 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1362_io_a),
    .io_b(FullAdder_1362_io_b),
    .io_ci(FullAdder_1362_io_ci),
    .io_s(FullAdder_1362_io_s),
    .io_co(FullAdder_1362_io_co)
  );
  FullAdder FullAdder_1363 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1363_io_a),
    .io_b(FullAdder_1363_io_b),
    .io_ci(FullAdder_1363_io_ci),
    .io_s(FullAdder_1363_io_s),
    .io_co(FullAdder_1363_io_co)
  );
  FullAdder FullAdder_1364 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1364_io_a),
    .io_b(FullAdder_1364_io_b),
    .io_ci(FullAdder_1364_io_ci),
    .io_s(FullAdder_1364_io_s),
    .io_co(FullAdder_1364_io_co)
  );
  FullAdder FullAdder_1365 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1365_io_a),
    .io_b(FullAdder_1365_io_b),
    .io_ci(FullAdder_1365_io_ci),
    .io_s(FullAdder_1365_io_s),
    .io_co(FullAdder_1365_io_co)
  );
  HalfAdder HalfAdder_40 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_40_io_a),
    .io_b(HalfAdder_40_io_b),
    .io_s(HalfAdder_40_io_s),
    .io_co(HalfAdder_40_io_co)
  );
  FullAdder FullAdder_1366 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1366_io_a),
    .io_b(FullAdder_1366_io_b),
    .io_ci(FullAdder_1366_io_ci),
    .io_s(FullAdder_1366_io_s),
    .io_co(FullAdder_1366_io_co)
  );
  FullAdder FullAdder_1367 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1367_io_a),
    .io_b(FullAdder_1367_io_b),
    .io_ci(FullAdder_1367_io_ci),
    .io_s(FullAdder_1367_io_s),
    .io_co(FullAdder_1367_io_co)
  );
  FullAdder FullAdder_1368 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1368_io_a),
    .io_b(FullAdder_1368_io_b),
    .io_ci(FullAdder_1368_io_ci),
    .io_s(FullAdder_1368_io_s),
    .io_co(FullAdder_1368_io_co)
  );
  FullAdder FullAdder_1369 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1369_io_a),
    .io_b(FullAdder_1369_io_b),
    .io_ci(FullAdder_1369_io_ci),
    .io_s(FullAdder_1369_io_s),
    .io_co(FullAdder_1369_io_co)
  );
  HalfAdder HalfAdder_41 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_41_io_a),
    .io_b(HalfAdder_41_io_b),
    .io_s(HalfAdder_41_io_s),
    .io_co(HalfAdder_41_io_co)
  );
  FullAdder FullAdder_1370 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1370_io_a),
    .io_b(FullAdder_1370_io_b),
    .io_ci(FullAdder_1370_io_ci),
    .io_s(FullAdder_1370_io_s),
    .io_co(FullAdder_1370_io_co)
  );
  FullAdder FullAdder_1371 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1371_io_a),
    .io_b(FullAdder_1371_io_b),
    .io_ci(FullAdder_1371_io_ci),
    .io_s(FullAdder_1371_io_s),
    .io_co(FullAdder_1371_io_co)
  );
  FullAdder FullAdder_1372 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1372_io_a),
    .io_b(FullAdder_1372_io_b),
    .io_ci(FullAdder_1372_io_ci),
    .io_s(FullAdder_1372_io_s),
    .io_co(FullAdder_1372_io_co)
  );
  FullAdder FullAdder_1373 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1373_io_a),
    .io_b(FullAdder_1373_io_b),
    .io_ci(FullAdder_1373_io_ci),
    .io_s(FullAdder_1373_io_s),
    .io_co(FullAdder_1373_io_co)
  );
  FullAdder FullAdder_1374 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1374_io_a),
    .io_b(FullAdder_1374_io_b),
    .io_ci(FullAdder_1374_io_ci),
    .io_s(FullAdder_1374_io_s),
    .io_co(FullAdder_1374_io_co)
  );
  FullAdder FullAdder_1375 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1375_io_a),
    .io_b(FullAdder_1375_io_b),
    .io_ci(FullAdder_1375_io_ci),
    .io_s(FullAdder_1375_io_s),
    .io_co(FullAdder_1375_io_co)
  );
  FullAdder FullAdder_1376 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1376_io_a),
    .io_b(FullAdder_1376_io_b),
    .io_ci(FullAdder_1376_io_ci),
    .io_s(FullAdder_1376_io_s),
    .io_co(FullAdder_1376_io_co)
  );
  FullAdder FullAdder_1377 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1377_io_a),
    .io_b(FullAdder_1377_io_b),
    .io_ci(FullAdder_1377_io_ci),
    .io_s(FullAdder_1377_io_s),
    .io_co(FullAdder_1377_io_co)
  );
  FullAdder FullAdder_1378 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1378_io_a),
    .io_b(FullAdder_1378_io_b),
    .io_ci(FullAdder_1378_io_ci),
    .io_s(FullAdder_1378_io_s),
    .io_co(FullAdder_1378_io_co)
  );
  FullAdder FullAdder_1379 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1379_io_a),
    .io_b(FullAdder_1379_io_b),
    .io_ci(FullAdder_1379_io_ci),
    .io_s(FullAdder_1379_io_s),
    .io_co(FullAdder_1379_io_co)
  );
  FullAdder FullAdder_1380 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1380_io_a),
    .io_b(FullAdder_1380_io_b),
    .io_ci(FullAdder_1380_io_ci),
    .io_s(FullAdder_1380_io_s),
    .io_co(FullAdder_1380_io_co)
  );
  FullAdder FullAdder_1381 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1381_io_a),
    .io_b(FullAdder_1381_io_b),
    .io_ci(FullAdder_1381_io_ci),
    .io_s(FullAdder_1381_io_s),
    .io_co(FullAdder_1381_io_co)
  );
  FullAdder FullAdder_1382 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1382_io_a),
    .io_b(FullAdder_1382_io_b),
    .io_ci(FullAdder_1382_io_ci),
    .io_s(FullAdder_1382_io_s),
    .io_co(FullAdder_1382_io_co)
  );
  FullAdder FullAdder_1383 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1383_io_a),
    .io_b(FullAdder_1383_io_b),
    .io_ci(FullAdder_1383_io_ci),
    .io_s(FullAdder_1383_io_s),
    .io_co(FullAdder_1383_io_co)
  );
  FullAdder FullAdder_1384 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1384_io_a),
    .io_b(FullAdder_1384_io_b),
    .io_ci(FullAdder_1384_io_ci),
    .io_s(FullAdder_1384_io_s),
    .io_co(FullAdder_1384_io_co)
  );
  FullAdder FullAdder_1385 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1385_io_a),
    .io_b(FullAdder_1385_io_b),
    .io_ci(FullAdder_1385_io_ci),
    .io_s(FullAdder_1385_io_s),
    .io_co(FullAdder_1385_io_co)
  );
  FullAdder FullAdder_1386 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1386_io_a),
    .io_b(FullAdder_1386_io_b),
    .io_ci(FullAdder_1386_io_ci),
    .io_s(FullAdder_1386_io_s),
    .io_co(FullAdder_1386_io_co)
  );
  FullAdder FullAdder_1387 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1387_io_a),
    .io_b(FullAdder_1387_io_b),
    .io_ci(FullAdder_1387_io_ci),
    .io_s(FullAdder_1387_io_s),
    .io_co(FullAdder_1387_io_co)
  );
  FullAdder FullAdder_1388 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1388_io_a),
    .io_b(FullAdder_1388_io_b),
    .io_ci(FullAdder_1388_io_ci),
    .io_s(FullAdder_1388_io_s),
    .io_co(FullAdder_1388_io_co)
  );
  FullAdder FullAdder_1389 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1389_io_a),
    .io_b(FullAdder_1389_io_b),
    .io_ci(FullAdder_1389_io_ci),
    .io_s(FullAdder_1389_io_s),
    .io_co(FullAdder_1389_io_co)
  );
  FullAdder FullAdder_1390 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1390_io_a),
    .io_b(FullAdder_1390_io_b),
    .io_ci(FullAdder_1390_io_ci),
    .io_s(FullAdder_1390_io_s),
    .io_co(FullAdder_1390_io_co)
  );
  FullAdder FullAdder_1391 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1391_io_a),
    .io_b(FullAdder_1391_io_b),
    .io_ci(FullAdder_1391_io_ci),
    .io_s(FullAdder_1391_io_s),
    .io_co(FullAdder_1391_io_co)
  );
  FullAdder FullAdder_1392 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1392_io_a),
    .io_b(FullAdder_1392_io_b),
    .io_ci(FullAdder_1392_io_ci),
    .io_s(FullAdder_1392_io_s),
    .io_co(FullAdder_1392_io_co)
  );
  FullAdder FullAdder_1393 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1393_io_a),
    .io_b(FullAdder_1393_io_b),
    .io_ci(FullAdder_1393_io_ci),
    .io_s(FullAdder_1393_io_s),
    .io_co(FullAdder_1393_io_co)
  );
  FullAdder FullAdder_1394 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1394_io_a),
    .io_b(FullAdder_1394_io_b),
    .io_ci(FullAdder_1394_io_ci),
    .io_s(FullAdder_1394_io_s),
    .io_co(FullAdder_1394_io_co)
  );
  FullAdder FullAdder_1395 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1395_io_a),
    .io_b(FullAdder_1395_io_b),
    .io_ci(FullAdder_1395_io_ci),
    .io_s(FullAdder_1395_io_s),
    .io_co(FullAdder_1395_io_co)
  );
  FullAdder FullAdder_1396 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1396_io_a),
    .io_b(FullAdder_1396_io_b),
    .io_ci(FullAdder_1396_io_ci),
    .io_s(FullAdder_1396_io_s),
    .io_co(FullAdder_1396_io_co)
  );
  FullAdder FullAdder_1397 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1397_io_a),
    .io_b(FullAdder_1397_io_b),
    .io_ci(FullAdder_1397_io_ci),
    .io_s(FullAdder_1397_io_s),
    .io_co(FullAdder_1397_io_co)
  );
  FullAdder FullAdder_1398 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1398_io_a),
    .io_b(FullAdder_1398_io_b),
    .io_ci(FullAdder_1398_io_ci),
    .io_s(FullAdder_1398_io_s),
    .io_co(FullAdder_1398_io_co)
  );
  FullAdder FullAdder_1399 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1399_io_a),
    .io_b(FullAdder_1399_io_b),
    .io_ci(FullAdder_1399_io_ci),
    .io_s(FullAdder_1399_io_s),
    .io_co(FullAdder_1399_io_co)
  );
  FullAdder FullAdder_1400 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1400_io_a),
    .io_b(FullAdder_1400_io_b),
    .io_ci(FullAdder_1400_io_ci),
    .io_s(FullAdder_1400_io_s),
    .io_co(FullAdder_1400_io_co)
  );
  FullAdder FullAdder_1401 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1401_io_a),
    .io_b(FullAdder_1401_io_b),
    .io_ci(FullAdder_1401_io_ci),
    .io_s(FullAdder_1401_io_s),
    .io_co(FullAdder_1401_io_co)
  );
  FullAdder FullAdder_1402 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1402_io_a),
    .io_b(FullAdder_1402_io_b),
    .io_ci(FullAdder_1402_io_ci),
    .io_s(FullAdder_1402_io_s),
    .io_co(FullAdder_1402_io_co)
  );
  FullAdder FullAdder_1403 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1403_io_a),
    .io_b(FullAdder_1403_io_b),
    .io_ci(FullAdder_1403_io_ci),
    .io_s(FullAdder_1403_io_s),
    .io_co(FullAdder_1403_io_co)
  );
  FullAdder FullAdder_1404 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1404_io_a),
    .io_b(FullAdder_1404_io_b),
    .io_ci(FullAdder_1404_io_ci),
    .io_s(FullAdder_1404_io_s),
    .io_co(FullAdder_1404_io_co)
  );
  FullAdder FullAdder_1405 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1405_io_a),
    .io_b(FullAdder_1405_io_b),
    .io_ci(FullAdder_1405_io_ci),
    .io_s(FullAdder_1405_io_s),
    .io_co(FullAdder_1405_io_co)
  );
  FullAdder FullAdder_1406 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1406_io_a),
    .io_b(FullAdder_1406_io_b),
    .io_ci(FullAdder_1406_io_ci),
    .io_s(FullAdder_1406_io_s),
    .io_co(FullAdder_1406_io_co)
  );
  FullAdder FullAdder_1407 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1407_io_a),
    .io_b(FullAdder_1407_io_b),
    .io_ci(FullAdder_1407_io_ci),
    .io_s(FullAdder_1407_io_s),
    .io_co(FullAdder_1407_io_co)
  );
  FullAdder FullAdder_1408 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1408_io_a),
    .io_b(FullAdder_1408_io_b),
    .io_ci(FullAdder_1408_io_ci),
    .io_s(FullAdder_1408_io_s),
    .io_co(FullAdder_1408_io_co)
  );
  FullAdder FullAdder_1409 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1409_io_a),
    .io_b(FullAdder_1409_io_b),
    .io_ci(FullAdder_1409_io_ci),
    .io_s(FullAdder_1409_io_s),
    .io_co(FullAdder_1409_io_co)
  );
  FullAdder FullAdder_1410 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1410_io_a),
    .io_b(FullAdder_1410_io_b),
    .io_ci(FullAdder_1410_io_ci),
    .io_s(FullAdder_1410_io_s),
    .io_co(FullAdder_1410_io_co)
  );
  FullAdder FullAdder_1411 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1411_io_a),
    .io_b(FullAdder_1411_io_b),
    .io_ci(FullAdder_1411_io_ci),
    .io_s(FullAdder_1411_io_s),
    .io_co(FullAdder_1411_io_co)
  );
  FullAdder FullAdder_1412 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1412_io_a),
    .io_b(FullAdder_1412_io_b),
    .io_ci(FullAdder_1412_io_ci),
    .io_s(FullAdder_1412_io_s),
    .io_co(FullAdder_1412_io_co)
  );
  FullAdder FullAdder_1413 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1413_io_a),
    .io_b(FullAdder_1413_io_b),
    .io_ci(FullAdder_1413_io_ci),
    .io_s(FullAdder_1413_io_s),
    .io_co(FullAdder_1413_io_co)
  );
  FullAdder FullAdder_1414 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1414_io_a),
    .io_b(FullAdder_1414_io_b),
    .io_ci(FullAdder_1414_io_ci),
    .io_s(FullAdder_1414_io_s),
    .io_co(FullAdder_1414_io_co)
  );
  FullAdder FullAdder_1415 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1415_io_a),
    .io_b(FullAdder_1415_io_b),
    .io_ci(FullAdder_1415_io_ci),
    .io_s(FullAdder_1415_io_s),
    .io_co(FullAdder_1415_io_co)
  );
  FullAdder FullAdder_1416 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1416_io_a),
    .io_b(FullAdder_1416_io_b),
    .io_ci(FullAdder_1416_io_ci),
    .io_s(FullAdder_1416_io_s),
    .io_co(FullAdder_1416_io_co)
  );
  FullAdder FullAdder_1417 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1417_io_a),
    .io_b(FullAdder_1417_io_b),
    .io_ci(FullAdder_1417_io_ci),
    .io_s(FullAdder_1417_io_s),
    .io_co(FullAdder_1417_io_co)
  );
  FullAdder FullAdder_1418 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1418_io_a),
    .io_b(FullAdder_1418_io_b),
    .io_ci(FullAdder_1418_io_ci),
    .io_s(FullAdder_1418_io_s),
    .io_co(FullAdder_1418_io_co)
  );
  FullAdder FullAdder_1419 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1419_io_a),
    .io_b(FullAdder_1419_io_b),
    .io_ci(FullAdder_1419_io_ci),
    .io_s(FullAdder_1419_io_s),
    .io_co(FullAdder_1419_io_co)
  );
  FullAdder FullAdder_1420 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1420_io_a),
    .io_b(FullAdder_1420_io_b),
    .io_ci(FullAdder_1420_io_ci),
    .io_s(FullAdder_1420_io_s),
    .io_co(FullAdder_1420_io_co)
  );
  HalfAdder HalfAdder_42 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_42_io_a),
    .io_b(HalfAdder_42_io_b),
    .io_s(HalfAdder_42_io_s),
    .io_co(HalfAdder_42_io_co)
  );
  FullAdder FullAdder_1421 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1421_io_a),
    .io_b(FullAdder_1421_io_b),
    .io_ci(FullAdder_1421_io_ci),
    .io_s(FullAdder_1421_io_s),
    .io_co(FullAdder_1421_io_co)
  );
  FullAdder FullAdder_1422 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1422_io_a),
    .io_b(FullAdder_1422_io_b),
    .io_ci(FullAdder_1422_io_ci),
    .io_s(FullAdder_1422_io_s),
    .io_co(FullAdder_1422_io_co)
  );
  FullAdder FullAdder_1423 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1423_io_a),
    .io_b(FullAdder_1423_io_b),
    .io_ci(FullAdder_1423_io_ci),
    .io_s(FullAdder_1423_io_s),
    .io_co(FullAdder_1423_io_co)
  );
  FullAdder FullAdder_1424 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1424_io_a),
    .io_b(FullAdder_1424_io_b),
    .io_ci(FullAdder_1424_io_ci),
    .io_s(FullAdder_1424_io_s),
    .io_co(FullAdder_1424_io_co)
  );
  FullAdder FullAdder_1425 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1425_io_a),
    .io_b(FullAdder_1425_io_b),
    .io_ci(FullAdder_1425_io_ci),
    .io_s(FullAdder_1425_io_s),
    .io_co(FullAdder_1425_io_co)
  );
  FullAdder FullAdder_1426 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1426_io_a),
    .io_b(FullAdder_1426_io_b),
    .io_ci(FullAdder_1426_io_ci),
    .io_s(FullAdder_1426_io_s),
    .io_co(FullAdder_1426_io_co)
  );
  FullAdder FullAdder_1427 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1427_io_a),
    .io_b(FullAdder_1427_io_b),
    .io_ci(FullAdder_1427_io_ci),
    .io_s(FullAdder_1427_io_s),
    .io_co(FullAdder_1427_io_co)
  );
  FullAdder FullAdder_1428 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1428_io_a),
    .io_b(FullAdder_1428_io_b),
    .io_ci(FullAdder_1428_io_ci),
    .io_s(FullAdder_1428_io_s),
    .io_co(FullAdder_1428_io_co)
  );
  FullAdder FullAdder_1429 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1429_io_a),
    .io_b(FullAdder_1429_io_b),
    .io_ci(FullAdder_1429_io_ci),
    .io_s(FullAdder_1429_io_s),
    .io_co(FullAdder_1429_io_co)
  );
  FullAdder FullAdder_1430 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1430_io_a),
    .io_b(FullAdder_1430_io_b),
    .io_ci(FullAdder_1430_io_ci),
    .io_s(FullAdder_1430_io_s),
    .io_co(FullAdder_1430_io_co)
  );
  FullAdder FullAdder_1431 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1431_io_a),
    .io_b(FullAdder_1431_io_b),
    .io_ci(FullAdder_1431_io_ci),
    .io_s(FullAdder_1431_io_s),
    .io_co(FullAdder_1431_io_co)
  );
  FullAdder FullAdder_1432 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1432_io_a),
    .io_b(FullAdder_1432_io_b),
    .io_ci(FullAdder_1432_io_ci),
    .io_s(FullAdder_1432_io_s),
    .io_co(FullAdder_1432_io_co)
  );
  FullAdder FullAdder_1433 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1433_io_a),
    .io_b(FullAdder_1433_io_b),
    .io_ci(FullAdder_1433_io_ci),
    .io_s(FullAdder_1433_io_s),
    .io_co(FullAdder_1433_io_co)
  );
  FullAdder FullAdder_1434 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1434_io_a),
    .io_b(FullAdder_1434_io_b),
    .io_ci(FullAdder_1434_io_ci),
    .io_s(FullAdder_1434_io_s),
    .io_co(FullAdder_1434_io_co)
  );
  FullAdder FullAdder_1435 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1435_io_a),
    .io_b(FullAdder_1435_io_b),
    .io_ci(FullAdder_1435_io_ci),
    .io_s(FullAdder_1435_io_s),
    .io_co(FullAdder_1435_io_co)
  );
  FullAdder FullAdder_1436 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1436_io_a),
    .io_b(FullAdder_1436_io_b),
    .io_ci(FullAdder_1436_io_ci),
    .io_s(FullAdder_1436_io_s),
    .io_co(FullAdder_1436_io_co)
  );
  FullAdder FullAdder_1437 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1437_io_a),
    .io_b(FullAdder_1437_io_b),
    .io_ci(FullAdder_1437_io_ci),
    .io_s(FullAdder_1437_io_s),
    .io_co(FullAdder_1437_io_co)
  );
  FullAdder FullAdder_1438 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1438_io_a),
    .io_b(FullAdder_1438_io_b),
    .io_ci(FullAdder_1438_io_ci),
    .io_s(FullAdder_1438_io_s),
    .io_co(FullAdder_1438_io_co)
  );
  FullAdder FullAdder_1439 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1439_io_a),
    .io_b(FullAdder_1439_io_b),
    .io_ci(FullAdder_1439_io_ci),
    .io_s(FullAdder_1439_io_s),
    .io_co(FullAdder_1439_io_co)
  );
  FullAdder FullAdder_1440 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1440_io_a),
    .io_b(FullAdder_1440_io_b),
    .io_ci(FullAdder_1440_io_ci),
    .io_s(FullAdder_1440_io_s),
    .io_co(FullAdder_1440_io_co)
  );
  FullAdder FullAdder_1441 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1441_io_a),
    .io_b(FullAdder_1441_io_b),
    .io_ci(FullAdder_1441_io_ci),
    .io_s(FullAdder_1441_io_s),
    .io_co(FullAdder_1441_io_co)
  );
  FullAdder FullAdder_1442 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1442_io_a),
    .io_b(FullAdder_1442_io_b),
    .io_ci(FullAdder_1442_io_ci),
    .io_s(FullAdder_1442_io_s),
    .io_co(FullAdder_1442_io_co)
  );
  FullAdder FullAdder_1443 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1443_io_a),
    .io_b(FullAdder_1443_io_b),
    .io_ci(FullAdder_1443_io_ci),
    .io_s(FullAdder_1443_io_s),
    .io_co(FullAdder_1443_io_co)
  );
  FullAdder FullAdder_1444 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1444_io_a),
    .io_b(FullAdder_1444_io_b),
    .io_ci(FullAdder_1444_io_ci),
    .io_s(FullAdder_1444_io_s),
    .io_co(FullAdder_1444_io_co)
  );
  FullAdder FullAdder_1445 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1445_io_a),
    .io_b(FullAdder_1445_io_b),
    .io_ci(FullAdder_1445_io_ci),
    .io_s(FullAdder_1445_io_s),
    .io_co(FullAdder_1445_io_co)
  );
  FullAdder FullAdder_1446 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1446_io_a),
    .io_b(FullAdder_1446_io_b),
    .io_ci(FullAdder_1446_io_ci),
    .io_s(FullAdder_1446_io_s),
    .io_co(FullAdder_1446_io_co)
  );
  FullAdder FullAdder_1447 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1447_io_a),
    .io_b(FullAdder_1447_io_b),
    .io_ci(FullAdder_1447_io_ci),
    .io_s(FullAdder_1447_io_s),
    .io_co(FullAdder_1447_io_co)
  );
  FullAdder FullAdder_1448 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1448_io_a),
    .io_b(FullAdder_1448_io_b),
    .io_ci(FullAdder_1448_io_ci),
    .io_s(FullAdder_1448_io_s),
    .io_co(FullAdder_1448_io_co)
  );
  FullAdder FullAdder_1449 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1449_io_a),
    .io_b(FullAdder_1449_io_b),
    .io_ci(FullAdder_1449_io_ci),
    .io_s(FullAdder_1449_io_s),
    .io_co(FullAdder_1449_io_co)
  );
  FullAdder FullAdder_1450 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1450_io_a),
    .io_b(FullAdder_1450_io_b),
    .io_ci(FullAdder_1450_io_ci),
    .io_s(FullAdder_1450_io_s),
    .io_co(FullAdder_1450_io_co)
  );
  FullAdder FullAdder_1451 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1451_io_a),
    .io_b(FullAdder_1451_io_b),
    .io_ci(FullAdder_1451_io_ci),
    .io_s(FullAdder_1451_io_s),
    .io_co(FullAdder_1451_io_co)
  );
  FullAdder FullAdder_1452 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1452_io_a),
    .io_b(FullAdder_1452_io_b),
    .io_ci(FullAdder_1452_io_ci),
    .io_s(FullAdder_1452_io_s),
    .io_co(FullAdder_1452_io_co)
  );
  FullAdder FullAdder_1453 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1453_io_a),
    .io_b(FullAdder_1453_io_b),
    .io_ci(FullAdder_1453_io_ci),
    .io_s(FullAdder_1453_io_s),
    .io_co(FullAdder_1453_io_co)
  );
  FullAdder FullAdder_1454 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1454_io_a),
    .io_b(FullAdder_1454_io_b),
    .io_ci(FullAdder_1454_io_ci),
    .io_s(FullAdder_1454_io_s),
    .io_co(FullAdder_1454_io_co)
  );
  FullAdder FullAdder_1455 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1455_io_a),
    .io_b(FullAdder_1455_io_b),
    .io_ci(FullAdder_1455_io_ci),
    .io_s(FullAdder_1455_io_s),
    .io_co(FullAdder_1455_io_co)
  );
  FullAdder FullAdder_1456 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1456_io_a),
    .io_b(FullAdder_1456_io_b),
    .io_ci(FullAdder_1456_io_ci),
    .io_s(FullAdder_1456_io_s),
    .io_co(FullAdder_1456_io_co)
  );
  FullAdder FullAdder_1457 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1457_io_a),
    .io_b(FullAdder_1457_io_b),
    .io_ci(FullAdder_1457_io_ci),
    .io_s(FullAdder_1457_io_s),
    .io_co(FullAdder_1457_io_co)
  );
  FullAdder FullAdder_1458 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1458_io_a),
    .io_b(FullAdder_1458_io_b),
    .io_ci(FullAdder_1458_io_ci),
    .io_s(FullAdder_1458_io_s),
    .io_co(FullAdder_1458_io_co)
  );
  FullAdder FullAdder_1459 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1459_io_a),
    .io_b(FullAdder_1459_io_b),
    .io_ci(FullAdder_1459_io_ci),
    .io_s(FullAdder_1459_io_s),
    .io_co(FullAdder_1459_io_co)
  );
  FullAdder FullAdder_1460 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1460_io_a),
    .io_b(FullAdder_1460_io_b),
    .io_ci(FullAdder_1460_io_ci),
    .io_s(FullAdder_1460_io_s),
    .io_co(FullAdder_1460_io_co)
  );
  FullAdder FullAdder_1461 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1461_io_a),
    .io_b(FullAdder_1461_io_b),
    .io_ci(FullAdder_1461_io_ci),
    .io_s(FullAdder_1461_io_s),
    .io_co(FullAdder_1461_io_co)
  );
  FullAdder FullAdder_1462 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1462_io_a),
    .io_b(FullAdder_1462_io_b),
    .io_ci(FullAdder_1462_io_ci),
    .io_s(FullAdder_1462_io_s),
    .io_co(FullAdder_1462_io_co)
  );
  FullAdder FullAdder_1463 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1463_io_a),
    .io_b(FullAdder_1463_io_b),
    .io_ci(FullAdder_1463_io_ci),
    .io_s(FullAdder_1463_io_s),
    .io_co(FullAdder_1463_io_co)
  );
  FullAdder FullAdder_1464 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1464_io_a),
    .io_b(FullAdder_1464_io_b),
    .io_ci(FullAdder_1464_io_ci),
    .io_s(FullAdder_1464_io_s),
    .io_co(FullAdder_1464_io_co)
  );
  FullAdder FullAdder_1465 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1465_io_a),
    .io_b(FullAdder_1465_io_b),
    .io_ci(FullAdder_1465_io_ci),
    .io_s(FullAdder_1465_io_s),
    .io_co(FullAdder_1465_io_co)
  );
  FullAdder FullAdder_1466 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1466_io_a),
    .io_b(FullAdder_1466_io_b),
    .io_ci(FullAdder_1466_io_ci),
    .io_s(FullAdder_1466_io_s),
    .io_co(FullAdder_1466_io_co)
  );
  FullAdder FullAdder_1467 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1467_io_a),
    .io_b(FullAdder_1467_io_b),
    .io_ci(FullAdder_1467_io_ci),
    .io_s(FullAdder_1467_io_s),
    .io_co(FullAdder_1467_io_co)
  );
  FullAdder FullAdder_1468 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1468_io_a),
    .io_b(FullAdder_1468_io_b),
    .io_ci(FullAdder_1468_io_ci),
    .io_s(FullAdder_1468_io_s),
    .io_co(FullAdder_1468_io_co)
  );
  FullAdder FullAdder_1469 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1469_io_a),
    .io_b(FullAdder_1469_io_b),
    .io_ci(FullAdder_1469_io_ci),
    .io_s(FullAdder_1469_io_s),
    .io_co(FullAdder_1469_io_co)
  );
  FullAdder FullAdder_1470 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1470_io_a),
    .io_b(FullAdder_1470_io_b),
    .io_ci(FullAdder_1470_io_ci),
    .io_s(FullAdder_1470_io_s),
    .io_co(FullAdder_1470_io_co)
  );
  FullAdder FullAdder_1471 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1471_io_a),
    .io_b(FullAdder_1471_io_b),
    .io_ci(FullAdder_1471_io_ci),
    .io_s(FullAdder_1471_io_s),
    .io_co(FullAdder_1471_io_co)
  );
  FullAdder FullAdder_1472 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1472_io_a),
    .io_b(FullAdder_1472_io_b),
    .io_ci(FullAdder_1472_io_ci),
    .io_s(FullAdder_1472_io_s),
    .io_co(FullAdder_1472_io_co)
  );
  FullAdder FullAdder_1473 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1473_io_a),
    .io_b(FullAdder_1473_io_b),
    .io_ci(FullAdder_1473_io_ci),
    .io_s(FullAdder_1473_io_s),
    .io_co(FullAdder_1473_io_co)
  );
  HalfAdder HalfAdder_43 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_43_io_a),
    .io_b(HalfAdder_43_io_b),
    .io_s(HalfAdder_43_io_s),
    .io_co(HalfAdder_43_io_co)
  );
  FullAdder FullAdder_1474 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1474_io_a),
    .io_b(FullAdder_1474_io_b),
    .io_ci(FullAdder_1474_io_ci),
    .io_s(FullAdder_1474_io_s),
    .io_co(FullAdder_1474_io_co)
  );
  FullAdder FullAdder_1475 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1475_io_a),
    .io_b(FullAdder_1475_io_b),
    .io_ci(FullAdder_1475_io_ci),
    .io_s(FullAdder_1475_io_s),
    .io_co(FullAdder_1475_io_co)
  );
  FullAdder FullAdder_1476 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1476_io_a),
    .io_b(FullAdder_1476_io_b),
    .io_ci(FullAdder_1476_io_ci),
    .io_s(FullAdder_1476_io_s),
    .io_co(FullAdder_1476_io_co)
  );
  FullAdder FullAdder_1477 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1477_io_a),
    .io_b(FullAdder_1477_io_b),
    .io_ci(FullAdder_1477_io_ci),
    .io_s(FullAdder_1477_io_s),
    .io_co(FullAdder_1477_io_co)
  );
  FullAdder FullAdder_1478 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1478_io_a),
    .io_b(FullAdder_1478_io_b),
    .io_ci(FullAdder_1478_io_ci),
    .io_s(FullAdder_1478_io_s),
    .io_co(FullAdder_1478_io_co)
  );
  FullAdder FullAdder_1479 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1479_io_a),
    .io_b(FullAdder_1479_io_b),
    .io_ci(FullAdder_1479_io_ci),
    .io_s(FullAdder_1479_io_s),
    .io_co(FullAdder_1479_io_co)
  );
  FullAdder FullAdder_1480 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1480_io_a),
    .io_b(FullAdder_1480_io_b),
    .io_ci(FullAdder_1480_io_ci),
    .io_s(FullAdder_1480_io_s),
    .io_co(FullAdder_1480_io_co)
  );
  FullAdder FullAdder_1481 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1481_io_a),
    .io_b(FullAdder_1481_io_b),
    .io_ci(FullAdder_1481_io_ci),
    .io_s(FullAdder_1481_io_s),
    .io_co(FullAdder_1481_io_co)
  );
  HalfAdder HalfAdder_44 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_44_io_a),
    .io_b(HalfAdder_44_io_b),
    .io_s(HalfAdder_44_io_s),
    .io_co(HalfAdder_44_io_co)
  );
  FullAdder FullAdder_1482 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1482_io_a),
    .io_b(FullAdder_1482_io_b),
    .io_ci(FullAdder_1482_io_ci),
    .io_s(FullAdder_1482_io_s),
    .io_co(FullAdder_1482_io_co)
  );
  FullAdder FullAdder_1483 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1483_io_a),
    .io_b(FullAdder_1483_io_b),
    .io_ci(FullAdder_1483_io_ci),
    .io_s(FullAdder_1483_io_s),
    .io_co(FullAdder_1483_io_co)
  );
  FullAdder FullAdder_1484 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1484_io_a),
    .io_b(FullAdder_1484_io_b),
    .io_ci(FullAdder_1484_io_ci),
    .io_s(FullAdder_1484_io_s),
    .io_co(FullAdder_1484_io_co)
  );
  FullAdder FullAdder_1485 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1485_io_a),
    .io_b(FullAdder_1485_io_b),
    .io_ci(FullAdder_1485_io_ci),
    .io_s(FullAdder_1485_io_s),
    .io_co(FullAdder_1485_io_co)
  );
  FullAdder FullAdder_1486 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1486_io_a),
    .io_b(FullAdder_1486_io_b),
    .io_ci(FullAdder_1486_io_ci),
    .io_s(FullAdder_1486_io_s),
    .io_co(FullAdder_1486_io_co)
  );
  FullAdder FullAdder_1487 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1487_io_a),
    .io_b(FullAdder_1487_io_b),
    .io_ci(FullAdder_1487_io_ci),
    .io_s(FullAdder_1487_io_s),
    .io_co(FullAdder_1487_io_co)
  );
  FullAdder FullAdder_1488 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1488_io_a),
    .io_b(FullAdder_1488_io_b),
    .io_ci(FullAdder_1488_io_ci),
    .io_s(FullAdder_1488_io_s),
    .io_co(FullAdder_1488_io_co)
  );
  FullAdder FullAdder_1489 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1489_io_a),
    .io_b(FullAdder_1489_io_b),
    .io_ci(FullAdder_1489_io_ci),
    .io_s(FullAdder_1489_io_s),
    .io_co(FullAdder_1489_io_co)
  );
  HalfAdder HalfAdder_45 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_45_io_a),
    .io_b(HalfAdder_45_io_b),
    .io_s(HalfAdder_45_io_s),
    .io_co(HalfAdder_45_io_co)
  );
  FullAdder FullAdder_1490 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1490_io_a),
    .io_b(FullAdder_1490_io_b),
    .io_ci(FullAdder_1490_io_ci),
    .io_s(FullAdder_1490_io_s),
    .io_co(FullAdder_1490_io_co)
  );
  FullAdder FullAdder_1491 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1491_io_a),
    .io_b(FullAdder_1491_io_b),
    .io_ci(FullAdder_1491_io_ci),
    .io_s(FullAdder_1491_io_s),
    .io_co(FullAdder_1491_io_co)
  );
  FullAdder FullAdder_1492 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1492_io_a),
    .io_b(FullAdder_1492_io_b),
    .io_ci(FullAdder_1492_io_ci),
    .io_s(FullAdder_1492_io_s),
    .io_co(FullAdder_1492_io_co)
  );
  FullAdder FullAdder_1493 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1493_io_a),
    .io_b(FullAdder_1493_io_b),
    .io_ci(FullAdder_1493_io_ci),
    .io_s(FullAdder_1493_io_s),
    .io_co(FullAdder_1493_io_co)
  );
  FullAdder FullAdder_1494 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1494_io_a),
    .io_b(FullAdder_1494_io_b),
    .io_ci(FullAdder_1494_io_ci),
    .io_s(FullAdder_1494_io_s),
    .io_co(FullAdder_1494_io_co)
  );
  FullAdder FullAdder_1495 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1495_io_a),
    .io_b(FullAdder_1495_io_b),
    .io_ci(FullAdder_1495_io_ci),
    .io_s(FullAdder_1495_io_s),
    .io_co(FullAdder_1495_io_co)
  );
  FullAdder FullAdder_1496 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1496_io_a),
    .io_b(FullAdder_1496_io_b),
    .io_ci(FullAdder_1496_io_ci),
    .io_s(FullAdder_1496_io_s),
    .io_co(FullAdder_1496_io_co)
  );
  FullAdder FullAdder_1497 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1497_io_a),
    .io_b(FullAdder_1497_io_b),
    .io_ci(FullAdder_1497_io_ci),
    .io_s(FullAdder_1497_io_s),
    .io_co(FullAdder_1497_io_co)
  );
  FullAdder FullAdder_1498 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1498_io_a),
    .io_b(FullAdder_1498_io_b),
    .io_ci(FullAdder_1498_io_ci),
    .io_s(FullAdder_1498_io_s),
    .io_co(FullAdder_1498_io_co)
  );
  FullAdder FullAdder_1499 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1499_io_a),
    .io_b(FullAdder_1499_io_b),
    .io_ci(FullAdder_1499_io_ci),
    .io_s(FullAdder_1499_io_s),
    .io_co(FullAdder_1499_io_co)
  );
  FullAdder FullAdder_1500 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1500_io_a),
    .io_b(FullAdder_1500_io_b),
    .io_ci(FullAdder_1500_io_ci),
    .io_s(FullAdder_1500_io_s),
    .io_co(FullAdder_1500_io_co)
  );
  FullAdder FullAdder_1501 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1501_io_a),
    .io_b(FullAdder_1501_io_b),
    .io_ci(FullAdder_1501_io_ci),
    .io_s(FullAdder_1501_io_s),
    .io_co(FullAdder_1501_io_co)
  );
  FullAdder FullAdder_1502 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1502_io_a),
    .io_b(FullAdder_1502_io_b),
    .io_ci(FullAdder_1502_io_ci),
    .io_s(FullAdder_1502_io_s),
    .io_co(FullAdder_1502_io_co)
  );
  FullAdder FullAdder_1503 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1503_io_a),
    .io_b(FullAdder_1503_io_b),
    .io_ci(FullAdder_1503_io_ci),
    .io_s(FullAdder_1503_io_s),
    .io_co(FullAdder_1503_io_co)
  );
  FullAdder FullAdder_1504 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1504_io_a),
    .io_b(FullAdder_1504_io_b),
    .io_ci(FullAdder_1504_io_ci),
    .io_s(FullAdder_1504_io_s),
    .io_co(FullAdder_1504_io_co)
  );
  FullAdder FullAdder_1505 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1505_io_a),
    .io_b(FullAdder_1505_io_b),
    .io_ci(FullAdder_1505_io_ci),
    .io_s(FullAdder_1505_io_s),
    .io_co(FullAdder_1505_io_co)
  );
  FullAdder FullAdder_1506 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1506_io_a),
    .io_b(FullAdder_1506_io_b),
    .io_ci(FullAdder_1506_io_ci),
    .io_s(FullAdder_1506_io_s),
    .io_co(FullAdder_1506_io_co)
  );
  FullAdder FullAdder_1507 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1507_io_a),
    .io_b(FullAdder_1507_io_b),
    .io_ci(FullAdder_1507_io_ci),
    .io_s(FullAdder_1507_io_s),
    .io_co(FullAdder_1507_io_co)
  );
  FullAdder FullAdder_1508 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1508_io_a),
    .io_b(FullAdder_1508_io_b),
    .io_ci(FullAdder_1508_io_ci),
    .io_s(FullAdder_1508_io_s),
    .io_co(FullAdder_1508_io_co)
  );
  FullAdder FullAdder_1509 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1509_io_a),
    .io_b(FullAdder_1509_io_b),
    .io_ci(FullAdder_1509_io_ci),
    .io_s(FullAdder_1509_io_s),
    .io_co(FullAdder_1509_io_co)
  );
  FullAdder FullAdder_1510 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1510_io_a),
    .io_b(FullAdder_1510_io_b),
    .io_ci(FullAdder_1510_io_ci),
    .io_s(FullAdder_1510_io_s),
    .io_co(FullAdder_1510_io_co)
  );
  FullAdder FullAdder_1511 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1511_io_a),
    .io_b(FullAdder_1511_io_b),
    .io_ci(FullAdder_1511_io_ci),
    .io_s(FullAdder_1511_io_s),
    .io_co(FullAdder_1511_io_co)
  );
  FullAdder FullAdder_1512 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1512_io_a),
    .io_b(FullAdder_1512_io_b),
    .io_ci(FullAdder_1512_io_ci),
    .io_s(FullAdder_1512_io_s),
    .io_co(FullAdder_1512_io_co)
  );
  FullAdder FullAdder_1513 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1513_io_a),
    .io_b(FullAdder_1513_io_b),
    .io_ci(FullAdder_1513_io_ci),
    .io_s(FullAdder_1513_io_s),
    .io_co(FullAdder_1513_io_co)
  );
  FullAdder FullAdder_1514 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1514_io_a),
    .io_b(FullAdder_1514_io_b),
    .io_ci(FullAdder_1514_io_ci),
    .io_s(FullAdder_1514_io_s),
    .io_co(FullAdder_1514_io_co)
  );
  FullAdder FullAdder_1515 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1515_io_a),
    .io_b(FullAdder_1515_io_b),
    .io_ci(FullAdder_1515_io_ci),
    .io_s(FullAdder_1515_io_s),
    .io_co(FullAdder_1515_io_co)
  );
  FullAdder FullAdder_1516 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1516_io_a),
    .io_b(FullAdder_1516_io_b),
    .io_ci(FullAdder_1516_io_ci),
    .io_s(FullAdder_1516_io_s),
    .io_co(FullAdder_1516_io_co)
  );
  FullAdder FullAdder_1517 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1517_io_a),
    .io_b(FullAdder_1517_io_b),
    .io_ci(FullAdder_1517_io_ci),
    .io_s(FullAdder_1517_io_s),
    .io_co(FullAdder_1517_io_co)
  );
  FullAdder FullAdder_1518 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1518_io_a),
    .io_b(FullAdder_1518_io_b),
    .io_ci(FullAdder_1518_io_ci),
    .io_s(FullAdder_1518_io_s),
    .io_co(FullAdder_1518_io_co)
  );
  FullAdder FullAdder_1519 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1519_io_a),
    .io_b(FullAdder_1519_io_b),
    .io_ci(FullAdder_1519_io_ci),
    .io_s(FullAdder_1519_io_s),
    .io_co(FullAdder_1519_io_co)
  );
  FullAdder FullAdder_1520 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1520_io_a),
    .io_b(FullAdder_1520_io_b),
    .io_ci(FullAdder_1520_io_ci),
    .io_s(FullAdder_1520_io_s),
    .io_co(FullAdder_1520_io_co)
  );
  FullAdder FullAdder_1521 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1521_io_a),
    .io_b(FullAdder_1521_io_b),
    .io_ci(FullAdder_1521_io_ci),
    .io_s(FullAdder_1521_io_s),
    .io_co(FullAdder_1521_io_co)
  );
  FullAdder FullAdder_1522 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1522_io_a),
    .io_b(FullAdder_1522_io_b),
    .io_ci(FullAdder_1522_io_ci),
    .io_s(FullAdder_1522_io_s),
    .io_co(FullAdder_1522_io_co)
  );
  FullAdder FullAdder_1523 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1523_io_a),
    .io_b(FullAdder_1523_io_b),
    .io_ci(FullAdder_1523_io_ci),
    .io_s(FullAdder_1523_io_s),
    .io_co(FullAdder_1523_io_co)
  );
  FullAdder FullAdder_1524 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1524_io_a),
    .io_b(FullAdder_1524_io_b),
    .io_ci(FullAdder_1524_io_ci),
    .io_s(FullAdder_1524_io_s),
    .io_co(FullAdder_1524_io_co)
  );
  FullAdder FullAdder_1525 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1525_io_a),
    .io_b(FullAdder_1525_io_b),
    .io_ci(FullAdder_1525_io_ci),
    .io_s(FullAdder_1525_io_s),
    .io_co(FullAdder_1525_io_co)
  );
  FullAdder FullAdder_1526 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1526_io_a),
    .io_b(FullAdder_1526_io_b),
    .io_ci(FullAdder_1526_io_ci),
    .io_s(FullAdder_1526_io_s),
    .io_co(FullAdder_1526_io_co)
  );
  FullAdder FullAdder_1527 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1527_io_a),
    .io_b(FullAdder_1527_io_b),
    .io_ci(FullAdder_1527_io_ci),
    .io_s(FullAdder_1527_io_s),
    .io_co(FullAdder_1527_io_co)
  );
  FullAdder FullAdder_1528 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1528_io_a),
    .io_b(FullAdder_1528_io_b),
    .io_ci(FullAdder_1528_io_ci),
    .io_s(FullAdder_1528_io_s),
    .io_co(FullAdder_1528_io_co)
  );
  FullAdder FullAdder_1529 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1529_io_a),
    .io_b(FullAdder_1529_io_b),
    .io_ci(FullAdder_1529_io_ci),
    .io_s(FullAdder_1529_io_s),
    .io_co(FullAdder_1529_io_co)
  );
  FullAdder FullAdder_1530 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1530_io_a),
    .io_b(FullAdder_1530_io_b),
    .io_ci(FullAdder_1530_io_ci),
    .io_s(FullAdder_1530_io_s),
    .io_co(FullAdder_1530_io_co)
  );
  FullAdder FullAdder_1531 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1531_io_a),
    .io_b(FullAdder_1531_io_b),
    .io_ci(FullAdder_1531_io_ci),
    .io_s(FullAdder_1531_io_s),
    .io_co(FullAdder_1531_io_co)
  );
  FullAdder FullAdder_1532 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1532_io_a),
    .io_b(FullAdder_1532_io_b),
    .io_ci(FullAdder_1532_io_ci),
    .io_s(FullAdder_1532_io_s),
    .io_co(FullAdder_1532_io_co)
  );
  FullAdder FullAdder_1533 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1533_io_a),
    .io_b(FullAdder_1533_io_b),
    .io_ci(FullAdder_1533_io_ci),
    .io_s(FullAdder_1533_io_s),
    .io_co(FullAdder_1533_io_co)
  );
  FullAdder FullAdder_1534 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1534_io_a),
    .io_b(FullAdder_1534_io_b),
    .io_ci(FullAdder_1534_io_ci),
    .io_s(FullAdder_1534_io_s),
    .io_co(FullAdder_1534_io_co)
  );
  FullAdder FullAdder_1535 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1535_io_a),
    .io_b(FullAdder_1535_io_b),
    .io_ci(FullAdder_1535_io_ci),
    .io_s(FullAdder_1535_io_s),
    .io_co(FullAdder_1535_io_co)
  );
  FullAdder FullAdder_1536 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1536_io_a),
    .io_b(FullAdder_1536_io_b),
    .io_ci(FullAdder_1536_io_ci),
    .io_s(FullAdder_1536_io_s),
    .io_co(FullAdder_1536_io_co)
  );
  FullAdder FullAdder_1537 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1537_io_a),
    .io_b(FullAdder_1537_io_b),
    .io_ci(FullAdder_1537_io_ci),
    .io_s(FullAdder_1537_io_s),
    .io_co(FullAdder_1537_io_co)
  );
  FullAdder FullAdder_1538 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1538_io_a),
    .io_b(FullAdder_1538_io_b),
    .io_ci(FullAdder_1538_io_ci),
    .io_s(FullAdder_1538_io_s),
    .io_co(FullAdder_1538_io_co)
  );
  FullAdder FullAdder_1539 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1539_io_a),
    .io_b(FullAdder_1539_io_b),
    .io_ci(FullAdder_1539_io_ci),
    .io_s(FullAdder_1539_io_s),
    .io_co(FullAdder_1539_io_co)
  );
  FullAdder FullAdder_1540 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1540_io_a),
    .io_b(FullAdder_1540_io_b),
    .io_ci(FullAdder_1540_io_ci),
    .io_s(FullAdder_1540_io_s),
    .io_co(FullAdder_1540_io_co)
  );
  FullAdder FullAdder_1541 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1541_io_a),
    .io_b(FullAdder_1541_io_b),
    .io_ci(FullAdder_1541_io_ci),
    .io_s(FullAdder_1541_io_s),
    .io_co(FullAdder_1541_io_co)
  );
  FullAdder FullAdder_1542 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1542_io_a),
    .io_b(FullAdder_1542_io_b),
    .io_ci(FullAdder_1542_io_ci),
    .io_s(FullAdder_1542_io_s),
    .io_co(FullAdder_1542_io_co)
  );
  FullAdder FullAdder_1543 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1543_io_a),
    .io_b(FullAdder_1543_io_b),
    .io_ci(FullAdder_1543_io_ci),
    .io_s(FullAdder_1543_io_s),
    .io_co(FullAdder_1543_io_co)
  );
  FullAdder FullAdder_1544 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1544_io_a),
    .io_b(FullAdder_1544_io_b),
    .io_ci(FullAdder_1544_io_ci),
    .io_s(FullAdder_1544_io_s),
    .io_co(FullAdder_1544_io_co)
  );
  FullAdder FullAdder_1545 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1545_io_a),
    .io_b(FullAdder_1545_io_b),
    .io_ci(FullAdder_1545_io_ci),
    .io_s(FullAdder_1545_io_s),
    .io_co(FullAdder_1545_io_co)
  );
  FullAdder FullAdder_1546 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1546_io_a),
    .io_b(FullAdder_1546_io_b),
    .io_ci(FullAdder_1546_io_ci),
    .io_s(FullAdder_1546_io_s),
    .io_co(FullAdder_1546_io_co)
  );
  FullAdder FullAdder_1547 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1547_io_a),
    .io_b(FullAdder_1547_io_b),
    .io_ci(FullAdder_1547_io_ci),
    .io_s(FullAdder_1547_io_s),
    .io_co(FullAdder_1547_io_co)
  );
  FullAdder FullAdder_1548 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1548_io_a),
    .io_b(FullAdder_1548_io_b),
    .io_ci(FullAdder_1548_io_ci),
    .io_s(FullAdder_1548_io_s),
    .io_co(FullAdder_1548_io_co)
  );
  FullAdder FullAdder_1549 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1549_io_a),
    .io_b(FullAdder_1549_io_b),
    .io_ci(FullAdder_1549_io_ci),
    .io_s(FullAdder_1549_io_s),
    .io_co(FullAdder_1549_io_co)
  );
  FullAdder FullAdder_1550 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1550_io_a),
    .io_b(FullAdder_1550_io_b),
    .io_ci(FullAdder_1550_io_ci),
    .io_s(FullAdder_1550_io_s),
    .io_co(FullAdder_1550_io_co)
  );
  FullAdder FullAdder_1551 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1551_io_a),
    .io_b(FullAdder_1551_io_b),
    .io_ci(FullAdder_1551_io_ci),
    .io_s(FullAdder_1551_io_s),
    .io_co(FullAdder_1551_io_co)
  );
  FullAdder FullAdder_1552 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1552_io_a),
    .io_b(FullAdder_1552_io_b),
    .io_ci(FullAdder_1552_io_ci),
    .io_s(FullAdder_1552_io_s),
    .io_co(FullAdder_1552_io_co)
  );
  FullAdder FullAdder_1553 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1553_io_a),
    .io_b(FullAdder_1553_io_b),
    .io_ci(FullAdder_1553_io_ci),
    .io_s(FullAdder_1553_io_s),
    .io_co(FullAdder_1553_io_co)
  );
  FullAdder FullAdder_1554 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1554_io_a),
    .io_b(FullAdder_1554_io_b),
    .io_ci(FullAdder_1554_io_ci),
    .io_s(FullAdder_1554_io_s),
    .io_co(FullAdder_1554_io_co)
  );
  FullAdder FullAdder_1555 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1555_io_a),
    .io_b(FullAdder_1555_io_b),
    .io_ci(FullAdder_1555_io_ci),
    .io_s(FullAdder_1555_io_s),
    .io_co(FullAdder_1555_io_co)
  );
  FullAdder FullAdder_1556 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1556_io_a),
    .io_b(FullAdder_1556_io_b),
    .io_ci(FullAdder_1556_io_ci),
    .io_s(FullAdder_1556_io_s),
    .io_co(FullAdder_1556_io_co)
  );
  FullAdder FullAdder_1557 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1557_io_a),
    .io_b(FullAdder_1557_io_b),
    .io_ci(FullAdder_1557_io_ci),
    .io_s(FullAdder_1557_io_s),
    .io_co(FullAdder_1557_io_co)
  );
  FullAdder FullAdder_1558 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1558_io_a),
    .io_b(FullAdder_1558_io_b),
    .io_ci(FullAdder_1558_io_ci),
    .io_s(FullAdder_1558_io_s),
    .io_co(FullAdder_1558_io_co)
  );
  FullAdder FullAdder_1559 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1559_io_a),
    .io_b(FullAdder_1559_io_b),
    .io_ci(FullAdder_1559_io_ci),
    .io_s(FullAdder_1559_io_s),
    .io_co(FullAdder_1559_io_co)
  );
  FullAdder FullAdder_1560 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1560_io_a),
    .io_b(FullAdder_1560_io_b),
    .io_ci(FullAdder_1560_io_ci),
    .io_s(FullAdder_1560_io_s),
    .io_co(FullAdder_1560_io_co)
  );
  FullAdder FullAdder_1561 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1561_io_a),
    .io_b(FullAdder_1561_io_b),
    .io_ci(FullAdder_1561_io_ci),
    .io_s(FullAdder_1561_io_s),
    .io_co(FullAdder_1561_io_co)
  );
  FullAdder FullAdder_1562 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1562_io_a),
    .io_b(FullAdder_1562_io_b),
    .io_ci(FullAdder_1562_io_ci),
    .io_s(FullAdder_1562_io_s),
    .io_co(FullAdder_1562_io_co)
  );
  FullAdder FullAdder_1563 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1563_io_a),
    .io_b(FullAdder_1563_io_b),
    .io_ci(FullAdder_1563_io_ci),
    .io_s(FullAdder_1563_io_s),
    .io_co(FullAdder_1563_io_co)
  );
  FullAdder FullAdder_1564 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1564_io_a),
    .io_b(FullAdder_1564_io_b),
    .io_ci(FullAdder_1564_io_ci),
    .io_s(FullAdder_1564_io_s),
    .io_co(FullAdder_1564_io_co)
  );
  FullAdder FullAdder_1565 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1565_io_a),
    .io_b(FullAdder_1565_io_b),
    .io_ci(FullAdder_1565_io_ci),
    .io_s(FullAdder_1565_io_s),
    .io_co(FullAdder_1565_io_co)
  );
  FullAdder FullAdder_1566 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1566_io_a),
    .io_b(FullAdder_1566_io_b),
    .io_ci(FullAdder_1566_io_ci),
    .io_s(FullAdder_1566_io_s),
    .io_co(FullAdder_1566_io_co)
  );
  FullAdder FullAdder_1567 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1567_io_a),
    .io_b(FullAdder_1567_io_b),
    .io_ci(FullAdder_1567_io_ci),
    .io_s(FullAdder_1567_io_s),
    .io_co(FullAdder_1567_io_co)
  );
  FullAdder FullAdder_1568 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1568_io_a),
    .io_b(FullAdder_1568_io_b),
    .io_ci(FullAdder_1568_io_ci),
    .io_s(FullAdder_1568_io_s),
    .io_co(FullAdder_1568_io_co)
  );
  FullAdder FullAdder_1569 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1569_io_a),
    .io_b(FullAdder_1569_io_b),
    .io_ci(FullAdder_1569_io_ci),
    .io_s(FullAdder_1569_io_s),
    .io_co(FullAdder_1569_io_co)
  );
  FullAdder FullAdder_1570 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1570_io_a),
    .io_b(FullAdder_1570_io_b),
    .io_ci(FullAdder_1570_io_ci),
    .io_s(FullAdder_1570_io_s),
    .io_co(FullAdder_1570_io_co)
  );
  FullAdder FullAdder_1571 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1571_io_a),
    .io_b(FullAdder_1571_io_b),
    .io_ci(FullAdder_1571_io_ci),
    .io_s(FullAdder_1571_io_s),
    .io_co(FullAdder_1571_io_co)
  );
  FullAdder FullAdder_1572 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1572_io_a),
    .io_b(FullAdder_1572_io_b),
    .io_ci(FullAdder_1572_io_ci),
    .io_s(FullAdder_1572_io_s),
    .io_co(FullAdder_1572_io_co)
  );
  FullAdder FullAdder_1573 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1573_io_a),
    .io_b(FullAdder_1573_io_b),
    .io_ci(FullAdder_1573_io_ci),
    .io_s(FullAdder_1573_io_s),
    .io_co(FullAdder_1573_io_co)
  );
  FullAdder FullAdder_1574 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1574_io_a),
    .io_b(FullAdder_1574_io_b),
    .io_ci(FullAdder_1574_io_ci),
    .io_s(FullAdder_1574_io_s),
    .io_co(FullAdder_1574_io_co)
  );
  FullAdder FullAdder_1575 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1575_io_a),
    .io_b(FullAdder_1575_io_b),
    .io_ci(FullAdder_1575_io_ci),
    .io_s(FullAdder_1575_io_s),
    .io_co(FullAdder_1575_io_co)
  );
  FullAdder FullAdder_1576 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1576_io_a),
    .io_b(FullAdder_1576_io_b),
    .io_ci(FullAdder_1576_io_ci),
    .io_s(FullAdder_1576_io_s),
    .io_co(FullAdder_1576_io_co)
  );
  HalfAdder HalfAdder_46 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_46_io_a),
    .io_b(HalfAdder_46_io_b),
    .io_s(HalfAdder_46_io_s),
    .io_co(HalfAdder_46_io_co)
  );
  FullAdder FullAdder_1577 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1577_io_a),
    .io_b(FullAdder_1577_io_b),
    .io_ci(FullAdder_1577_io_ci),
    .io_s(FullAdder_1577_io_s),
    .io_co(FullAdder_1577_io_co)
  );
  FullAdder FullAdder_1578 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1578_io_a),
    .io_b(FullAdder_1578_io_b),
    .io_ci(FullAdder_1578_io_ci),
    .io_s(FullAdder_1578_io_s),
    .io_co(FullAdder_1578_io_co)
  );
  FullAdder FullAdder_1579 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1579_io_a),
    .io_b(FullAdder_1579_io_b),
    .io_ci(FullAdder_1579_io_ci),
    .io_s(FullAdder_1579_io_s),
    .io_co(FullAdder_1579_io_co)
  );
  FullAdder FullAdder_1580 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1580_io_a),
    .io_b(FullAdder_1580_io_b),
    .io_ci(FullAdder_1580_io_ci),
    .io_s(FullAdder_1580_io_s),
    .io_co(FullAdder_1580_io_co)
  );
  FullAdder FullAdder_1581 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1581_io_a),
    .io_b(FullAdder_1581_io_b),
    .io_ci(FullAdder_1581_io_ci),
    .io_s(FullAdder_1581_io_s),
    .io_co(FullAdder_1581_io_co)
  );
  FullAdder FullAdder_1582 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1582_io_a),
    .io_b(FullAdder_1582_io_b),
    .io_ci(FullAdder_1582_io_ci),
    .io_s(FullAdder_1582_io_s),
    .io_co(FullAdder_1582_io_co)
  );
  FullAdder FullAdder_1583 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1583_io_a),
    .io_b(FullAdder_1583_io_b),
    .io_ci(FullAdder_1583_io_ci),
    .io_s(FullAdder_1583_io_s),
    .io_co(FullAdder_1583_io_co)
  );
  FullAdder FullAdder_1584 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1584_io_a),
    .io_b(FullAdder_1584_io_b),
    .io_ci(FullAdder_1584_io_ci),
    .io_s(FullAdder_1584_io_s),
    .io_co(FullAdder_1584_io_co)
  );
  FullAdder FullAdder_1585 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1585_io_a),
    .io_b(FullAdder_1585_io_b),
    .io_ci(FullAdder_1585_io_ci),
    .io_s(FullAdder_1585_io_s),
    .io_co(FullAdder_1585_io_co)
  );
  FullAdder FullAdder_1586 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1586_io_a),
    .io_b(FullAdder_1586_io_b),
    .io_ci(FullAdder_1586_io_ci),
    .io_s(FullAdder_1586_io_s),
    .io_co(FullAdder_1586_io_co)
  );
  FullAdder FullAdder_1587 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1587_io_a),
    .io_b(FullAdder_1587_io_b),
    .io_ci(FullAdder_1587_io_ci),
    .io_s(FullAdder_1587_io_s),
    .io_co(FullAdder_1587_io_co)
  );
  FullAdder FullAdder_1588 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1588_io_a),
    .io_b(FullAdder_1588_io_b),
    .io_ci(FullAdder_1588_io_ci),
    .io_s(FullAdder_1588_io_s),
    .io_co(FullAdder_1588_io_co)
  );
  FullAdder FullAdder_1589 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1589_io_a),
    .io_b(FullAdder_1589_io_b),
    .io_ci(FullAdder_1589_io_ci),
    .io_s(FullAdder_1589_io_s),
    .io_co(FullAdder_1589_io_co)
  );
  FullAdder FullAdder_1590 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1590_io_a),
    .io_b(FullAdder_1590_io_b),
    .io_ci(FullAdder_1590_io_ci),
    .io_s(FullAdder_1590_io_s),
    .io_co(FullAdder_1590_io_co)
  );
  FullAdder FullAdder_1591 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1591_io_a),
    .io_b(FullAdder_1591_io_b),
    .io_ci(FullAdder_1591_io_ci),
    .io_s(FullAdder_1591_io_s),
    .io_co(FullAdder_1591_io_co)
  );
  FullAdder FullAdder_1592 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1592_io_a),
    .io_b(FullAdder_1592_io_b),
    .io_ci(FullAdder_1592_io_ci),
    .io_s(FullAdder_1592_io_s),
    .io_co(FullAdder_1592_io_co)
  );
  FullAdder FullAdder_1593 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1593_io_a),
    .io_b(FullAdder_1593_io_b),
    .io_ci(FullAdder_1593_io_ci),
    .io_s(FullAdder_1593_io_s),
    .io_co(FullAdder_1593_io_co)
  );
  FullAdder FullAdder_1594 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1594_io_a),
    .io_b(FullAdder_1594_io_b),
    .io_ci(FullAdder_1594_io_ci),
    .io_s(FullAdder_1594_io_s),
    .io_co(FullAdder_1594_io_co)
  );
  FullAdder FullAdder_1595 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1595_io_a),
    .io_b(FullAdder_1595_io_b),
    .io_ci(FullAdder_1595_io_ci),
    .io_s(FullAdder_1595_io_s),
    .io_co(FullAdder_1595_io_co)
  );
  FullAdder FullAdder_1596 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1596_io_a),
    .io_b(FullAdder_1596_io_b),
    .io_ci(FullAdder_1596_io_ci),
    .io_s(FullAdder_1596_io_s),
    .io_co(FullAdder_1596_io_co)
  );
  FullAdder FullAdder_1597 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1597_io_a),
    .io_b(FullAdder_1597_io_b),
    .io_ci(FullAdder_1597_io_ci),
    .io_s(FullAdder_1597_io_s),
    .io_co(FullAdder_1597_io_co)
  );
  FullAdder FullAdder_1598 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1598_io_a),
    .io_b(FullAdder_1598_io_b),
    .io_ci(FullAdder_1598_io_ci),
    .io_s(FullAdder_1598_io_s),
    .io_co(FullAdder_1598_io_co)
  );
  FullAdder FullAdder_1599 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1599_io_a),
    .io_b(FullAdder_1599_io_b),
    .io_ci(FullAdder_1599_io_ci),
    .io_s(FullAdder_1599_io_s),
    .io_co(FullAdder_1599_io_co)
  );
  FullAdder FullAdder_1600 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1600_io_a),
    .io_b(FullAdder_1600_io_b),
    .io_ci(FullAdder_1600_io_ci),
    .io_s(FullAdder_1600_io_s),
    .io_co(FullAdder_1600_io_co)
  );
  FullAdder FullAdder_1601 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1601_io_a),
    .io_b(FullAdder_1601_io_b),
    .io_ci(FullAdder_1601_io_ci),
    .io_s(FullAdder_1601_io_s),
    .io_co(FullAdder_1601_io_co)
  );
  FullAdder FullAdder_1602 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1602_io_a),
    .io_b(FullAdder_1602_io_b),
    .io_ci(FullAdder_1602_io_ci),
    .io_s(FullAdder_1602_io_s),
    .io_co(FullAdder_1602_io_co)
  );
  FullAdder FullAdder_1603 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1603_io_a),
    .io_b(FullAdder_1603_io_b),
    .io_ci(FullAdder_1603_io_ci),
    .io_s(FullAdder_1603_io_s),
    .io_co(FullAdder_1603_io_co)
  );
  FullAdder FullAdder_1604 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1604_io_a),
    .io_b(FullAdder_1604_io_b),
    .io_ci(FullAdder_1604_io_ci),
    .io_s(FullAdder_1604_io_s),
    .io_co(FullAdder_1604_io_co)
  );
  FullAdder FullAdder_1605 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1605_io_a),
    .io_b(FullAdder_1605_io_b),
    .io_ci(FullAdder_1605_io_ci),
    .io_s(FullAdder_1605_io_s),
    .io_co(FullAdder_1605_io_co)
  );
  FullAdder FullAdder_1606 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1606_io_a),
    .io_b(FullAdder_1606_io_b),
    .io_ci(FullAdder_1606_io_ci),
    .io_s(FullAdder_1606_io_s),
    .io_co(FullAdder_1606_io_co)
  );
  FullAdder FullAdder_1607 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1607_io_a),
    .io_b(FullAdder_1607_io_b),
    .io_ci(FullAdder_1607_io_ci),
    .io_s(FullAdder_1607_io_s),
    .io_co(FullAdder_1607_io_co)
  );
  FullAdder FullAdder_1608 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1608_io_a),
    .io_b(FullAdder_1608_io_b),
    .io_ci(FullAdder_1608_io_ci),
    .io_s(FullAdder_1608_io_s),
    .io_co(FullAdder_1608_io_co)
  );
  FullAdder FullAdder_1609 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1609_io_a),
    .io_b(FullAdder_1609_io_b),
    .io_ci(FullAdder_1609_io_ci),
    .io_s(FullAdder_1609_io_s),
    .io_co(FullAdder_1609_io_co)
  );
  FullAdder FullAdder_1610 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1610_io_a),
    .io_b(FullAdder_1610_io_b),
    .io_ci(FullAdder_1610_io_ci),
    .io_s(FullAdder_1610_io_s),
    .io_co(FullAdder_1610_io_co)
  );
  FullAdder FullAdder_1611 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1611_io_a),
    .io_b(FullAdder_1611_io_b),
    .io_ci(FullAdder_1611_io_ci),
    .io_s(FullAdder_1611_io_s),
    .io_co(FullAdder_1611_io_co)
  );
  FullAdder FullAdder_1612 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1612_io_a),
    .io_b(FullAdder_1612_io_b),
    .io_ci(FullAdder_1612_io_ci),
    .io_s(FullAdder_1612_io_s),
    .io_co(FullAdder_1612_io_co)
  );
  FullAdder FullAdder_1613 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1613_io_a),
    .io_b(FullAdder_1613_io_b),
    .io_ci(FullAdder_1613_io_ci),
    .io_s(FullAdder_1613_io_s),
    .io_co(FullAdder_1613_io_co)
  );
  FullAdder FullAdder_1614 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1614_io_a),
    .io_b(FullAdder_1614_io_b),
    .io_ci(FullAdder_1614_io_ci),
    .io_s(FullAdder_1614_io_s),
    .io_co(FullAdder_1614_io_co)
  );
  FullAdder FullAdder_1615 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1615_io_a),
    .io_b(FullAdder_1615_io_b),
    .io_ci(FullAdder_1615_io_ci),
    .io_s(FullAdder_1615_io_s),
    .io_co(FullAdder_1615_io_co)
  );
  FullAdder FullAdder_1616 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1616_io_a),
    .io_b(FullAdder_1616_io_b),
    .io_ci(FullAdder_1616_io_ci),
    .io_s(FullAdder_1616_io_s),
    .io_co(FullAdder_1616_io_co)
  );
  FullAdder FullAdder_1617 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1617_io_a),
    .io_b(FullAdder_1617_io_b),
    .io_ci(FullAdder_1617_io_ci),
    .io_s(FullAdder_1617_io_s),
    .io_co(FullAdder_1617_io_co)
  );
  FullAdder FullAdder_1618 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1618_io_a),
    .io_b(FullAdder_1618_io_b),
    .io_ci(FullAdder_1618_io_ci),
    .io_s(FullAdder_1618_io_s),
    .io_co(FullAdder_1618_io_co)
  );
  FullAdder FullAdder_1619 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1619_io_a),
    .io_b(FullAdder_1619_io_b),
    .io_ci(FullAdder_1619_io_ci),
    .io_s(FullAdder_1619_io_s),
    .io_co(FullAdder_1619_io_co)
  );
  FullAdder FullAdder_1620 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1620_io_a),
    .io_b(FullAdder_1620_io_b),
    .io_ci(FullAdder_1620_io_ci),
    .io_s(FullAdder_1620_io_s),
    .io_co(FullAdder_1620_io_co)
  );
  FullAdder FullAdder_1621 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1621_io_a),
    .io_b(FullAdder_1621_io_b),
    .io_ci(FullAdder_1621_io_ci),
    .io_s(FullAdder_1621_io_s),
    .io_co(FullAdder_1621_io_co)
  );
  FullAdder FullAdder_1622 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1622_io_a),
    .io_b(FullAdder_1622_io_b),
    .io_ci(FullAdder_1622_io_ci),
    .io_s(FullAdder_1622_io_s),
    .io_co(FullAdder_1622_io_co)
  );
  FullAdder FullAdder_1623 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1623_io_a),
    .io_b(FullAdder_1623_io_b),
    .io_ci(FullAdder_1623_io_ci),
    .io_s(FullAdder_1623_io_s),
    .io_co(FullAdder_1623_io_co)
  );
  FullAdder FullAdder_1624 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1624_io_a),
    .io_b(FullAdder_1624_io_b),
    .io_ci(FullAdder_1624_io_ci),
    .io_s(FullAdder_1624_io_s),
    .io_co(FullAdder_1624_io_co)
  );
  FullAdder FullAdder_1625 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1625_io_a),
    .io_b(FullAdder_1625_io_b),
    .io_ci(FullAdder_1625_io_ci),
    .io_s(FullAdder_1625_io_s),
    .io_co(FullAdder_1625_io_co)
  );
  FullAdder FullAdder_1626 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1626_io_a),
    .io_b(FullAdder_1626_io_b),
    .io_ci(FullAdder_1626_io_ci),
    .io_s(FullAdder_1626_io_s),
    .io_co(FullAdder_1626_io_co)
  );
  FullAdder FullAdder_1627 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1627_io_a),
    .io_b(FullAdder_1627_io_b),
    .io_ci(FullAdder_1627_io_ci),
    .io_s(FullAdder_1627_io_s),
    .io_co(FullAdder_1627_io_co)
  );
  FullAdder FullAdder_1628 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1628_io_a),
    .io_b(FullAdder_1628_io_b),
    .io_ci(FullAdder_1628_io_ci),
    .io_s(FullAdder_1628_io_s),
    .io_co(FullAdder_1628_io_co)
  );
  FullAdder FullAdder_1629 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1629_io_a),
    .io_b(FullAdder_1629_io_b),
    .io_ci(FullAdder_1629_io_ci),
    .io_s(FullAdder_1629_io_s),
    .io_co(FullAdder_1629_io_co)
  );
  FullAdder FullAdder_1630 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1630_io_a),
    .io_b(FullAdder_1630_io_b),
    .io_ci(FullAdder_1630_io_ci),
    .io_s(FullAdder_1630_io_s),
    .io_co(FullAdder_1630_io_co)
  );
  FullAdder FullAdder_1631 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1631_io_a),
    .io_b(FullAdder_1631_io_b),
    .io_ci(FullAdder_1631_io_ci),
    .io_s(FullAdder_1631_io_s),
    .io_co(FullAdder_1631_io_co)
  );
  FullAdder FullAdder_1632 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1632_io_a),
    .io_b(FullAdder_1632_io_b),
    .io_ci(FullAdder_1632_io_ci),
    .io_s(FullAdder_1632_io_s),
    .io_co(FullAdder_1632_io_co)
  );
  FullAdder FullAdder_1633 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1633_io_a),
    .io_b(FullAdder_1633_io_b),
    .io_ci(FullAdder_1633_io_ci),
    .io_s(FullAdder_1633_io_s),
    .io_co(FullAdder_1633_io_co)
  );
  FullAdder FullAdder_1634 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1634_io_a),
    .io_b(FullAdder_1634_io_b),
    .io_ci(FullAdder_1634_io_ci),
    .io_s(FullAdder_1634_io_s),
    .io_co(FullAdder_1634_io_co)
  );
  FullAdder FullAdder_1635 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1635_io_a),
    .io_b(FullAdder_1635_io_b),
    .io_ci(FullAdder_1635_io_ci),
    .io_s(FullAdder_1635_io_s),
    .io_co(FullAdder_1635_io_co)
  );
  FullAdder FullAdder_1636 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1636_io_a),
    .io_b(FullAdder_1636_io_b),
    .io_ci(FullAdder_1636_io_ci),
    .io_s(FullAdder_1636_io_s),
    .io_co(FullAdder_1636_io_co)
  );
  FullAdder FullAdder_1637 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1637_io_a),
    .io_b(FullAdder_1637_io_b),
    .io_ci(FullAdder_1637_io_ci),
    .io_s(FullAdder_1637_io_s),
    .io_co(FullAdder_1637_io_co)
  );
  FullAdder FullAdder_1638 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1638_io_a),
    .io_b(FullAdder_1638_io_b),
    .io_ci(FullAdder_1638_io_ci),
    .io_s(FullAdder_1638_io_s),
    .io_co(FullAdder_1638_io_co)
  );
  FullAdder FullAdder_1639 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1639_io_a),
    .io_b(FullAdder_1639_io_b),
    .io_ci(FullAdder_1639_io_ci),
    .io_s(FullAdder_1639_io_s),
    .io_co(FullAdder_1639_io_co)
  );
  FullAdder FullAdder_1640 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1640_io_a),
    .io_b(FullAdder_1640_io_b),
    .io_ci(FullAdder_1640_io_ci),
    .io_s(FullAdder_1640_io_s),
    .io_co(FullAdder_1640_io_co)
  );
  FullAdder FullAdder_1641 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1641_io_a),
    .io_b(FullAdder_1641_io_b),
    .io_ci(FullAdder_1641_io_ci),
    .io_s(FullAdder_1641_io_s),
    .io_co(FullAdder_1641_io_co)
  );
  FullAdder FullAdder_1642 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1642_io_a),
    .io_b(FullAdder_1642_io_b),
    .io_ci(FullAdder_1642_io_ci),
    .io_s(FullAdder_1642_io_s),
    .io_co(FullAdder_1642_io_co)
  );
  FullAdder FullAdder_1643 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1643_io_a),
    .io_b(FullAdder_1643_io_b),
    .io_ci(FullAdder_1643_io_ci),
    .io_s(FullAdder_1643_io_s),
    .io_co(FullAdder_1643_io_co)
  );
  FullAdder FullAdder_1644 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1644_io_a),
    .io_b(FullAdder_1644_io_b),
    .io_ci(FullAdder_1644_io_ci),
    .io_s(FullAdder_1644_io_s),
    .io_co(FullAdder_1644_io_co)
  );
  FullAdder FullAdder_1645 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1645_io_a),
    .io_b(FullAdder_1645_io_b),
    .io_ci(FullAdder_1645_io_ci),
    .io_s(FullAdder_1645_io_s),
    .io_co(FullAdder_1645_io_co)
  );
  FullAdder FullAdder_1646 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1646_io_a),
    .io_b(FullAdder_1646_io_b),
    .io_ci(FullAdder_1646_io_ci),
    .io_s(FullAdder_1646_io_s),
    .io_co(FullAdder_1646_io_co)
  );
  FullAdder FullAdder_1647 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1647_io_a),
    .io_b(FullAdder_1647_io_b),
    .io_ci(FullAdder_1647_io_ci),
    .io_s(FullAdder_1647_io_s),
    .io_co(FullAdder_1647_io_co)
  );
  FullAdder FullAdder_1648 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1648_io_a),
    .io_b(FullAdder_1648_io_b),
    .io_ci(FullAdder_1648_io_ci),
    .io_s(FullAdder_1648_io_s),
    .io_co(FullAdder_1648_io_co)
  );
  FullAdder FullAdder_1649 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1649_io_a),
    .io_b(FullAdder_1649_io_b),
    .io_ci(FullAdder_1649_io_ci),
    .io_s(FullAdder_1649_io_s),
    .io_co(FullAdder_1649_io_co)
  );
  FullAdder FullAdder_1650 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1650_io_a),
    .io_b(FullAdder_1650_io_b),
    .io_ci(FullAdder_1650_io_ci),
    .io_s(FullAdder_1650_io_s),
    .io_co(FullAdder_1650_io_co)
  );
  FullAdder FullAdder_1651 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1651_io_a),
    .io_b(FullAdder_1651_io_b),
    .io_ci(FullAdder_1651_io_ci),
    .io_s(FullAdder_1651_io_s),
    .io_co(FullAdder_1651_io_co)
  );
  FullAdder FullAdder_1652 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1652_io_a),
    .io_b(FullAdder_1652_io_b),
    .io_ci(FullAdder_1652_io_ci),
    .io_s(FullAdder_1652_io_s),
    .io_co(FullAdder_1652_io_co)
  );
  FullAdder FullAdder_1653 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1653_io_a),
    .io_b(FullAdder_1653_io_b),
    .io_ci(FullAdder_1653_io_ci),
    .io_s(FullAdder_1653_io_s),
    .io_co(FullAdder_1653_io_co)
  );
  FullAdder FullAdder_1654 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1654_io_a),
    .io_b(FullAdder_1654_io_b),
    .io_ci(FullAdder_1654_io_ci),
    .io_s(FullAdder_1654_io_s),
    .io_co(FullAdder_1654_io_co)
  );
  FullAdder FullAdder_1655 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1655_io_a),
    .io_b(FullAdder_1655_io_b),
    .io_ci(FullAdder_1655_io_ci),
    .io_s(FullAdder_1655_io_s),
    .io_co(FullAdder_1655_io_co)
  );
  FullAdder FullAdder_1656 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1656_io_a),
    .io_b(FullAdder_1656_io_b),
    .io_ci(FullAdder_1656_io_ci),
    .io_s(FullAdder_1656_io_s),
    .io_co(FullAdder_1656_io_co)
  );
  FullAdder FullAdder_1657 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1657_io_a),
    .io_b(FullAdder_1657_io_b),
    .io_ci(FullAdder_1657_io_ci),
    .io_s(FullAdder_1657_io_s),
    .io_co(FullAdder_1657_io_co)
  );
  HalfAdder HalfAdder_47 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_47_io_a),
    .io_b(HalfAdder_47_io_b),
    .io_s(HalfAdder_47_io_s),
    .io_co(HalfAdder_47_io_co)
  );
  FullAdder FullAdder_1658 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1658_io_a),
    .io_b(FullAdder_1658_io_b),
    .io_ci(FullAdder_1658_io_ci),
    .io_s(FullAdder_1658_io_s),
    .io_co(FullAdder_1658_io_co)
  );
  FullAdder FullAdder_1659 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1659_io_a),
    .io_b(FullAdder_1659_io_b),
    .io_ci(FullAdder_1659_io_ci),
    .io_s(FullAdder_1659_io_s),
    .io_co(FullAdder_1659_io_co)
  );
  FullAdder FullAdder_1660 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1660_io_a),
    .io_b(FullAdder_1660_io_b),
    .io_ci(FullAdder_1660_io_ci),
    .io_s(FullAdder_1660_io_s),
    .io_co(FullAdder_1660_io_co)
  );
  FullAdder FullAdder_1661 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1661_io_a),
    .io_b(FullAdder_1661_io_b),
    .io_ci(FullAdder_1661_io_ci),
    .io_s(FullAdder_1661_io_s),
    .io_co(FullAdder_1661_io_co)
  );
  FullAdder FullAdder_1662 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1662_io_a),
    .io_b(FullAdder_1662_io_b),
    .io_ci(FullAdder_1662_io_ci),
    .io_s(FullAdder_1662_io_s),
    .io_co(FullAdder_1662_io_co)
  );
  FullAdder FullAdder_1663 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1663_io_a),
    .io_b(FullAdder_1663_io_b),
    .io_ci(FullAdder_1663_io_ci),
    .io_s(FullAdder_1663_io_s),
    .io_co(FullAdder_1663_io_co)
  );
  FullAdder FullAdder_1664 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1664_io_a),
    .io_b(FullAdder_1664_io_b),
    .io_ci(FullAdder_1664_io_ci),
    .io_s(FullAdder_1664_io_s),
    .io_co(FullAdder_1664_io_co)
  );
  FullAdder FullAdder_1665 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1665_io_a),
    .io_b(FullAdder_1665_io_b),
    .io_ci(FullAdder_1665_io_ci),
    .io_s(FullAdder_1665_io_s),
    .io_co(FullAdder_1665_io_co)
  );
  FullAdder FullAdder_1666 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1666_io_a),
    .io_b(FullAdder_1666_io_b),
    .io_ci(FullAdder_1666_io_ci),
    .io_s(FullAdder_1666_io_s),
    .io_co(FullAdder_1666_io_co)
  );
  FullAdder FullAdder_1667 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1667_io_a),
    .io_b(FullAdder_1667_io_b),
    .io_ci(FullAdder_1667_io_ci),
    .io_s(FullAdder_1667_io_s),
    .io_co(FullAdder_1667_io_co)
  );
  FullAdder FullAdder_1668 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1668_io_a),
    .io_b(FullAdder_1668_io_b),
    .io_ci(FullAdder_1668_io_ci),
    .io_s(FullAdder_1668_io_s),
    .io_co(FullAdder_1668_io_co)
  );
  FullAdder FullAdder_1669 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1669_io_a),
    .io_b(FullAdder_1669_io_b),
    .io_ci(FullAdder_1669_io_ci),
    .io_s(FullAdder_1669_io_s),
    .io_co(FullAdder_1669_io_co)
  );
  HalfAdder HalfAdder_48 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_48_io_a),
    .io_b(HalfAdder_48_io_b),
    .io_s(HalfAdder_48_io_s),
    .io_co(HalfAdder_48_io_co)
  );
  FullAdder FullAdder_1670 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1670_io_a),
    .io_b(FullAdder_1670_io_b),
    .io_ci(FullAdder_1670_io_ci),
    .io_s(FullAdder_1670_io_s),
    .io_co(FullAdder_1670_io_co)
  );
  FullAdder FullAdder_1671 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1671_io_a),
    .io_b(FullAdder_1671_io_b),
    .io_ci(FullAdder_1671_io_ci),
    .io_s(FullAdder_1671_io_s),
    .io_co(FullAdder_1671_io_co)
  );
  FullAdder FullAdder_1672 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1672_io_a),
    .io_b(FullAdder_1672_io_b),
    .io_ci(FullAdder_1672_io_ci),
    .io_s(FullAdder_1672_io_s),
    .io_co(FullAdder_1672_io_co)
  );
  FullAdder FullAdder_1673 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1673_io_a),
    .io_b(FullAdder_1673_io_b),
    .io_ci(FullAdder_1673_io_ci),
    .io_s(FullAdder_1673_io_s),
    .io_co(FullAdder_1673_io_co)
  );
  FullAdder FullAdder_1674 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1674_io_a),
    .io_b(FullAdder_1674_io_b),
    .io_ci(FullAdder_1674_io_ci),
    .io_s(FullAdder_1674_io_s),
    .io_co(FullAdder_1674_io_co)
  );
  FullAdder FullAdder_1675 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1675_io_a),
    .io_b(FullAdder_1675_io_b),
    .io_ci(FullAdder_1675_io_ci),
    .io_s(FullAdder_1675_io_s),
    .io_co(FullAdder_1675_io_co)
  );
  FullAdder FullAdder_1676 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1676_io_a),
    .io_b(FullAdder_1676_io_b),
    .io_ci(FullAdder_1676_io_ci),
    .io_s(FullAdder_1676_io_s),
    .io_co(FullAdder_1676_io_co)
  );
  FullAdder FullAdder_1677 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1677_io_a),
    .io_b(FullAdder_1677_io_b),
    .io_ci(FullAdder_1677_io_ci),
    .io_s(FullAdder_1677_io_s),
    .io_co(FullAdder_1677_io_co)
  );
  FullAdder FullAdder_1678 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1678_io_a),
    .io_b(FullAdder_1678_io_b),
    .io_ci(FullAdder_1678_io_ci),
    .io_s(FullAdder_1678_io_s),
    .io_co(FullAdder_1678_io_co)
  );
  FullAdder FullAdder_1679 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1679_io_a),
    .io_b(FullAdder_1679_io_b),
    .io_ci(FullAdder_1679_io_ci),
    .io_s(FullAdder_1679_io_s),
    .io_co(FullAdder_1679_io_co)
  );
  FullAdder FullAdder_1680 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1680_io_a),
    .io_b(FullAdder_1680_io_b),
    .io_ci(FullAdder_1680_io_ci),
    .io_s(FullAdder_1680_io_s),
    .io_co(FullAdder_1680_io_co)
  );
  FullAdder FullAdder_1681 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1681_io_a),
    .io_b(FullAdder_1681_io_b),
    .io_ci(FullAdder_1681_io_ci),
    .io_s(FullAdder_1681_io_s),
    .io_co(FullAdder_1681_io_co)
  );
  FullAdder FullAdder_1682 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1682_io_a),
    .io_b(FullAdder_1682_io_b),
    .io_ci(FullAdder_1682_io_ci),
    .io_s(FullAdder_1682_io_s),
    .io_co(FullAdder_1682_io_co)
  );
  FullAdder FullAdder_1683 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1683_io_a),
    .io_b(FullAdder_1683_io_b),
    .io_ci(FullAdder_1683_io_ci),
    .io_s(FullAdder_1683_io_s),
    .io_co(FullAdder_1683_io_co)
  );
  FullAdder FullAdder_1684 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1684_io_a),
    .io_b(FullAdder_1684_io_b),
    .io_ci(FullAdder_1684_io_ci),
    .io_s(FullAdder_1684_io_s),
    .io_co(FullAdder_1684_io_co)
  );
  FullAdder FullAdder_1685 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1685_io_a),
    .io_b(FullAdder_1685_io_b),
    .io_ci(FullAdder_1685_io_ci),
    .io_s(FullAdder_1685_io_s),
    .io_co(FullAdder_1685_io_co)
  );
  FullAdder FullAdder_1686 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1686_io_a),
    .io_b(FullAdder_1686_io_b),
    .io_ci(FullAdder_1686_io_ci),
    .io_s(FullAdder_1686_io_s),
    .io_co(FullAdder_1686_io_co)
  );
  FullAdder FullAdder_1687 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1687_io_a),
    .io_b(FullAdder_1687_io_b),
    .io_ci(FullAdder_1687_io_ci),
    .io_s(FullAdder_1687_io_s),
    .io_co(FullAdder_1687_io_co)
  );
  FullAdder FullAdder_1688 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1688_io_a),
    .io_b(FullAdder_1688_io_b),
    .io_ci(FullAdder_1688_io_ci),
    .io_s(FullAdder_1688_io_s),
    .io_co(FullAdder_1688_io_co)
  );
  FullAdder FullAdder_1689 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1689_io_a),
    .io_b(FullAdder_1689_io_b),
    .io_ci(FullAdder_1689_io_ci),
    .io_s(FullAdder_1689_io_s),
    .io_co(FullAdder_1689_io_co)
  );
  FullAdder FullAdder_1690 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1690_io_a),
    .io_b(FullAdder_1690_io_b),
    .io_ci(FullAdder_1690_io_ci),
    .io_s(FullAdder_1690_io_s),
    .io_co(FullAdder_1690_io_co)
  );
  FullAdder FullAdder_1691 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1691_io_a),
    .io_b(FullAdder_1691_io_b),
    .io_ci(FullAdder_1691_io_ci),
    .io_s(FullAdder_1691_io_s),
    .io_co(FullAdder_1691_io_co)
  );
  FullAdder FullAdder_1692 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1692_io_a),
    .io_b(FullAdder_1692_io_b),
    .io_ci(FullAdder_1692_io_ci),
    .io_s(FullAdder_1692_io_s),
    .io_co(FullAdder_1692_io_co)
  );
  FullAdder FullAdder_1693 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1693_io_a),
    .io_b(FullAdder_1693_io_b),
    .io_ci(FullAdder_1693_io_ci),
    .io_s(FullAdder_1693_io_s),
    .io_co(FullAdder_1693_io_co)
  );
  FullAdder FullAdder_1694 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1694_io_a),
    .io_b(FullAdder_1694_io_b),
    .io_ci(FullAdder_1694_io_ci),
    .io_s(FullAdder_1694_io_s),
    .io_co(FullAdder_1694_io_co)
  );
  FullAdder FullAdder_1695 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1695_io_a),
    .io_b(FullAdder_1695_io_b),
    .io_ci(FullAdder_1695_io_ci),
    .io_s(FullAdder_1695_io_s),
    .io_co(FullAdder_1695_io_co)
  );
  FullAdder FullAdder_1696 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1696_io_a),
    .io_b(FullAdder_1696_io_b),
    .io_ci(FullAdder_1696_io_ci),
    .io_s(FullAdder_1696_io_s),
    .io_co(FullAdder_1696_io_co)
  );
  FullAdder FullAdder_1697 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1697_io_a),
    .io_b(FullAdder_1697_io_b),
    .io_ci(FullAdder_1697_io_ci),
    .io_s(FullAdder_1697_io_s),
    .io_co(FullAdder_1697_io_co)
  );
  FullAdder FullAdder_1698 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1698_io_a),
    .io_b(FullAdder_1698_io_b),
    .io_ci(FullAdder_1698_io_ci),
    .io_s(FullAdder_1698_io_s),
    .io_co(FullAdder_1698_io_co)
  );
  FullAdder FullAdder_1699 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1699_io_a),
    .io_b(FullAdder_1699_io_b),
    .io_ci(FullAdder_1699_io_ci),
    .io_s(FullAdder_1699_io_s),
    .io_co(FullAdder_1699_io_co)
  );
  FullAdder FullAdder_1700 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1700_io_a),
    .io_b(FullAdder_1700_io_b),
    .io_ci(FullAdder_1700_io_ci),
    .io_s(FullAdder_1700_io_s),
    .io_co(FullAdder_1700_io_co)
  );
  FullAdder FullAdder_1701 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1701_io_a),
    .io_b(FullAdder_1701_io_b),
    .io_ci(FullAdder_1701_io_ci),
    .io_s(FullAdder_1701_io_s),
    .io_co(FullAdder_1701_io_co)
  );
  FullAdder FullAdder_1702 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1702_io_a),
    .io_b(FullAdder_1702_io_b),
    .io_ci(FullAdder_1702_io_ci),
    .io_s(FullAdder_1702_io_s),
    .io_co(FullAdder_1702_io_co)
  );
  FullAdder FullAdder_1703 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1703_io_a),
    .io_b(FullAdder_1703_io_b),
    .io_ci(FullAdder_1703_io_ci),
    .io_s(FullAdder_1703_io_s),
    .io_co(FullAdder_1703_io_co)
  );
  FullAdder FullAdder_1704 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1704_io_a),
    .io_b(FullAdder_1704_io_b),
    .io_ci(FullAdder_1704_io_ci),
    .io_s(FullAdder_1704_io_s),
    .io_co(FullAdder_1704_io_co)
  );
  FullAdder FullAdder_1705 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1705_io_a),
    .io_b(FullAdder_1705_io_b),
    .io_ci(FullAdder_1705_io_ci),
    .io_s(FullAdder_1705_io_s),
    .io_co(FullAdder_1705_io_co)
  );
  FullAdder FullAdder_1706 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1706_io_a),
    .io_b(FullAdder_1706_io_b),
    .io_ci(FullAdder_1706_io_ci),
    .io_s(FullAdder_1706_io_s),
    .io_co(FullAdder_1706_io_co)
  );
  FullAdder FullAdder_1707 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1707_io_a),
    .io_b(FullAdder_1707_io_b),
    .io_ci(FullAdder_1707_io_ci),
    .io_s(FullAdder_1707_io_s),
    .io_co(FullAdder_1707_io_co)
  );
  FullAdder FullAdder_1708 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1708_io_a),
    .io_b(FullAdder_1708_io_b),
    .io_ci(FullAdder_1708_io_ci),
    .io_s(FullAdder_1708_io_s),
    .io_co(FullAdder_1708_io_co)
  );
  FullAdder FullAdder_1709 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1709_io_a),
    .io_b(FullAdder_1709_io_b),
    .io_ci(FullAdder_1709_io_ci),
    .io_s(FullAdder_1709_io_s),
    .io_co(FullAdder_1709_io_co)
  );
  FullAdder FullAdder_1710 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1710_io_a),
    .io_b(FullAdder_1710_io_b),
    .io_ci(FullAdder_1710_io_ci),
    .io_s(FullAdder_1710_io_s),
    .io_co(FullAdder_1710_io_co)
  );
  FullAdder FullAdder_1711 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1711_io_a),
    .io_b(FullAdder_1711_io_b),
    .io_ci(FullAdder_1711_io_ci),
    .io_s(FullAdder_1711_io_s),
    .io_co(FullAdder_1711_io_co)
  );
  FullAdder FullAdder_1712 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1712_io_a),
    .io_b(FullAdder_1712_io_b),
    .io_ci(FullAdder_1712_io_ci),
    .io_s(FullAdder_1712_io_s),
    .io_co(FullAdder_1712_io_co)
  );
  FullAdder FullAdder_1713 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1713_io_a),
    .io_b(FullAdder_1713_io_b),
    .io_ci(FullAdder_1713_io_ci),
    .io_s(FullAdder_1713_io_s),
    .io_co(FullAdder_1713_io_co)
  );
  FullAdder FullAdder_1714 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1714_io_a),
    .io_b(FullAdder_1714_io_b),
    .io_ci(FullAdder_1714_io_ci),
    .io_s(FullAdder_1714_io_s),
    .io_co(FullAdder_1714_io_co)
  );
  FullAdder FullAdder_1715 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1715_io_a),
    .io_b(FullAdder_1715_io_b),
    .io_ci(FullAdder_1715_io_ci),
    .io_s(FullAdder_1715_io_s),
    .io_co(FullAdder_1715_io_co)
  );
  FullAdder FullAdder_1716 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1716_io_a),
    .io_b(FullAdder_1716_io_b),
    .io_ci(FullAdder_1716_io_ci),
    .io_s(FullAdder_1716_io_s),
    .io_co(FullAdder_1716_io_co)
  );
  FullAdder FullAdder_1717 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1717_io_a),
    .io_b(FullAdder_1717_io_b),
    .io_ci(FullAdder_1717_io_ci),
    .io_s(FullAdder_1717_io_s),
    .io_co(FullAdder_1717_io_co)
  );
  FullAdder FullAdder_1718 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1718_io_a),
    .io_b(FullAdder_1718_io_b),
    .io_ci(FullAdder_1718_io_ci),
    .io_s(FullAdder_1718_io_s),
    .io_co(FullAdder_1718_io_co)
  );
  FullAdder FullAdder_1719 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1719_io_a),
    .io_b(FullAdder_1719_io_b),
    .io_ci(FullAdder_1719_io_ci),
    .io_s(FullAdder_1719_io_s),
    .io_co(FullAdder_1719_io_co)
  );
  FullAdder FullAdder_1720 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1720_io_a),
    .io_b(FullAdder_1720_io_b),
    .io_ci(FullAdder_1720_io_ci),
    .io_s(FullAdder_1720_io_s),
    .io_co(FullAdder_1720_io_co)
  );
  FullAdder FullAdder_1721 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1721_io_a),
    .io_b(FullAdder_1721_io_b),
    .io_ci(FullAdder_1721_io_ci),
    .io_s(FullAdder_1721_io_s),
    .io_co(FullAdder_1721_io_co)
  );
  FullAdder FullAdder_1722 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1722_io_a),
    .io_b(FullAdder_1722_io_b),
    .io_ci(FullAdder_1722_io_ci),
    .io_s(FullAdder_1722_io_s),
    .io_co(FullAdder_1722_io_co)
  );
  FullAdder FullAdder_1723 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1723_io_a),
    .io_b(FullAdder_1723_io_b),
    .io_ci(FullAdder_1723_io_ci),
    .io_s(FullAdder_1723_io_s),
    .io_co(FullAdder_1723_io_co)
  );
  FullAdder FullAdder_1724 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1724_io_a),
    .io_b(FullAdder_1724_io_b),
    .io_ci(FullAdder_1724_io_ci),
    .io_s(FullAdder_1724_io_s),
    .io_co(FullAdder_1724_io_co)
  );
  FullAdder FullAdder_1725 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1725_io_a),
    .io_b(FullAdder_1725_io_b),
    .io_ci(FullAdder_1725_io_ci),
    .io_s(FullAdder_1725_io_s),
    .io_co(FullAdder_1725_io_co)
  );
  FullAdder FullAdder_1726 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1726_io_a),
    .io_b(FullAdder_1726_io_b),
    .io_ci(FullAdder_1726_io_ci),
    .io_s(FullAdder_1726_io_s),
    .io_co(FullAdder_1726_io_co)
  );
  FullAdder FullAdder_1727 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1727_io_a),
    .io_b(FullAdder_1727_io_b),
    .io_ci(FullAdder_1727_io_ci),
    .io_s(FullAdder_1727_io_s),
    .io_co(FullAdder_1727_io_co)
  );
  FullAdder FullAdder_1728 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1728_io_a),
    .io_b(FullAdder_1728_io_b),
    .io_ci(FullAdder_1728_io_ci),
    .io_s(FullAdder_1728_io_s),
    .io_co(FullAdder_1728_io_co)
  );
  FullAdder FullAdder_1729 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1729_io_a),
    .io_b(FullAdder_1729_io_b),
    .io_ci(FullAdder_1729_io_ci),
    .io_s(FullAdder_1729_io_s),
    .io_co(FullAdder_1729_io_co)
  );
  FullAdder FullAdder_1730 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1730_io_a),
    .io_b(FullAdder_1730_io_b),
    .io_ci(FullAdder_1730_io_ci),
    .io_s(FullAdder_1730_io_s),
    .io_co(FullAdder_1730_io_co)
  );
  FullAdder FullAdder_1731 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1731_io_a),
    .io_b(FullAdder_1731_io_b),
    .io_ci(FullAdder_1731_io_ci),
    .io_s(FullAdder_1731_io_s),
    .io_co(FullAdder_1731_io_co)
  );
  FullAdder FullAdder_1732 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1732_io_a),
    .io_b(FullAdder_1732_io_b),
    .io_ci(FullAdder_1732_io_ci),
    .io_s(FullAdder_1732_io_s),
    .io_co(FullAdder_1732_io_co)
  );
  FullAdder FullAdder_1733 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1733_io_a),
    .io_b(FullAdder_1733_io_b),
    .io_ci(FullAdder_1733_io_ci),
    .io_s(FullAdder_1733_io_s),
    .io_co(FullAdder_1733_io_co)
  );
  FullAdder FullAdder_1734 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1734_io_a),
    .io_b(FullAdder_1734_io_b),
    .io_ci(FullAdder_1734_io_ci),
    .io_s(FullAdder_1734_io_s),
    .io_co(FullAdder_1734_io_co)
  );
  FullAdder FullAdder_1735 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1735_io_a),
    .io_b(FullAdder_1735_io_b),
    .io_ci(FullAdder_1735_io_ci),
    .io_s(FullAdder_1735_io_s),
    .io_co(FullAdder_1735_io_co)
  );
  FullAdder FullAdder_1736 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1736_io_a),
    .io_b(FullAdder_1736_io_b),
    .io_ci(FullAdder_1736_io_ci),
    .io_s(FullAdder_1736_io_s),
    .io_co(FullAdder_1736_io_co)
  );
  FullAdder FullAdder_1737 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1737_io_a),
    .io_b(FullAdder_1737_io_b),
    .io_ci(FullAdder_1737_io_ci),
    .io_s(FullAdder_1737_io_s),
    .io_co(FullAdder_1737_io_co)
  );
  FullAdder FullAdder_1738 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1738_io_a),
    .io_b(FullAdder_1738_io_b),
    .io_ci(FullAdder_1738_io_ci),
    .io_s(FullAdder_1738_io_s),
    .io_co(FullAdder_1738_io_co)
  );
  FullAdder FullAdder_1739 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1739_io_a),
    .io_b(FullAdder_1739_io_b),
    .io_ci(FullAdder_1739_io_ci),
    .io_s(FullAdder_1739_io_s),
    .io_co(FullAdder_1739_io_co)
  );
  FullAdder FullAdder_1740 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1740_io_a),
    .io_b(FullAdder_1740_io_b),
    .io_ci(FullAdder_1740_io_ci),
    .io_s(FullAdder_1740_io_s),
    .io_co(FullAdder_1740_io_co)
  );
  FullAdder FullAdder_1741 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1741_io_a),
    .io_b(FullAdder_1741_io_b),
    .io_ci(FullAdder_1741_io_ci),
    .io_s(FullAdder_1741_io_s),
    .io_co(FullAdder_1741_io_co)
  );
  FullAdder FullAdder_1742 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1742_io_a),
    .io_b(FullAdder_1742_io_b),
    .io_ci(FullAdder_1742_io_ci),
    .io_s(FullAdder_1742_io_s),
    .io_co(FullAdder_1742_io_co)
  );
  FullAdder FullAdder_1743 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1743_io_a),
    .io_b(FullAdder_1743_io_b),
    .io_ci(FullAdder_1743_io_ci),
    .io_s(FullAdder_1743_io_s),
    .io_co(FullAdder_1743_io_co)
  );
  FullAdder FullAdder_1744 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1744_io_a),
    .io_b(FullAdder_1744_io_b),
    .io_ci(FullAdder_1744_io_ci),
    .io_s(FullAdder_1744_io_s),
    .io_co(FullAdder_1744_io_co)
  );
  FullAdder FullAdder_1745 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1745_io_a),
    .io_b(FullAdder_1745_io_b),
    .io_ci(FullAdder_1745_io_ci),
    .io_s(FullAdder_1745_io_s),
    .io_co(FullAdder_1745_io_co)
  );
  FullAdder FullAdder_1746 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1746_io_a),
    .io_b(FullAdder_1746_io_b),
    .io_ci(FullAdder_1746_io_ci),
    .io_s(FullAdder_1746_io_s),
    .io_co(FullAdder_1746_io_co)
  );
  FullAdder FullAdder_1747 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1747_io_a),
    .io_b(FullAdder_1747_io_b),
    .io_ci(FullAdder_1747_io_ci),
    .io_s(FullAdder_1747_io_s),
    .io_co(FullAdder_1747_io_co)
  );
  FullAdder FullAdder_1748 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1748_io_a),
    .io_b(FullAdder_1748_io_b),
    .io_ci(FullAdder_1748_io_ci),
    .io_s(FullAdder_1748_io_s),
    .io_co(FullAdder_1748_io_co)
  );
  FullAdder FullAdder_1749 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1749_io_a),
    .io_b(FullAdder_1749_io_b),
    .io_ci(FullAdder_1749_io_ci),
    .io_s(FullAdder_1749_io_s),
    .io_co(FullAdder_1749_io_co)
  );
  FullAdder FullAdder_1750 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1750_io_a),
    .io_b(FullAdder_1750_io_b),
    .io_ci(FullAdder_1750_io_ci),
    .io_s(FullAdder_1750_io_s),
    .io_co(FullAdder_1750_io_co)
  );
  FullAdder FullAdder_1751 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1751_io_a),
    .io_b(FullAdder_1751_io_b),
    .io_ci(FullAdder_1751_io_ci),
    .io_s(FullAdder_1751_io_s),
    .io_co(FullAdder_1751_io_co)
  );
  FullAdder FullAdder_1752 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1752_io_a),
    .io_b(FullAdder_1752_io_b),
    .io_ci(FullAdder_1752_io_ci),
    .io_s(FullAdder_1752_io_s),
    .io_co(FullAdder_1752_io_co)
  );
  FullAdder FullAdder_1753 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1753_io_a),
    .io_b(FullAdder_1753_io_b),
    .io_ci(FullAdder_1753_io_ci),
    .io_s(FullAdder_1753_io_s),
    .io_co(FullAdder_1753_io_co)
  );
  FullAdder FullAdder_1754 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1754_io_a),
    .io_b(FullAdder_1754_io_b),
    .io_ci(FullAdder_1754_io_ci),
    .io_s(FullAdder_1754_io_s),
    .io_co(FullAdder_1754_io_co)
  );
  FullAdder FullAdder_1755 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1755_io_a),
    .io_b(FullAdder_1755_io_b),
    .io_ci(FullAdder_1755_io_ci),
    .io_s(FullAdder_1755_io_s),
    .io_co(FullAdder_1755_io_co)
  );
  FullAdder FullAdder_1756 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1756_io_a),
    .io_b(FullAdder_1756_io_b),
    .io_ci(FullAdder_1756_io_ci),
    .io_s(FullAdder_1756_io_s),
    .io_co(FullAdder_1756_io_co)
  );
  FullAdder FullAdder_1757 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1757_io_a),
    .io_b(FullAdder_1757_io_b),
    .io_ci(FullAdder_1757_io_ci),
    .io_s(FullAdder_1757_io_s),
    .io_co(FullAdder_1757_io_co)
  );
  FullAdder FullAdder_1758 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1758_io_a),
    .io_b(FullAdder_1758_io_b),
    .io_ci(FullAdder_1758_io_ci),
    .io_s(FullAdder_1758_io_s),
    .io_co(FullAdder_1758_io_co)
  );
  FullAdder FullAdder_1759 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1759_io_a),
    .io_b(FullAdder_1759_io_b),
    .io_ci(FullAdder_1759_io_ci),
    .io_s(FullAdder_1759_io_s),
    .io_co(FullAdder_1759_io_co)
  );
  FullAdder FullAdder_1760 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1760_io_a),
    .io_b(FullAdder_1760_io_b),
    .io_ci(FullAdder_1760_io_ci),
    .io_s(FullAdder_1760_io_s),
    .io_co(FullAdder_1760_io_co)
  );
  FullAdder FullAdder_1761 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1761_io_a),
    .io_b(FullAdder_1761_io_b),
    .io_ci(FullAdder_1761_io_ci),
    .io_s(FullAdder_1761_io_s),
    .io_co(FullAdder_1761_io_co)
  );
  FullAdder FullAdder_1762 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1762_io_a),
    .io_b(FullAdder_1762_io_b),
    .io_ci(FullAdder_1762_io_ci),
    .io_s(FullAdder_1762_io_s),
    .io_co(FullAdder_1762_io_co)
  );
  FullAdder FullAdder_1763 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1763_io_a),
    .io_b(FullAdder_1763_io_b),
    .io_ci(FullAdder_1763_io_ci),
    .io_s(FullAdder_1763_io_s),
    .io_co(FullAdder_1763_io_co)
  );
  FullAdder FullAdder_1764 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1764_io_a),
    .io_b(FullAdder_1764_io_b),
    .io_ci(FullAdder_1764_io_ci),
    .io_s(FullAdder_1764_io_s),
    .io_co(FullAdder_1764_io_co)
  );
  FullAdder FullAdder_1765 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1765_io_a),
    .io_b(FullAdder_1765_io_b),
    .io_ci(FullAdder_1765_io_ci),
    .io_s(FullAdder_1765_io_s),
    .io_co(FullAdder_1765_io_co)
  );
  FullAdder FullAdder_1766 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1766_io_a),
    .io_b(FullAdder_1766_io_b),
    .io_ci(FullAdder_1766_io_ci),
    .io_s(FullAdder_1766_io_s),
    .io_co(FullAdder_1766_io_co)
  );
  FullAdder FullAdder_1767 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1767_io_a),
    .io_b(FullAdder_1767_io_b),
    .io_ci(FullAdder_1767_io_ci),
    .io_s(FullAdder_1767_io_s),
    .io_co(FullAdder_1767_io_co)
  );
  FullAdder FullAdder_1768 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1768_io_a),
    .io_b(FullAdder_1768_io_b),
    .io_ci(FullAdder_1768_io_ci),
    .io_s(FullAdder_1768_io_s),
    .io_co(FullAdder_1768_io_co)
  );
  FullAdder FullAdder_1769 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1769_io_a),
    .io_b(FullAdder_1769_io_b),
    .io_ci(FullAdder_1769_io_ci),
    .io_s(FullAdder_1769_io_s),
    .io_co(FullAdder_1769_io_co)
  );
  FullAdder FullAdder_1770 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1770_io_a),
    .io_b(FullAdder_1770_io_b),
    .io_ci(FullAdder_1770_io_ci),
    .io_s(FullAdder_1770_io_s),
    .io_co(FullAdder_1770_io_co)
  );
  FullAdder FullAdder_1771 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1771_io_a),
    .io_b(FullAdder_1771_io_b),
    .io_ci(FullAdder_1771_io_ci),
    .io_s(FullAdder_1771_io_s),
    .io_co(FullAdder_1771_io_co)
  );
  FullAdder FullAdder_1772 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1772_io_a),
    .io_b(FullAdder_1772_io_b),
    .io_ci(FullAdder_1772_io_ci),
    .io_s(FullAdder_1772_io_s),
    .io_co(FullAdder_1772_io_co)
  );
  FullAdder FullAdder_1773 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1773_io_a),
    .io_b(FullAdder_1773_io_b),
    .io_ci(FullAdder_1773_io_ci),
    .io_s(FullAdder_1773_io_s),
    .io_co(FullAdder_1773_io_co)
  );
  FullAdder FullAdder_1774 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1774_io_a),
    .io_b(FullAdder_1774_io_b),
    .io_ci(FullAdder_1774_io_ci),
    .io_s(FullAdder_1774_io_s),
    .io_co(FullAdder_1774_io_co)
  );
  FullAdder FullAdder_1775 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1775_io_a),
    .io_b(FullAdder_1775_io_b),
    .io_ci(FullAdder_1775_io_ci),
    .io_s(FullAdder_1775_io_s),
    .io_co(FullAdder_1775_io_co)
  );
  FullAdder FullAdder_1776 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1776_io_a),
    .io_b(FullAdder_1776_io_b),
    .io_ci(FullAdder_1776_io_ci),
    .io_s(FullAdder_1776_io_s),
    .io_co(FullAdder_1776_io_co)
  );
  FullAdder FullAdder_1777 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1777_io_a),
    .io_b(FullAdder_1777_io_b),
    .io_ci(FullAdder_1777_io_ci),
    .io_s(FullAdder_1777_io_s),
    .io_co(FullAdder_1777_io_co)
  );
  FullAdder FullAdder_1778 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1778_io_a),
    .io_b(FullAdder_1778_io_b),
    .io_ci(FullAdder_1778_io_ci),
    .io_s(FullAdder_1778_io_s),
    .io_co(FullAdder_1778_io_co)
  );
  FullAdder FullAdder_1779 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1779_io_a),
    .io_b(FullAdder_1779_io_b),
    .io_ci(FullAdder_1779_io_ci),
    .io_s(FullAdder_1779_io_s),
    .io_co(FullAdder_1779_io_co)
  );
  FullAdder FullAdder_1780 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1780_io_a),
    .io_b(FullAdder_1780_io_b),
    .io_ci(FullAdder_1780_io_ci),
    .io_s(FullAdder_1780_io_s),
    .io_co(FullAdder_1780_io_co)
  );
  FullAdder FullAdder_1781 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1781_io_a),
    .io_b(FullAdder_1781_io_b),
    .io_ci(FullAdder_1781_io_ci),
    .io_s(FullAdder_1781_io_s),
    .io_co(FullAdder_1781_io_co)
  );
  FullAdder FullAdder_1782 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1782_io_a),
    .io_b(FullAdder_1782_io_b),
    .io_ci(FullAdder_1782_io_ci),
    .io_s(FullAdder_1782_io_s),
    .io_co(FullAdder_1782_io_co)
  );
  FullAdder FullAdder_1783 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1783_io_a),
    .io_b(FullAdder_1783_io_b),
    .io_ci(FullAdder_1783_io_ci),
    .io_s(FullAdder_1783_io_s),
    .io_co(FullAdder_1783_io_co)
  );
  FullAdder FullAdder_1784 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1784_io_a),
    .io_b(FullAdder_1784_io_b),
    .io_ci(FullAdder_1784_io_ci),
    .io_s(FullAdder_1784_io_s),
    .io_co(FullAdder_1784_io_co)
  );
  FullAdder FullAdder_1785 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1785_io_a),
    .io_b(FullAdder_1785_io_b),
    .io_ci(FullAdder_1785_io_ci),
    .io_s(FullAdder_1785_io_s),
    .io_co(FullAdder_1785_io_co)
  );
  FullAdder FullAdder_1786 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1786_io_a),
    .io_b(FullAdder_1786_io_b),
    .io_ci(FullAdder_1786_io_ci),
    .io_s(FullAdder_1786_io_s),
    .io_co(FullAdder_1786_io_co)
  );
  FullAdder FullAdder_1787 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1787_io_a),
    .io_b(FullAdder_1787_io_b),
    .io_ci(FullAdder_1787_io_ci),
    .io_s(FullAdder_1787_io_s),
    .io_co(FullAdder_1787_io_co)
  );
  FullAdder FullAdder_1788 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1788_io_a),
    .io_b(FullAdder_1788_io_b),
    .io_ci(FullAdder_1788_io_ci),
    .io_s(FullAdder_1788_io_s),
    .io_co(FullAdder_1788_io_co)
  );
  FullAdder FullAdder_1789 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1789_io_a),
    .io_b(FullAdder_1789_io_b),
    .io_ci(FullAdder_1789_io_ci),
    .io_s(FullAdder_1789_io_s),
    .io_co(FullAdder_1789_io_co)
  );
  FullAdder FullAdder_1790 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1790_io_a),
    .io_b(FullAdder_1790_io_b),
    .io_ci(FullAdder_1790_io_ci),
    .io_s(FullAdder_1790_io_s),
    .io_co(FullAdder_1790_io_co)
  );
  FullAdder FullAdder_1791 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1791_io_a),
    .io_b(FullAdder_1791_io_b),
    .io_ci(FullAdder_1791_io_ci),
    .io_s(FullAdder_1791_io_s),
    .io_co(FullAdder_1791_io_co)
  );
  FullAdder FullAdder_1792 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1792_io_a),
    .io_b(FullAdder_1792_io_b),
    .io_ci(FullAdder_1792_io_ci),
    .io_s(FullAdder_1792_io_s),
    .io_co(FullAdder_1792_io_co)
  );
  FullAdder FullAdder_1793 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1793_io_a),
    .io_b(FullAdder_1793_io_b),
    .io_ci(FullAdder_1793_io_ci),
    .io_s(FullAdder_1793_io_s),
    .io_co(FullAdder_1793_io_co)
  );
  FullAdder FullAdder_1794 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1794_io_a),
    .io_b(FullAdder_1794_io_b),
    .io_ci(FullAdder_1794_io_ci),
    .io_s(FullAdder_1794_io_s),
    .io_co(FullAdder_1794_io_co)
  );
  FullAdder FullAdder_1795 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1795_io_a),
    .io_b(FullAdder_1795_io_b),
    .io_ci(FullAdder_1795_io_ci),
    .io_s(FullAdder_1795_io_s),
    .io_co(FullAdder_1795_io_co)
  );
  FullAdder FullAdder_1796 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1796_io_a),
    .io_b(FullAdder_1796_io_b),
    .io_ci(FullAdder_1796_io_ci),
    .io_s(FullAdder_1796_io_s),
    .io_co(FullAdder_1796_io_co)
  );
  FullAdder FullAdder_1797 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1797_io_a),
    .io_b(FullAdder_1797_io_b),
    .io_ci(FullAdder_1797_io_ci),
    .io_s(FullAdder_1797_io_s),
    .io_co(FullAdder_1797_io_co)
  );
  FullAdder FullAdder_1798 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1798_io_a),
    .io_b(FullAdder_1798_io_b),
    .io_ci(FullAdder_1798_io_ci),
    .io_s(FullAdder_1798_io_s),
    .io_co(FullAdder_1798_io_co)
  );
  FullAdder FullAdder_1799 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1799_io_a),
    .io_b(FullAdder_1799_io_b),
    .io_ci(FullAdder_1799_io_ci),
    .io_s(FullAdder_1799_io_s),
    .io_co(FullAdder_1799_io_co)
  );
  FullAdder FullAdder_1800 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1800_io_a),
    .io_b(FullAdder_1800_io_b),
    .io_ci(FullAdder_1800_io_ci),
    .io_s(FullAdder_1800_io_s),
    .io_co(FullAdder_1800_io_co)
  );
  FullAdder FullAdder_1801 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1801_io_a),
    .io_b(FullAdder_1801_io_b),
    .io_ci(FullAdder_1801_io_ci),
    .io_s(FullAdder_1801_io_s),
    .io_co(FullAdder_1801_io_co)
  );
  FullAdder FullAdder_1802 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1802_io_a),
    .io_b(FullAdder_1802_io_b),
    .io_ci(FullAdder_1802_io_ci),
    .io_s(FullAdder_1802_io_s),
    .io_co(FullAdder_1802_io_co)
  );
  FullAdder FullAdder_1803 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1803_io_a),
    .io_b(FullAdder_1803_io_b),
    .io_ci(FullAdder_1803_io_ci),
    .io_s(FullAdder_1803_io_s),
    .io_co(FullAdder_1803_io_co)
  );
  HalfAdder HalfAdder_49 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_49_io_a),
    .io_b(HalfAdder_49_io_b),
    .io_s(HalfAdder_49_io_s),
    .io_co(HalfAdder_49_io_co)
  );
  FullAdder FullAdder_1804 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1804_io_a),
    .io_b(FullAdder_1804_io_b),
    .io_ci(FullAdder_1804_io_ci),
    .io_s(FullAdder_1804_io_s),
    .io_co(FullAdder_1804_io_co)
  );
  FullAdder FullAdder_1805 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1805_io_a),
    .io_b(FullAdder_1805_io_b),
    .io_ci(FullAdder_1805_io_ci),
    .io_s(FullAdder_1805_io_s),
    .io_co(FullAdder_1805_io_co)
  );
  FullAdder FullAdder_1806 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1806_io_a),
    .io_b(FullAdder_1806_io_b),
    .io_ci(FullAdder_1806_io_ci),
    .io_s(FullAdder_1806_io_s),
    .io_co(FullAdder_1806_io_co)
  );
  FullAdder FullAdder_1807 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1807_io_a),
    .io_b(FullAdder_1807_io_b),
    .io_ci(FullAdder_1807_io_ci),
    .io_s(FullAdder_1807_io_s),
    .io_co(FullAdder_1807_io_co)
  );
  FullAdder FullAdder_1808 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1808_io_a),
    .io_b(FullAdder_1808_io_b),
    .io_ci(FullAdder_1808_io_ci),
    .io_s(FullAdder_1808_io_s),
    .io_co(FullAdder_1808_io_co)
  );
  FullAdder FullAdder_1809 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1809_io_a),
    .io_b(FullAdder_1809_io_b),
    .io_ci(FullAdder_1809_io_ci),
    .io_s(FullAdder_1809_io_s),
    .io_co(FullAdder_1809_io_co)
  );
  FullAdder FullAdder_1810 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1810_io_a),
    .io_b(FullAdder_1810_io_b),
    .io_ci(FullAdder_1810_io_ci),
    .io_s(FullAdder_1810_io_s),
    .io_co(FullAdder_1810_io_co)
  );
  FullAdder FullAdder_1811 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1811_io_a),
    .io_b(FullAdder_1811_io_b),
    .io_ci(FullAdder_1811_io_ci),
    .io_s(FullAdder_1811_io_s),
    .io_co(FullAdder_1811_io_co)
  );
  FullAdder FullAdder_1812 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1812_io_a),
    .io_b(FullAdder_1812_io_b),
    .io_ci(FullAdder_1812_io_ci),
    .io_s(FullAdder_1812_io_s),
    .io_co(FullAdder_1812_io_co)
  );
  FullAdder FullAdder_1813 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1813_io_a),
    .io_b(FullAdder_1813_io_b),
    .io_ci(FullAdder_1813_io_ci),
    .io_s(FullAdder_1813_io_s),
    .io_co(FullAdder_1813_io_co)
  );
  FullAdder FullAdder_1814 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1814_io_a),
    .io_b(FullAdder_1814_io_b),
    .io_ci(FullAdder_1814_io_ci),
    .io_s(FullAdder_1814_io_s),
    .io_co(FullAdder_1814_io_co)
  );
  FullAdder FullAdder_1815 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1815_io_a),
    .io_b(FullAdder_1815_io_b),
    .io_ci(FullAdder_1815_io_ci),
    .io_s(FullAdder_1815_io_s),
    .io_co(FullAdder_1815_io_co)
  );
  FullAdder FullAdder_1816 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1816_io_a),
    .io_b(FullAdder_1816_io_b),
    .io_ci(FullAdder_1816_io_ci),
    .io_s(FullAdder_1816_io_s),
    .io_co(FullAdder_1816_io_co)
  );
  FullAdder FullAdder_1817 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1817_io_a),
    .io_b(FullAdder_1817_io_b),
    .io_ci(FullAdder_1817_io_ci),
    .io_s(FullAdder_1817_io_s),
    .io_co(FullAdder_1817_io_co)
  );
  FullAdder FullAdder_1818 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1818_io_a),
    .io_b(FullAdder_1818_io_b),
    .io_ci(FullAdder_1818_io_ci),
    .io_s(FullAdder_1818_io_s),
    .io_co(FullAdder_1818_io_co)
  );
  FullAdder FullAdder_1819 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1819_io_a),
    .io_b(FullAdder_1819_io_b),
    .io_ci(FullAdder_1819_io_ci),
    .io_s(FullAdder_1819_io_s),
    .io_co(FullAdder_1819_io_co)
  );
  FullAdder FullAdder_1820 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1820_io_a),
    .io_b(FullAdder_1820_io_b),
    .io_ci(FullAdder_1820_io_ci),
    .io_s(FullAdder_1820_io_s),
    .io_co(FullAdder_1820_io_co)
  );
  FullAdder FullAdder_1821 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1821_io_a),
    .io_b(FullAdder_1821_io_b),
    .io_ci(FullAdder_1821_io_ci),
    .io_s(FullAdder_1821_io_s),
    .io_co(FullAdder_1821_io_co)
  );
  FullAdder FullAdder_1822 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1822_io_a),
    .io_b(FullAdder_1822_io_b),
    .io_ci(FullAdder_1822_io_ci),
    .io_s(FullAdder_1822_io_s),
    .io_co(FullAdder_1822_io_co)
  );
  FullAdder FullAdder_1823 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1823_io_a),
    .io_b(FullAdder_1823_io_b),
    .io_ci(FullAdder_1823_io_ci),
    .io_s(FullAdder_1823_io_s),
    .io_co(FullAdder_1823_io_co)
  );
  FullAdder FullAdder_1824 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1824_io_a),
    .io_b(FullAdder_1824_io_b),
    .io_ci(FullAdder_1824_io_ci),
    .io_s(FullAdder_1824_io_s),
    .io_co(FullAdder_1824_io_co)
  );
  FullAdder FullAdder_1825 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1825_io_a),
    .io_b(FullAdder_1825_io_b),
    .io_ci(FullAdder_1825_io_ci),
    .io_s(FullAdder_1825_io_s),
    .io_co(FullAdder_1825_io_co)
  );
  FullAdder FullAdder_1826 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1826_io_a),
    .io_b(FullAdder_1826_io_b),
    .io_ci(FullAdder_1826_io_ci),
    .io_s(FullAdder_1826_io_s),
    .io_co(FullAdder_1826_io_co)
  );
  FullAdder FullAdder_1827 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1827_io_a),
    .io_b(FullAdder_1827_io_b),
    .io_ci(FullAdder_1827_io_ci),
    .io_s(FullAdder_1827_io_s),
    .io_co(FullAdder_1827_io_co)
  );
  FullAdder FullAdder_1828 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1828_io_a),
    .io_b(FullAdder_1828_io_b),
    .io_ci(FullAdder_1828_io_ci),
    .io_s(FullAdder_1828_io_s),
    .io_co(FullAdder_1828_io_co)
  );
  FullAdder FullAdder_1829 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1829_io_a),
    .io_b(FullAdder_1829_io_b),
    .io_ci(FullAdder_1829_io_ci),
    .io_s(FullAdder_1829_io_s),
    .io_co(FullAdder_1829_io_co)
  );
  FullAdder FullAdder_1830 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1830_io_a),
    .io_b(FullAdder_1830_io_b),
    .io_ci(FullAdder_1830_io_ci),
    .io_s(FullAdder_1830_io_s),
    .io_co(FullAdder_1830_io_co)
  );
  FullAdder FullAdder_1831 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1831_io_a),
    .io_b(FullAdder_1831_io_b),
    .io_ci(FullAdder_1831_io_ci),
    .io_s(FullAdder_1831_io_s),
    .io_co(FullAdder_1831_io_co)
  );
  FullAdder FullAdder_1832 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1832_io_a),
    .io_b(FullAdder_1832_io_b),
    .io_ci(FullAdder_1832_io_ci),
    .io_s(FullAdder_1832_io_s),
    .io_co(FullAdder_1832_io_co)
  );
  FullAdder FullAdder_1833 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1833_io_a),
    .io_b(FullAdder_1833_io_b),
    .io_ci(FullAdder_1833_io_ci),
    .io_s(FullAdder_1833_io_s),
    .io_co(FullAdder_1833_io_co)
  );
  FullAdder FullAdder_1834 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1834_io_a),
    .io_b(FullAdder_1834_io_b),
    .io_ci(FullAdder_1834_io_ci),
    .io_s(FullAdder_1834_io_s),
    .io_co(FullAdder_1834_io_co)
  );
  FullAdder FullAdder_1835 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1835_io_a),
    .io_b(FullAdder_1835_io_b),
    .io_ci(FullAdder_1835_io_ci),
    .io_s(FullAdder_1835_io_s),
    .io_co(FullAdder_1835_io_co)
  );
  FullAdder FullAdder_1836 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1836_io_a),
    .io_b(FullAdder_1836_io_b),
    .io_ci(FullAdder_1836_io_ci),
    .io_s(FullAdder_1836_io_s),
    .io_co(FullAdder_1836_io_co)
  );
  FullAdder FullAdder_1837 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1837_io_a),
    .io_b(FullAdder_1837_io_b),
    .io_ci(FullAdder_1837_io_ci),
    .io_s(FullAdder_1837_io_s),
    .io_co(FullAdder_1837_io_co)
  );
  FullAdder FullAdder_1838 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1838_io_a),
    .io_b(FullAdder_1838_io_b),
    .io_ci(FullAdder_1838_io_ci),
    .io_s(FullAdder_1838_io_s),
    .io_co(FullAdder_1838_io_co)
  );
  FullAdder FullAdder_1839 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1839_io_a),
    .io_b(FullAdder_1839_io_b),
    .io_ci(FullAdder_1839_io_ci),
    .io_s(FullAdder_1839_io_s),
    .io_co(FullAdder_1839_io_co)
  );
  FullAdder FullAdder_1840 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1840_io_a),
    .io_b(FullAdder_1840_io_b),
    .io_ci(FullAdder_1840_io_ci),
    .io_s(FullAdder_1840_io_s),
    .io_co(FullAdder_1840_io_co)
  );
  FullAdder FullAdder_1841 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1841_io_a),
    .io_b(FullAdder_1841_io_b),
    .io_ci(FullAdder_1841_io_ci),
    .io_s(FullAdder_1841_io_s),
    .io_co(FullAdder_1841_io_co)
  );
  FullAdder FullAdder_1842 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1842_io_a),
    .io_b(FullAdder_1842_io_b),
    .io_ci(FullAdder_1842_io_ci),
    .io_s(FullAdder_1842_io_s),
    .io_co(FullAdder_1842_io_co)
  );
  FullAdder FullAdder_1843 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1843_io_a),
    .io_b(FullAdder_1843_io_b),
    .io_ci(FullAdder_1843_io_ci),
    .io_s(FullAdder_1843_io_s),
    .io_co(FullAdder_1843_io_co)
  );
  FullAdder FullAdder_1844 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1844_io_a),
    .io_b(FullAdder_1844_io_b),
    .io_ci(FullAdder_1844_io_ci),
    .io_s(FullAdder_1844_io_s),
    .io_co(FullAdder_1844_io_co)
  );
  FullAdder FullAdder_1845 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1845_io_a),
    .io_b(FullAdder_1845_io_b),
    .io_ci(FullAdder_1845_io_ci),
    .io_s(FullAdder_1845_io_s),
    .io_co(FullAdder_1845_io_co)
  );
  FullAdder FullAdder_1846 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1846_io_a),
    .io_b(FullAdder_1846_io_b),
    .io_ci(FullAdder_1846_io_ci),
    .io_s(FullAdder_1846_io_s),
    .io_co(FullAdder_1846_io_co)
  );
  FullAdder FullAdder_1847 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1847_io_a),
    .io_b(FullAdder_1847_io_b),
    .io_ci(FullAdder_1847_io_ci),
    .io_s(FullAdder_1847_io_s),
    .io_co(FullAdder_1847_io_co)
  );
  FullAdder FullAdder_1848 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1848_io_a),
    .io_b(FullAdder_1848_io_b),
    .io_ci(FullAdder_1848_io_ci),
    .io_s(FullAdder_1848_io_s),
    .io_co(FullAdder_1848_io_co)
  );
  FullAdder FullAdder_1849 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1849_io_a),
    .io_b(FullAdder_1849_io_b),
    .io_ci(FullAdder_1849_io_ci),
    .io_s(FullAdder_1849_io_s),
    .io_co(FullAdder_1849_io_co)
  );
  FullAdder FullAdder_1850 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1850_io_a),
    .io_b(FullAdder_1850_io_b),
    .io_ci(FullAdder_1850_io_ci),
    .io_s(FullAdder_1850_io_s),
    .io_co(FullAdder_1850_io_co)
  );
  FullAdder FullAdder_1851 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1851_io_a),
    .io_b(FullAdder_1851_io_b),
    .io_ci(FullAdder_1851_io_ci),
    .io_s(FullAdder_1851_io_s),
    .io_co(FullAdder_1851_io_co)
  );
  FullAdder FullAdder_1852 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1852_io_a),
    .io_b(FullAdder_1852_io_b),
    .io_ci(FullAdder_1852_io_ci),
    .io_s(FullAdder_1852_io_s),
    .io_co(FullAdder_1852_io_co)
  );
  FullAdder FullAdder_1853 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1853_io_a),
    .io_b(FullAdder_1853_io_b),
    .io_ci(FullAdder_1853_io_ci),
    .io_s(FullAdder_1853_io_s),
    .io_co(FullAdder_1853_io_co)
  );
  FullAdder FullAdder_1854 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1854_io_a),
    .io_b(FullAdder_1854_io_b),
    .io_ci(FullAdder_1854_io_ci),
    .io_s(FullAdder_1854_io_s),
    .io_co(FullAdder_1854_io_co)
  );
  FullAdder FullAdder_1855 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1855_io_a),
    .io_b(FullAdder_1855_io_b),
    .io_ci(FullAdder_1855_io_ci),
    .io_s(FullAdder_1855_io_s),
    .io_co(FullAdder_1855_io_co)
  );
  FullAdder FullAdder_1856 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1856_io_a),
    .io_b(FullAdder_1856_io_b),
    .io_ci(FullAdder_1856_io_ci),
    .io_s(FullAdder_1856_io_s),
    .io_co(FullAdder_1856_io_co)
  );
  FullAdder FullAdder_1857 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1857_io_a),
    .io_b(FullAdder_1857_io_b),
    .io_ci(FullAdder_1857_io_ci),
    .io_s(FullAdder_1857_io_s),
    .io_co(FullAdder_1857_io_co)
  );
  FullAdder FullAdder_1858 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1858_io_a),
    .io_b(FullAdder_1858_io_b),
    .io_ci(FullAdder_1858_io_ci),
    .io_s(FullAdder_1858_io_s),
    .io_co(FullAdder_1858_io_co)
  );
  FullAdder FullAdder_1859 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1859_io_a),
    .io_b(FullAdder_1859_io_b),
    .io_ci(FullAdder_1859_io_ci),
    .io_s(FullAdder_1859_io_s),
    .io_co(FullAdder_1859_io_co)
  );
  FullAdder FullAdder_1860 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1860_io_a),
    .io_b(FullAdder_1860_io_b),
    .io_ci(FullAdder_1860_io_ci),
    .io_s(FullAdder_1860_io_s),
    .io_co(FullAdder_1860_io_co)
  );
  FullAdder FullAdder_1861 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1861_io_a),
    .io_b(FullAdder_1861_io_b),
    .io_ci(FullAdder_1861_io_ci),
    .io_s(FullAdder_1861_io_s),
    .io_co(FullAdder_1861_io_co)
  );
  FullAdder FullAdder_1862 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1862_io_a),
    .io_b(FullAdder_1862_io_b),
    .io_ci(FullAdder_1862_io_ci),
    .io_s(FullAdder_1862_io_s),
    .io_co(FullAdder_1862_io_co)
  );
  FullAdder FullAdder_1863 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1863_io_a),
    .io_b(FullAdder_1863_io_b),
    .io_ci(FullAdder_1863_io_ci),
    .io_s(FullAdder_1863_io_s),
    .io_co(FullAdder_1863_io_co)
  );
  FullAdder FullAdder_1864 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1864_io_a),
    .io_b(FullAdder_1864_io_b),
    .io_ci(FullAdder_1864_io_ci),
    .io_s(FullAdder_1864_io_s),
    .io_co(FullAdder_1864_io_co)
  );
  FullAdder FullAdder_1865 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1865_io_a),
    .io_b(FullAdder_1865_io_b),
    .io_ci(FullAdder_1865_io_ci),
    .io_s(FullAdder_1865_io_s),
    .io_co(FullAdder_1865_io_co)
  );
  FullAdder FullAdder_1866 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1866_io_a),
    .io_b(FullAdder_1866_io_b),
    .io_ci(FullAdder_1866_io_ci),
    .io_s(FullAdder_1866_io_s),
    .io_co(FullAdder_1866_io_co)
  );
  FullAdder FullAdder_1867 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1867_io_a),
    .io_b(FullAdder_1867_io_b),
    .io_ci(FullAdder_1867_io_ci),
    .io_s(FullAdder_1867_io_s),
    .io_co(FullAdder_1867_io_co)
  );
  FullAdder FullAdder_1868 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1868_io_a),
    .io_b(FullAdder_1868_io_b),
    .io_ci(FullAdder_1868_io_ci),
    .io_s(FullAdder_1868_io_s),
    .io_co(FullAdder_1868_io_co)
  );
  FullAdder FullAdder_1869 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1869_io_a),
    .io_b(FullAdder_1869_io_b),
    .io_ci(FullAdder_1869_io_ci),
    .io_s(FullAdder_1869_io_s),
    .io_co(FullAdder_1869_io_co)
  );
  FullAdder FullAdder_1870 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1870_io_a),
    .io_b(FullAdder_1870_io_b),
    .io_ci(FullAdder_1870_io_ci),
    .io_s(FullAdder_1870_io_s),
    .io_co(FullAdder_1870_io_co)
  );
  FullAdder FullAdder_1871 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1871_io_a),
    .io_b(FullAdder_1871_io_b),
    .io_ci(FullAdder_1871_io_ci),
    .io_s(FullAdder_1871_io_s),
    .io_co(FullAdder_1871_io_co)
  );
  FullAdder FullAdder_1872 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1872_io_a),
    .io_b(FullAdder_1872_io_b),
    .io_ci(FullAdder_1872_io_ci),
    .io_s(FullAdder_1872_io_s),
    .io_co(FullAdder_1872_io_co)
  );
  FullAdder FullAdder_1873 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1873_io_a),
    .io_b(FullAdder_1873_io_b),
    .io_ci(FullAdder_1873_io_ci),
    .io_s(FullAdder_1873_io_s),
    .io_co(FullAdder_1873_io_co)
  );
  FullAdder FullAdder_1874 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1874_io_a),
    .io_b(FullAdder_1874_io_b),
    .io_ci(FullAdder_1874_io_ci),
    .io_s(FullAdder_1874_io_s),
    .io_co(FullAdder_1874_io_co)
  );
  FullAdder FullAdder_1875 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1875_io_a),
    .io_b(FullAdder_1875_io_b),
    .io_ci(FullAdder_1875_io_ci),
    .io_s(FullAdder_1875_io_s),
    .io_co(FullAdder_1875_io_co)
  );
  FullAdder FullAdder_1876 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1876_io_a),
    .io_b(FullAdder_1876_io_b),
    .io_ci(FullAdder_1876_io_ci),
    .io_s(FullAdder_1876_io_s),
    .io_co(FullAdder_1876_io_co)
  );
  FullAdder FullAdder_1877 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1877_io_a),
    .io_b(FullAdder_1877_io_b),
    .io_ci(FullAdder_1877_io_ci),
    .io_s(FullAdder_1877_io_s),
    .io_co(FullAdder_1877_io_co)
  );
  FullAdder FullAdder_1878 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1878_io_a),
    .io_b(FullAdder_1878_io_b),
    .io_ci(FullAdder_1878_io_ci),
    .io_s(FullAdder_1878_io_s),
    .io_co(FullAdder_1878_io_co)
  );
  FullAdder FullAdder_1879 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1879_io_a),
    .io_b(FullAdder_1879_io_b),
    .io_ci(FullAdder_1879_io_ci),
    .io_s(FullAdder_1879_io_s),
    .io_co(FullAdder_1879_io_co)
  );
  FullAdder FullAdder_1880 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1880_io_a),
    .io_b(FullAdder_1880_io_b),
    .io_ci(FullAdder_1880_io_ci),
    .io_s(FullAdder_1880_io_s),
    .io_co(FullAdder_1880_io_co)
  );
  FullAdder FullAdder_1881 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1881_io_a),
    .io_b(FullAdder_1881_io_b),
    .io_ci(FullAdder_1881_io_ci),
    .io_s(FullAdder_1881_io_s),
    .io_co(FullAdder_1881_io_co)
  );
  FullAdder FullAdder_1882 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1882_io_a),
    .io_b(FullAdder_1882_io_b),
    .io_ci(FullAdder_1882_io_ci),
    .io_s(FullAdder_1882_io_s),
    .io_co(FullAdder_1882_io_co)
  );
  FullAdder FullAdder_1883 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1883_io_a),
    .io_b(FullAdder_1883_io_b),
    .io_ci(FullAdder_1883_io_ci),
    .io_s(FullAdder_1883_io_s),
    .io_co(FullAdder_1883_io_co)
  );
  FullAdder FullAdder_1884 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1884_io_a),
    .io_b(FullAdder_1884_io_b),
    .io_ci(FullAdder_1884_io_ci),
    .io_s(FullAdder_1884_io_s),
    .io_co(FullAdder_1884_io_co)
  );
  FullAdder FullAdder_1885 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1885_io_a),
    .io_b(FullAdder_1885_io_b),
    .io_ci(FullAdder_1885_io_ci),
    .io_s(FullAdder_1885_io_s),
    .io_co(FullAdder_1885_io_co)
  );
  FullAdder FullAdder_1886 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1886_io_a),
    .io_b(FullAdder_1886_io_b),
    .io_ci(FullAdder_1886_io_ci),
    .io_s(FullAdder_1886_io_s),
    .io_co(FullAdder_1886_io_co)
  );
  FullAdder FullAdder_1887 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1887_io_a),
    .io_b(FullAdder_1887_io_b),
    .io_ci(FullAdder_1887_io_ci),
    .io_s(FullAdder_1887_io_s),
    .io_co(FullAdder_1887_io_co)
  );
  FullAdder FullAdder_1888 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1888_io_a),
    .io_b(FullAdder_1888_io_b),
    .io_ci(FullAdder_1888_io_ci),
    .io_s(FullAdder_1888_io_s),
    .io_co(FullAdder_1888_io_co)
  );
  FullAdder FullAdder_1889 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1889_io_a),
    .io_b(FullAdder_1889_io_b),
    .io_ci(FullAdder_1889_io_ci),
    .io_s(FullAdder_1889_io_s),
    .io_co(FullAdder_1889_io_co)
  );
  FullAdder FullAdder_1890 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1890_io_a),
    .io_b(FullAdder_1890_io_b),
    .io_ci(FullAdder_1890_io_ci),
    .io_s(FullAdder_1890_io_s),
    .io_co(FullAdder_1890_io_co)
  );
  FullAdder FullAdder_1891 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1891_io_a),
    .io_b(FullAdder_1891_io_b),
    .io_ci(FullAdder_1891_io_ci),
    .io_s(FullAdder_1891_io_s),
    .io_co(FullAdder_1891_io_co)
  );
  FullAdder FullAdder_1892 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1892_io_a),
    .io_b(FullAdder_1892_io_b),
    .io_ci(FullAdder_1892_io_ci),
    .io_s(FullAdder_1892_io_s),
    .io_co(FullAdder_1892_io_co)
  );
  FullAdder FullAdder_1893 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1893_io_a),
    .io_b(FullAdder_1893_io_b),
    .io_ci(FullAdder_1893_io_ci),
    .io_s(FullAdder_1893_io_s),
    .io_co(FullAdder_1893_io_co)
  );
  FullAdder FullAdder_1894 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1894_io_a),
    .io_b(FullAdder_1894_io_b),
    .io_ci(FullAdder_1894_io_ci),
    .io_s(FullAdder_1894_io_s),
    .io_co(FullAdder_1894_io_co)
  );
  FullAdder FullAdder_1895 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1895_io_a),
    .io_b(FullAdder_1895_io_b),
    .io_ci(FullAdder_1895_io_ci),
    .io_s(FullAdder_1895_io_s),
    .io_co(FullAdder_1895_io_co)
  );
  FullAdder FullAdder_1896 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1896_io_a),
    .io_b(FullAdder_1896_io_b),
    .io_ci(FullAdder_1896_io_ci),
    .io_s(FullAdder_1896_io_s),
    .io_co(FullAdder_1896_io_co)
  );
  FullAdder FullAdder_1897 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1897_io_a),
    .io_b(FullAdder_1897_io_b),
    .io_ci(FullAdder_1897_io_ci),
    .io_s(FullAdder_1897_io_s),
    .io_co(FullAdder_1897_io_co)
  );
  FullAdder FullAdder_1898 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1898_io_a),
    .io_b(FullAdder_1898_io_b),
    .io_ci(FullAdder_1898_io_ci),
    .io_s(FullAdder_1898_io_s),
    .io_co(FullAdder_1898_io_co)
  );
  FullAdder FullAdder_1899 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1899_io_a),
    .io_b(FullAdder_1899_io_b),
    .io_ci(FullAdder_1899_io_ci),
    .io_s(FullAdder_1899_io_s),
    .io_co(FullAdder_1899_io_co)
  );
  FullAdder FullAdder_1900 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1900_io_a),
    .io_b(FullAdder_1900_io_b),
    .io_ci(FullAdder_1900_io_ci),
    .io_s(FullAdder_1900_io_s),
    .io_co(FullAdder_1900_io_co)
  );
  FullAdder FullAdder_1901 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1901_io_a),
    .io_b(FullAdder_1901_io_b),
    .io_ci(FullAdder_1901_io_ci),
    .io_s(FullAdder_1901_io_s),
    .io_co(FullAdder_1901_io_co)
  );
  FullAdder FullAdder_1902 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1902_io_a),
    .io_b(FullAdder_1902_io_b),
    .io_ci(FullAdder_1902_io_ci),
    .io_s(FullAdder_1902_io_s),
    .io_co(FullAdder_1902_io_co)
  );
  FullAdder FullAdder_1903 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1903_io_a),
    .io_b(FullAdder_1903_io_b),
    .io_ci(FullAdder_1903_io_ci),
    .io_s(FullAdder_1903_io_s),
    .io_co(FullAdder_1903_io_co)
  );
  FullAdder FullAdder_1904 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1904_io_a),
    .io_b(FullAdder_1904_io_b),
    .io_ci(FullAdder_1904_io_ci),
    .io_s(FullAdder_1904_io_s),
    .io_co(FullAdder_1904_io_co)
  );
  FullAdder FullAdder_1905 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1905_io_a),
    .io_b(FullAdder_1905_io_b),
    .io_ci(FullAdder_1905_io_ci),
    .io_s(FullAdder_1905_io_s),
    .io_co(FullAdder_1905_io_co)
  );
  FullAdder FullAdder_1906 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1906_io_a),
    .io_b(FullAdder_1906_io_b),
    .io_ci(FullAdder_1906_io_ci),
    .io_s(FullAdder_1906_io_s),
    .io_co(FullAdder_1906_io_co)
  );
  FullAdder FullAdder_1907 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1907_io_a),
    .io_b(FullAdder_1907_io_b),
    .io_ci(FullAdder_1907_io_ci),
    .io_s(FullAdder_1907_io_s),
    .io_co(FullAdder_1907_io_co)
  );
  FullAdder FullAdder_1908 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1908_io_a),
    .io_b(FullAdder_1908_io_b),
    .io_ci(FullAdder_1908_io_ci),
    .io_s(FullAdder_1908_io_s),
    .io_co(FullAdder_1908_io_co)
  );
  FullAdder FullAdder_1909 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1909_io_a),
    .io_b(FullAdder_1909_io_b),
    .io_ci(FullAdder_1909_io_ci),
    .io_s(FullAdder_1909_io_s),
    .io_co(FullAdder_1909_io_co)
  );
  FullAdder FullAdder_1910 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1910_io_a),
    .io_b(FullAdder_1910_io_b),
    .io_ci(FullAdder_1910_io_ci),
    .io_s(FullAdder_1910_io_s),
    .io_co(FullAdder_1910_io_co)
  );
  FullAdder FullAdder_1911 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1911_io_a),
    .io_b(FullAdder_1911_io_b),
    .io_ci(FullAdder_1911_io_ci),
    .io_s(FullAdder_1911_io_s),
    .io_co(FullAdder_1911_io_co)
  );
  FullAdder FullAdder_1912 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1912_io_a),
    .io_b(FullAdder_1912_io_b),
    .io_ci(FullAdder_1912_io_ci),
    .io_s(FullAdder_1912_io_s),
    .io_co(FullAdder_1912_io_co)
  );
  FullAdder FullAdder_1913 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1913_io_a),
    .io_b(FullAdder_1913_io_b),
    .io_ci(FullAdder_1913_io_ci),
    .io_s(FullAdder_1913_io_s),
    .io_co(FullAdder_1913_io_co)
  );
  FullAdder FullAdder_1914 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1914_io_a),
    .io_b(FullAdder_1914_io_b),
    .io_ci(FullAdder_1914_io_ci),
    .io_s(FullAdder_1914_io_s),
    .io_co(FullAdder_1914_io_co)
  );
  FullAdder FullAdder_1915 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1915_io_a),
    .io_b(FullAdder_1915_io_b),
    .io_ci(FullAdder_1915_io_ci),
    .io_s(FullAdder_1915_io_s),
    .io_co(FullAdder_1915_io_co)
  );
  FullAdder FullAdder_1916 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1916_io_a),
    .io_b(FullAdder_1916_io_b),
    .io_ci(FullAdder_1916_io_ci),
    .io_s(FullAdder_1916_io_s),
    .io_co(FullAdder_1916_io_co)
  );
  FullAdder FullAdder_1917 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1917_io_a),
    .io_b(FullAdder_1917_io_b),
    .io_ci(FullAdder_1917_io_ci),
    .io_s(FullAdder_1917_io_s),
    .io_co(FullAdder_1917_io_co)
  );
  FullAdder FullAdder_1918 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1918_io_a),
    .io_b(FullAdder_1918_io_b),
    .io_ci(FullAdder_1918_io_ci),
    .io_s(FullAdder_1918_io_s),
    .io_co(FullAdder_1918_io_co)
  );
  FullAdder FullAdder_1919 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1919_io_a),
    .io_b(FullAdder_1919_io_b),
    .io_ci(FullAdder_1919_io_ci),
    .io_s(FullAdder_1919_io_s),
    .io_co(FullAdder_1919_io_co)
  );
  FullAdder FullAdder_1920 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1920_io_a),
    .io_b(FullAdder_1920_io_b),
    .io_ci(FullAdder_1920_io_ci),
    .io_s(FullAdder_1920_io_s),
    .io_co(FullAdder_1920_io_co)
  );
  FullAdder FullAdder_1921 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1921_io_a),
    .io_b(FullAdder_1921_io_b),
    .io_ci(FullAdder_1921_io_ci),
    .io_s(FullAdder_1921_io_s),
    .io_co(FullAdder_1921_io_co)
  );
  FullAdder FullAdder_1922 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1922_io_a),
    .io_b(FullAdder_1922_io_b),
    .io_ci(FullAdder_1922_io_ci),
    .io_s(FullAdder_1922_io_s),
    .io_co(FullAdder_1922_io_co)
  );
  FullAdder FullAdder_1923 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1923_io_a),
    .io_b(FullAdder_1923_io_b),
    .io_ci(FullAdder_1923_io_ci),
    .io_s(FullAdder_1923_io_s),
    .io_co(FullAdder_1923_io_co)
  );
  FullAdder FullAdder_1924 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1924_io_a),
    .io_b(FullAdder_1924_io_b),
    .io_ci(FullAdder_1924_io_ci),
    .io_s(FullAdder_1924_io_s),
    .io_co(FullAdder_1924_io_co)
  );
  FullAdder FullAdder_1925 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1925_io_a),
    .io_b(FullAdder_1925_io_b),
    .io_ci(FullAdder_1925_io_ci),
    .io_s(FullAdder_1925_io_s),
    .io_co(FullAdder_1925_io_co)
  );
  HalfAdder HalfAdder_50 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_50_io_a),
    .io_b(HalfAdder_50_io_b),
    .io_s(HalfAdder_50_io_s),
    .io_co(HalfAdder_50_io_co)
  );
  FullAdder FullAdder_1926 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1926_io_a),
    .io_b(FullAdder_1926_io_b),
    .io_ci(FullAdder_1926_io_ci),
    .io_s(FullAdder_1926_io_s),
    .io_co(FullAdder_1926_io_co)
  );
  FullAdder FullAdder_1927 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1927_io_a),
    .io_b(FullAdder_1927_io_b),
    .io_ci(FullAdder_1927_io_ci),
    .io_s(FullAdder_1927_io_s),
    .io_co(FullAdder_1927_io_co)
  );
  FullAdder FullAdder_1928 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1928_io_a),
    .io_b(FullAdder_1928_io_b),
    .io_ci(FullAdder_1928_io_ci),
    .io_s(FullAdder_1928_io_s),
    .io_co(FullAdder_1928_io_co)
  );
  FullAdder FullAdder_1929 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1929_io_a),
    .io_b(FullAdder_1929_io_b),
    .io_ci(FullAdder_1929_io_ci),
    .io_s(FullAdder_1929_io_s),
    .io_co(FullAdder_1929_io_co)
  );
  FullAdder FullAdder_1930 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1930_io_a),
    .io_b(FullAdder_1930_io_b),
    .io_ci(FullAdder_1930_io_ci),
    .io_s(FullAdder_1930_io_s),
    .io_co(FullAdder_1930_io_co)
  );
  FullAdder FullAdder_1931 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1931_io_a),
    .io_b(FullAdder_1931_io_b),
    .io_ci(FullAdder_1931_io_ci),
    .io_s(FullAdder_1931_io_s),
    .io_co(FullAdder_1931_io_co)
  );
  FullAdder FullAdder_1932 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1932_io_a),
    .io_b(FullAdder_1932_io_b),
    .io_ci(FullAdder_1932_io_ci),
    .io_s(FullAdder_1932_io_s),
    .io_co(FullAdder_1932_io_co)
  );
  FullAdder FullAdder_1933 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1933_io_a),
    .io_b(FullAdder_1933_io_b),
    .io_ci(FullAdder_1933_io_ci),
    .io_s(FullAdder_1933_io_s),
    .io_co(FullAdder_1933_io_co)
  );
  FullAdder FullAdder_1934 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1934_io_a),
    .io_b(FullAdder_1934_io_b),
    .io_ci(FullAdder_1934_io_ci),
    .io_s(FullAdder_1934_io_s),
    .io_co(FullAdder_1934_io_co)
  );
  FullAdder FullAdder_1935 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1935_io_a),
    .io_b(FullAdder_1935_io_b),
    .io_ci(FullAdder_1935_io_ci),
    .io_s(FullAdder_1935_io_s),
    .io_co(FullAdder_1935_io_co)
  );
  FullAdder FullAdder_1936 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1936_io_a),
    .io_b(FullAdder_1936_io_b),
    .io_ci(FullAdder_1936_io_ci),
    .io_s(FullAdder_1936_io_s),
    .io_co(FullAdder_1936_io_co)
  );
  FullAdder FullAdder_1937 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1937_io_a),
    .io_b(FullAdder_1937_io_b),
    .io_ci(FullAdder_1937_io_ci),
    .io_s(FullAdder_1937_io_s),
    .io_co(FullAdder_1937_io_co)
  );
  FullAdder FullAdder_1938 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1938_io_a),
    .io_b(FullAdder_1938_io_b),
    .io_ci(FullAdder_1938_io_ci),
    .io_s(FullAdder_1938_io_s),
    .io_co(FullAdder_1938_io_co)
  );
  FullAdder FullAdder_1939 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1939_io_a),
    .io_b(FullAdder_1939_io_b),
    .io_ci(FullAdder_1939_io_ci),
    .io_s(FullAdder_1939_io_s),
    .io_co(FullAdder_1939_io_co)
  );
  FullAdder FullAdder_1940 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1940_io_a),
    .io_b(FullAdder_1940_io_b),
    .io_ci(FullAdder_1940_io_ci),
    .io_s(FullAdder_1940_io_s),
    .io_co(FullAdder_1940_io_co)
  );
  FullAdder FullAdder_1941 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1941_io_a),
    .io_b(FullAdder_1941_io_b),
    .io_ci(FullAdder_1941_io_ci),
    .io_s(FullAdder_1941_io_s),
    .io_co(FullAdder_1941_io_co)
  );
  FullAdder FullAdder_1942 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1942_io_a),
    .io_b(FullAdder_1942_io_b),
    .io_ci(FullAdder_1942_io_ci),
    .io_s(FullAdder_1942_io_s),
    .io_co(FullAdder_1942_io_co)
  );
  FullAdder FullAdder_1943 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1943_io_a),
    .io_b(FullAdder_1943_io_b),
    .io_ci(FullAdder_1943_io_ci),
    .io_s(FullAdder_1943_io_s),
    .io_co(FullAdder_1943_io_co)
  );
  FullAdder FullAdder_1944 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1944_io_a),
    .io_b(FullAdder_1944_io_b),
    .io_ci(FullAdder_1944_io_ci),
    .io_s(FullAdder_1944_io_s),
    .io_co(FullAdder_1944_io_co)
  );
  FullAdder FullAdder_1945 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1945_io_a),
    .io_b(FullAdder_1945_io_b),
    .io_ci(FullAdder_1945_io_ci),
    .io_s(FullAdder_1945_io_s),
    .io_co(FullAdder_1945_io_co)
  );
  FullAdder FullAdder_1946 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1946_io_a),
    .io_b(FullAdder_1946_io_b),
    .io_ci(FullAdder_1946_io_ci),
    .io_s(FullAdder_1946_io_s),
    .io_co(FullAdder_1946_io_co)
  );
  FullAdder FullAdder_1947 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1947_io_a),
    .io_b(FullAdder_1947_io_b),
    .io_ci(FullAdder_1947_io_ci),
    .io_s(FullAdder_1947_io_s),
    .io_co(FullAdder_1947_io_co)
  );
  FullAdder FullAdder_1948 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1948_io_a),
    .io_b(FullAdder_1948_io_b),
    .io_ci(FullAdder_1948_io_ci),
    .io_s(FullAdder_1948_io_s),
    .io_co(FullAdder_1948_io_co)
  );
  FullAdder FullAdder_1949 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1949_io_a),
    .io_b(FullAdder_1949_io_b),
    .io_ci(FullAdder_1949_io_ci),
    .io_s(FullAdder_1949_io_s),
    .io_co(FullAdder_1949_io_co)
  );
  FullAdder FullAdder_1950 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1950_io_a),
    .io_b(FullAdder_1950_io_b),
    .io_ci(FullAdder_1950_io_ci),
    .io_s(FullAdder_1950_io_s),
    .io_co(FullAdder_1950_io_co)
  );
  FullAdder FullAdder_1951 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1951_io_a),
    .io_b(FullAdder_1951_io_b),
    .io_ci(FullAdder_1951_io_ci),
    .io_s(FullAdder_1951_io_s),
    .io_co(FullAdder_1951_io_co)
  );
  FullAdder FullAdder_1952 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1952_io_a),
    .io_b(FullAdder_1952_io_b),
    .io_ci(FullAdder_1952_io_ci),
    .io_s(FullAdder_1952_io_s),
    .io_co(FullAdder_1952_io_co)
  );
  FullAdder FullAdder_1953 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1953_io_a),
    .io_b(FullAdder_1953_io_b),
    .io_ci(FullAdder_1953_io_ci),
    .io_s(FullAdder_1953_io_s),
    .io_co(FullAdder_1953_io_co)
  );
  FullAdder FullAdder_1954 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1954_io_a),
    .io_b(FullAdder_1954_io_b),
    .io_ci(FullAdder_1954_io_ci),
    .io_s(FullAdder_1954_io_s),
    .io_co(FullAdder_1954_io_co)
  );
  FullAdder FullAdder_1955 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1955_io_a),
    .io_b(FullAdder_1955_io_b),
    .io_ci(FullAdder_1955_io_ci),
    .io_s(FullAdder_1955_io_s),
    .io_co(FullAdder_1955_io_co)
  );
  FullAdder FullAdder_1956 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1956_io_a),
    .io_b(FullAdder_1956_io_b),
    .io_ci(FullAdder_1956_io_ci),
    .io_s(FullAdder_1956_io_s),
    .io_co(FullAdder_1956_io_co)
  );
  FullAdder FullAdder_1957 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1957_io_a),
    .io_b(FullAdder_1957_io_b),
    .io_ci(FullAdder_1957_io_ci),
    .io_s(FullAdder_1957_io_s),
    .io_co(FullAdder_1957_io_co)
  );
  FullAdder FullAdder_1958 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1958_io_a),
    .io_b(FullAdder_1958_io_b),
    .io_ci(FullAdder_1958_io_ci),
    .io_s(FullAdder_1958_io_s),
    .io_co(FullAdder_1958_io_co)
  );
  FullAdder FullAdder_1959 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1959_io_a),
    .io_b(FullAdder_1959_io_b),
    .io_ci(FullAdder_1959_io_ci),
    .io_s(FullAdder_1959_io_s),
    .io_co(FullAdder_1959_io_co)
  );
  FullAdder FullAdder_1960 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1960_io_a),
    .io_b(FullAdder_1960_io_b),
    .io_ci(FullAdder_1960_io_ci),
    .io_s(FullAdder_1960_io_s),
    .io_co(FullAdder_1960_io_co)
  );
  FullAdder FullAdder_1961 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1961_io_a),
    .io_b(FullAdder_1961_io_b),
    .io_ci(FullAdder_1961_io_ci),
    .io_s(FullAdder_1961_io_s),
    .io_co(FullAdder_1961_io_co)
  );
  FullAdder FullAdder_1962 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1962_io_a),
    .io_b(FullAdder_1962_io_b),
    .io_ci(FullAdder_1962_io_ci),
    .io_s(FullAdder_1962_io_s),
    .io_co(FullAdder_1962_io_co)
  );
  FullAdder FullAdder_1963 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1963_io_a),
    .io_b(FullAdder_1963_io_b),
    .io_ci(FullAdder_1963_io_ci),
    .io_s(FullAdder_1963_io_s),
    .io_co(FullAdder_1963_io_co)
  );
  FullAdder FullAdder_1964 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1964_io_a),
    .io_b(FullAdder_1964_io_b),
    .io_ci(FullAdder_1964_io_ci),
    .io_s(FullAdder_1964_io_s),
    .io_co(FullAdder_1964_io_co)
  );
  FullAdder FullAdder_1965 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1965_io_a),
    .io_b(FullAdder_1965_io_b),
    .io_ci(FullAdder_1965_io_ci),
    .io_s(FullAdder_1965_io_s),
    .io_co(FullAdder_1965_io_co)
  );
  FullAdder FullAdder_1966 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1966_io_a),
    .io_b(FullAdder_1966_io_b),
    .io_ci(FullAdder_1966_io_ci),
    .io_s(FullAdder_1966_io_s),
    .io_co(FullAdder_1966_io_co)
  );
  FullAdder FullAdder_1967 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1967_io_a),
    .io_b(FullAdder_1967_io_b),
    .io_ci(FullAdder_1967_io_ci),
    .io_s(FullAdder_1967_io_s),
    .io_co(FullAdder_1967_io_co)
  );
  FullAdder FullAdder_1968 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1968_io_a),
    .io_b(FullAdder_1968_io_b),
    .io_ci(FullAdder_1968_io_ci),
    .io_s(FullAdder_1968_io_s),
    .io_co(FullAdder_1968_io_co)
  );
  HalfAdder HalfAdder_51 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_51_io_a),
    .io_b(HalfAdder_51_io_b),
    .io_s(HalfAdder_51_io_s),
    .io_co(HalfAdder_51_io_co)
  );
  FullAdder FullAdder_1969 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1969_io_a),
    .io_b(FullAdder_1969_io_b),
    .io_ci(FullAdder_1969_io_ci),
    .io_s(FullAdder_1969_io_s),
    .io_co(FullAdder_1969_io_co)
  );
  FullAdder FullAdder_1970 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1970_io_a),
    .io_b(FullAdder_1970_io_b),
    .io_ci(FullAdder_1970_io_ci),
    .io_s(FullAdder_1970_io_s),
    .io_co(FullAdder_1970_io_co)
  );
  FullAdder FullAdder_1971 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1971_io_a),
    .io_b(FullAdder_1971_io_b),
    .io_ci(FullAdder_1971_io_ci),
    .io_s(FullAdder_1971_io_s),
    .io_co(FullAdder_1971_io_co)
  );
  FullAdder FullAdder_1972 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1972_io_a),
    .io_b(FullAdder_1972_io_b),
    .io_ci(FullAdder_1972_io_ci),
    .io_s(FullAdder_1972_io_s),
    .io_co(FullAdder_1972_io_co)
  );
  FullAdder FullAdder_1973 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1973_io_a),
    .io_b(FullAdder_1973_io_b),
    .io_ci(FullAdder_1973_io_ci),
    .io_s(FullAdder_1973_io_s),
    .io_co(FullAdder_1973_io_co)
  );
  FullAdder FullAdder_1974 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1974_io_a),
    .io_b(FullAdder_1974_io_b),
    .io_ci(FullAdder_1974_io_ci),
    .io_s(FullAdder_1974_io_s),
    .io_co(FullAdder_1974_io_co)
  );
  FullAdder FullAdder_1975 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1975_io_a),
    .io_b(FullAdder_1975_io_b),
    .io_ci(FullAdder_1975_io_ci),
    .io_s(FullAdder_1975_io_s),
    .io_co(FullAdder_1975_io_co)
  );
  FullAdder FullAdder_1976 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1976_io_a),
    .io_b(FullAdder_1976_io_b),
    .io_ci(FullAdder_1976_io_ci),
    .io_s(FullAdder_1976_io_s),
    .io_co(FullAdder_1976_io_co)
  );
  FullAdder FullAdder_1977 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1977_io_a),
    .io_b(FullAdder_1977_io_b),
    .io_ci(FullAdder_1977_io_ci),
    .io_s(FullAdder_1977_io_s),
    .io_co(FullAdder_1977_io_co)
  );
  FullAdder FullAdder_1978 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1978_io_a),
    .io_b(FullAdder_1978_io_b),
    .io_ci(FullAdder_1978_io_ci),
    .io_s(FullAdder_1978_io_s),
    .io_co(FullAdder_1978_io_co)
  );
  FullAdder FullAdder_1979 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1979_io_a),
    .io_b(FullAdder_1979_io_b),
    .io_ci(FullAdder_1979_io_ci),
    .io_s(FullAdder_1979_io_s),
    .io_co(FullAdder_1979_io_co)
  );
  FullAdder FullAdder_1980 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1980_io_a),
    .io_b(FullAdder_1980_io_b),
    .io_ci(FullAdder_1980_io_ci),
    .io_s(FullAdder_1980_io_s),
    .io_co(FullAdder_1980_io_co)
  );
  FullAdder FullAdder_1981 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1981_io_a),
    .io_b(FullAdder_1981_io_b),
    .io_ci(FullAdder_1981_io_ci),
    .io_s(FullAdder_1981_io_s),
    .io_co(FullAdder_1981_io_co)
  );
  FullAdder FullAdder_1982 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1982_io_a),
    .io_b(FullAdder_1982_io_b),
    .io_ci(FullAdder_1982_io_ci),
    .io_s(FullAdder_1982_io_s),
    .io_co(FullAdder_1982_io_co)
  );
  FullAdder FullAdder_1983 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1983_io_a),
    .io_b(FullAdder_1983_io_b),
    .io_ci(FullAdder_1983_io_ci),
    .io_s(FullAdder_1983_io_s),
    .io_co(FullAdder_1983_io_co)
  );
  FullAdder FullAdder_1984 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1984_io_a),
    .io_b(FullAdder_1984_io_b),
    .io_ci(FullAdder_1984_io_ci),
    .io_s(FullAdder_1984_io_s),
    .io_co(FullAdder_1984_io_co)
  );
  FullAdder FullAdder_1985 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1985_io_a),
    .io_b(FullAdder_1985_io_b),
    .io_ci(FullAdder_1985_io_ci),
    .io_s(FullAdder_1985_io_s),
    .io_co(FullAdder_1985_io_co)
  );
  FullAdder FullAdder_1986 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1986_io_a),
    .io_b(FullAdder_1986_io_b),
    .io_ci(FullAdder_1986_io_ci),
    .io_s(FullAdder_1986_io_s),
    .io_co(FullAdder_1986_io_co)
  );
  FullAdder FullAdder_1987 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1987_io_a),
    .io_b(FullAdder_1987_io_b),
    .io_ci(FullAdder_1987_io_ci),
    .io_s(FullAdder_1987_io_s),
    .io_co(FullAdder_1987_io_co)
  );
  FullAdder FullAdder_1988 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1988_io_a),
    .io_b(FullAdder_1988_io_b),
    .io_ci(FullAdder_1988_io_ci),
    .io_s(FullAdder_1988_io_s),
    .io_co(FullAdder_1988_io_co)
  );
  FullAdder FullAdder_1989 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1989_io_a),
    .io_b(FullAdder_1989_io_b),
    .io_ci(FullAdder_1989_io_ci),
    .io_s(FullAdder_1989_io_s),
    .io_co(FullAdder_1989_io_co)
  );
  FullAdder FullAdder_1990 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1990_io_a),
    .io_b(FullAdder_1990_io_b),
    .io_ci(FullAdder_1990_io_ci),
    .io_s(FullAdder_1990_io_s),
    .io_co(FullAdder_1990_io_co)
  );
  FullAdder FullAdder_1991 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1991_io_a),
    .io_b(FullAdder_1991_io_b),
    .io_ci(FullAdder_1991_io_ci),
    .io_s(FullAdder_1991_io_s),
    .io_co(FullAdder_1991_io_co)
  );
  FullAdder FullAdder_1992 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1992_io_a),
    .io_b(FullAdder_1992_io_b),
    .io_ci(FullAdder_1992_io_ci),
    .io_s(FullAdder_1992_io_s),
    .io_co(FullAdder_1992_io_co)
  );
  FullAdder FullAdder_1993 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1993_io_a),
    .io_b(FullAdder_1993_io_b),
    .io_ci(FullAdder_1993_io_ci),
    .io_s(FullAdder_1993_io_s),
    .io_co(FullAdder_1993_io_co)
  );
  FullAdder FullAdder_1994 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1994_io_a),
    .io_b(FullAdder_1994_io_b),
    .io_ci(FullAdder_1994_io_ci),
    .io_s(FullAdder_1994_io_s),
    .io_co(FullAdder_1994_io_co)
  );
  FullAdder FullAdder_1995 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1995_io_a),
    .io_b(FullAdder_1995_io_b),
    .io_ci(FullAdder_1995_io_ci),
    .io_s(FullAdder_1995_io_s),
    .io_co(FullAdder_1995_io_co)
  );
  FullAdder FullAdder_1996 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1996_io_a),
    .io_b(FullAdder_1996_io_b),
    .io_ci(FullAdder_1996_io_ci),
    .io_s(FullAdder_1996_io_s),
    .io_co(FullAdder_1996_io_co)
  );
  FullAdder FullAdder_1997 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1997_io_a),
    .io_b(FullAdder_1997_io_b),
    .io_ci(FullAdder_1997_io_ci),
    .io_s(FullAdder_1997_io_s),
    .io_co(FullAdder_1997_io_co)
  );
  FullAdder FullAdder_1998 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1998_io_a),
    .io_b(FullAdder_1998_io_b),
    .io_ci(FullAdder_1998_io_ci),
    .io_s(FullAdder_1998_io_s),
    .io_co(FullAdder_1998_io_co)
  );
  FullAdder FullAdder_1999 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_1999_io_a),
    .io_b(FullAdder_1999_io_b),
    .io_ci(FullAdder_1999_io_ci),
    .io_s(FullAdder_1999_io_s),
    .io_co(FullAdder_1999_io_co)
  );
  FullAdder FullAdder_2000 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2000_io_a),
    .io_b(FullAdder_2000_io_b),
    .io_ci(FullAdder_2000_io_ci),
    .io_s(FullAdder_2000_io_s),
    .io_co(FullAdder_2000_io_co)
  );
  FullAdder FullAdder_2001 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2001_io_a),
    .io_b(FullAdder_2001_io_b),
    .io_ci(FullAdder_2001_io_ci),
    .io_s(FullAdder_2001_io_s),
    .io_co(FullAdder_2001_io_co)
  );
  FullAdder FullAdder_2002 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2002_io_a),
    .io_b(FullAdder_2002_io_b),
    .io_ci(FullAdder_2002_io_ci),
    .io_s(FullAdder_2002_io_s),
    .io_co(FullAdder_2002_io_co)
  );
  FullAdder FullAdder_2003 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2003_io_a),
    .io_b(FullAdder_2003_io_b),
    .io_ci(FullAdder_2003_io_ci),
    .io_s(FullAdder_2003_io_s),
    .io_co(FullAdder_2003_io_co)
  );
  FullAdder FullAdder_2004 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2004_io_a),
    .io_b(FullAdder_2004_io_b),
    .io_ci(FullAdder_2004_io_ci),
    .io_s(FullAdder_2004_io_s),
    .io_co(FullAdder_2004_io_co)
  );
  FullAdder FullAdder_2005 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2005_io_a),
    .io_b(FullAdder_2005_io_b),
    .io_ci(FullAdder_2005_io_ci),
    .io_s(FullAdder_2005_io_s),
    .io_co(FullAdder_2005_io_co)
  );
  FullAdder FullAdder_2006 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2006_io_a),
    .io_b(FullAdder_2006_io_b),
    .io_ci(FullAdder_2006_io_ci),
    .io_s(FullAdder_2006_io_s),
    .io_co(FullAdder_2006_io_co)
  );
  FullAdder FullAdder_2007 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2007_io_a),
    .io_b(FullAdder_2007_io_b),
    .io_ci(FullAdder_2007_io_ci),
    .io_s(FullAdder_2007_io_s),
    .io_co(FullAdder_2007_io_co)
  );
  FullAdder FullAdder_2008 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2008_io_a),
    .io_b(FullAdder_2008_io_b),
    .io_ci(FullAdder_2008_io_ci),
    .io_s(FullAdder_2008_io_s),
    .io_co(FullAdder_2008_io_co)
  );
  FullAdder FullAdder_2009 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2009_io_a),
    .io_b(FullAdder_2009_io_b),
    .io_ci(FullAdder_2009_io_ci),
    .io_s(FullAdder_2009_io_s),
    .io_co(FullAdder_2009_io_co)
  );
  FullAdder FullAdder_2010 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2010_io_a),
    .io_b(FullAdder_2010_io_b),
    .io_ci(FullAdder_2010_io_ci),
    .io_s(FullAdder_2010_io_s),
    .io_co(FullAdder_2010_io_co)
  );
  FullAdder FullAdder_2011 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2011_io_a),
    .io_b(FullAdder_2011_io_b),
    .io_ci(FullAdder_2011_io_ci),
    .io_s(FullAdder_2011_io_s),
    .io_co(FullAdder_2011_io_co)
  );
  FullAdder FullAdder_2012 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2012_io_a),
    .io_b(FullAdder_2012_io_b),
    .io_ci(FullAdder_2012_io_ci),
    .io_s(FullAdder_2012_io_s),
    .io_co(FullAdder_2012_io_co)
  );
  FullAdder FullAdder_2013 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2013_io_a),
    .io_b(FullAdder_2013_io_b),
    .io_ci(FullAdder_2013_io_ci),
    .io_s(FullAdder_2013_io_s),
    .io_co(FullAdder_2013_io_co)
  );
  FullAdder FullAdder_2014 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2014_io_a),
    .io_b(FullAdder_2014_io_b),
    .io_ci(FullAdder_2014_io_ci),
    .io_s(FullAdder_2014_io_s),
    .io_co(FullAdder_2014_io_co)
  );
  FullAdder FullAdder_2015 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2015_io_a),
    .io_b(FullAdder_2015_io_b),
    .io_ci(FullAdder_2015_io_ci),
    .io_s(FullAdder_2015_io_s),
    .io_co(FullAdder_2015_io_co)
  );
  FullAdder FullAdder_2016 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2016_io_a),
    .io_b(FullAdder_2016_io_b),
    .io_ci(FullAdder_2016_io_ci),
    .io_s(FullAdder_2016_io_s),
    .io_co(FullAdder_2016_io_co)
  );
  HalfAdder HalfAdder_52 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_52_io_a),
    .io_b(HalfAdder_52_io_b),
    .io_s(HalfAdder_52_io_s),
    .io_co(HalfAdder_52_io_co)
  );
  FullAdder FullAdder_2017 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2017_io_a),
    .io_b(FullAdder_2017_io_b),
    .io_ci(FullAdder_2017_io_ci),
    .io_s(FullAdder_2017_io_s),
    .io_co(FullAdder_2017_io_co)
  );
  FullAdder FullAdder_2018 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2018_io_a),
    .io_b(FullAdder_2018_io_b),
    .io_ci(FullAdder_2018_io_ci),
    .io_s(FullAdder_2018_io_s),
    .io_co(FullAdder_2018_io_co)
  );
  FullAdder FullAdder_2019 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2019_io_a),
    .io_b(FullAdder_2019_io_b),
    .io_ci(FullAdder_2019_io_ci),
    .io_s(FullAdder_2019_io_s),
    .io_co(FullAdder_2019_io_co)
  );
  FullAdder FullAdder_2020 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2020_io_a),
    .io_b(FullAdder_2020_io_b),
    .io_ci(FullAdder_2020_io_ci),
    .io_s(FullAdder_2020_io_s),
    .io_co(FullAdder_2020_io_co)
  );
  FullAdder FullAdder_2021 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2021_io_a),
    .io_b(FullAdder_2021_io_b),
    .io_ci(FullAdder_2021_io_ci),
    .io_s(FullAdder_2021_io_s),
    .io_co(FullAdder_2021_io_co)
  );
  FullAdder FullAdder_2022 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2022_io_a),
    .io_b(FullAdder_2022_io_b),
    .io_ci(FullAdder_2022_io_ci),
    .io_s(FullAdder_2022_io_s),
    .io_co(FullAdder_2022_io_co)
  );
  FullAdder FullAdder_2023 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2023_io_a),
    .io_b(FullAdder_2023_io_b),
    .io_ci(FullAdder_2023_io_ci),
    .io_s(FullAdder_2023_io_s),
    .io_co(FullAdder_2023_io_co)
  );
  FullAdder FullAdder_2024 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2024_io_a),
    .io_b(FullAdder_2024_io_b),
    .io_ci(FullAdder_2024_io_ci),
    .io_s(FullAdder_2024_io_s),
    .io_co(FullAdder_2024_io_co)
  );
  FullAdder FullAdder_2025 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2025_io_a),
    .io_b(FullAdder_2025_io_b),
    .io_ci(FullAdder_2025_io_ci),
    .io_s(FullAdder_2025_io_s),
    .io_co(FullAdder_2025_io_co)
  );
  FullAdder FullAdder_2026 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2026_io_a),
    .io_b(FullAdder_2026_io_b),
    .io_ci(FullAdder_2026_io_ci),
    .io_s(FullAdder_2026_io_s),
    .io_co(FullAdder_2026_io_co)
  );
  FullAdder FullAdder_2027 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2027_io_a),
    .io_b(FullAdder_2027_io_b),
    .io_ci(FullAdder_2027_io_ci),
    .io_s(FullAdder_2027_io_s),
    .io_co(FullAdder_2027_io_co)
  );
  FullAdder FullAdder_2028 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2028_io_a),
    .io_b(FullAdder_2028_io_b),
    .io_ci(FullAdder_2028_io_ci),
    .io_s(FullAdder_2028_io_s),
    .io_co(FullAdder_2028_io_co)
  );
  FullAdder FullAdder_2029 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2029_io_a),
    .io_b(FullAdder_2029_io_b),
    .io_ci(FullAdder_2029_io_ci),
    .io_s(FullAdder_2029_io_s),
    .io_co(FullAdder_2029_io_co)
  );
  FullAdder FullAdder_2030 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2030_io_a),
    .io_b(FullAdder_2030_io_b),
    .io_ci(FullAdder_2030_io_ci),
    .io_s(FullAdder_2030_io_s),
    .io_co(FullAdder_2030_io_co)
  );
  FullAdder FullAdder_2031 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2031_io_a),
    .io_b(FullAdder_2031_io_b),
    .io_ci(FullAdder_2031_io_ci),
    .io_s(FullAdder_2031_io_s),
    .io_co(FullAdder_2031_io_co)
  );
  FullAdder FullAdder_2032 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2032_io_a),
    .io_b(FullAdder_2032_io_b),
    .io_ci(FullAdder_2032_io_ci),
    .io_s(FullAdder_2032_io_s),
    .io_co(FullAdder_2032_io_co)
  );
  FullAdder FullAdder_2033 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2033_io_a),
    .io_b(FullAdder_2033_io_b),
    .io_ci(FullAdder_2033_io_ci),
    .io_s(FullAdder_2033_io_s),
    .io_co(FullAdder_2033_io_co)
  );
  FullAdder FullAdder_2034 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2034_io_a),
    .io_b(FullAdder_2034_io_b),
    .io_ci(FullAdder_2034_io_ci),
    .io_s(FullAdder_2034_io_s),
    .io_co(FullAdder_2034_io_co)
  );
  FullAdder FullAdder_2035 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2035_io_a),
    .io_b(FullAdder_2035_io_b),
    .io_ci(FullAdder_2035_io_ci),
    .io_s(FullAdder_2035_io_s),
    .io_co(FullAdder_2035_io_co)
  );
  FullAdder FullAdder_2036 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2036_io_a),
    .io_b(FullAdder_2036_io_b),
    .io_ci(FullAdder_2036_io_ci),
    .io_s(FullAdder_2036_io_s),
    .io_co(FullAdder_2036_io_co)
  );
  FullAdder FullAdder_2037 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2037_io_a),
    .io_b(FullAdder_2037_io_b),
    .io_ci(FullAdder_2037_io_ci),
    .io_s(FullAdder_2037_io_s),
    .io_co(FullAdder_2037_io_co)
  );
  FullAdder FullAdder_2038 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2038_io_a),
    .io_b(FullAdder_2038_io_b),
    .io_ci(FullAdder_2038_io_ci),
    .io_s(FullAdder_2038_io_s),
    .io_co(FullAdder_2038_io_co)
  );
  FullAdder FullAdder_2039 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2039_io_a),
    .io_b(FullAdder_2039_io_b),
    .io_ci(FullAdder_2039_io_ci),
    .io_s(FullAdder_2039_io_s),
    .io_co(FullAdder_2039_io_co)
  );
  FullAdder FullAdder_2040 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2040_io_a),
    .io_b(FullAdder_2040_io_b),
    .io_ci(FullAdder_2040_io_ci),
    .io_s(FullAdder_2040_io_s),
    .io_co(FullAdder_2040_io_co)
  );
  FullAdder FullAdder_2041 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2041_io_a),
    .io_b(FullAdder_2041_io_b),
    .io_ci(FullAdder_2041_io_ci),
    .io_s(FullAdder_2041_io_s),
    .io_co(FullAdder_2041_io_co)
  );
  FullAdder FullAdder_2042 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2042_io_a),
    .io_b(FullAdder_2042_io_b),
    .io_ci(FullAdder_2042_io_ci),
    .io_s(FullAdder_2042_io_s),
    .io_co(FullAdder_2042_io_co)
  );
  FullAdder FullAdder_2043 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2043_io_a),
    .io_b(FullAdder_2043_io_b),
    .io_ci(FullAdder_2043_io_ci),
    .io_s(FullAdder_2043_io_s),
    .io_co(FullAdder_2043_io_co)
  );
  FullAdder FullAdder_2044 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2044_io_a),
    .io_b(FullAdder_2044_io_b),
    .io_ci(FullAdder_2044_io_ci),
    .io_s(FullAdder_2044_io_s),
    .io_co(FullAdder_2044_io_co)
  );
  FullAdder FullAdder_2045 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2045_io_a),
    .io_b(FullAdder_2045_io_b),
    .io_ci(FullAdder_2045_io_ci),
    .io_s(FullAdder_2045_io_s),
    .io_co(FullAdder_2045_io_co)
  );
  FullAdder FullAdder_2046 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2046_io_a),
    .io_b(FullAdder_2046_io_b),
    .io_ci(FullAdder_2046_io_ci),
    .io_s(FullAdder_2046_io_s),
    .io_co(FullAdder_2046_io_co)
  );
  FullAdder FullAdder_2047 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2047_io_a),
    .io_b(FullAdder_2047_io_b),
    .io_ci(FullAdder_2047_io_ci),
    .io_s(FullAdder_2047_io_s),
    .io_co(FullAdder_2047_io_co)
  );
  FullAdder FullAdder_2048 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2048_io_a),
    .io_b(FullAdder_2048_io_b),
    .io_ci(FullAdder_2048_io_ci),
    .io_s(FullAdder_2048_io_s),
    .io_co(FullAdder_2048_io_co)
  );
  FullAdder FullAdder_2049 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2049_io_a),
    .io_b(FullAdder_2049_io_b),
    .io_ci(FullAdder_2049_io_ci),
    .io_s(FullAdder_2049_io_s),
    .io_co(FullAdder_2049_io_co)
  );
  FullAdder FullAdder_2050 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2050_io_a),
    .io_b(FullAdder_2050_io_b),
    .io_ci(FullAdder_2050_io_ci),
    .io_s(FullAdder_2050_io_s),
    .io_co(FullAdder_2050_io_co)
  );
  FullAdder FullAdder_2051 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2051_io_a),
    .io_b(FullAdder_2051_io_b),
    .io_ci(FullAdder_2051_io_ci),
    .io_s(FullAdder_2051_io_s),
    .io_co(FullAdder_2051_io_co)
  );
  HalfAdder HalfAdder_53 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_53_io_a),
    .io_b(HalfAdder_53_io_b),
    .io_s(HalfAdder_53_io_s),
    .io_co(HalfAdder_53_io_co)
  );
  FullAdder FullAdder_2052 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2052_io_a),
    .io_b(FullAdder_2052_io_b),
    .io_ci(FullAdder_2052_io_ci),
    .io_s(FullAdder_2052_io_s),
    .io_co(FullAdder_2052_io_co)
  );
  FullAdder FullAdder_2053 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2053_io_a),
    .io_b(FullAdder_2053_io_b),
    .io_ci(FullAdder_2053_io_ci),
    .io_s(FullAdder_2053_io_s),
    .io_co(FullAdder_2053_io_co)
  );
  FullAdder FullAdder_2054 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2054_io_a),
    .io_b(FullAdder_2054_io_b),
    .io_ci(FullAdder_2054_io_ci),
    .io_s(FullAdder_2054_io_s),
    .io_co(FullAdder_2054_io_co)
  );
  FullAdder FullAdder_2055 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2055_io_a),
    .io_b(FullAdder_2055_io_b),
    .io_ci(FullAdder_2055_io_ci),
    .io_s(FullAdder_2055_io_s),
    .io_co(FullAdder_2055_io_co)
  );
  FullAdder FullAdder_2056 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2056_io_a),
    .io_b(FullAdder_2056_io_b),
    .io_ci(FullAdder_2056_io_ci),
    .io_s(FullAdder_2056_io_s),
    .io_co(FullAdder_2056_io_co)
  );
  FullAdder FullAdder_2057 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2057_io_a),
    .io_b(FullAdder_2057_io_b),
    .io_ci(FullAdder_2057_io_ci),
    .io_s(FullAdder_2057_io_s),
    .io_co(FullAdder_2057_io_co)
  );
  FullAdder FullAdder_2058 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2058_io_a),
    .io_b(FullAdder_2058_io_b),
    .io_ci(FullAdder_2058_io_ci),
    .io_s(FullAdder_2058_io_s),
    .io_co(FullAdder_2058_io_co)
  );
  FullAdder FullAdder_2059 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2059_io_a),
    .io_b(FullAdder_2059_io_b),
    .io_ci(FullAdder_2059_io_ci),
    .io_s(FullAdder_2059_io_s),
    .io_co(FullAdder_2059_io_co)
  );
  FullAdder FullAdder_2060 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2060_io_a),
    .io_b(FullAdder_2060_io_b),
    .io_ci(FullAdder_2060_io_ci),
    .io_s(FullAdder_2060_io_s),
    .io_co(FullAdder_2060_io_co)
  );
  FullAdder FullAdder_2061 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2061_io_a),
    .io_b(FullAdder_2061_io_b),
    .io_ci(FullAdder_2061_io_ci),
    .io_s(FullAdder_2061_io_s),
    .io_co(FullAdder_2061_io_co)
  );
  FullAdder FullAdder_2062 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2062_io_a),
    .io_b(FullAdder_2062_io_b),
    .io_ci(FullAdder_2062_io_ci),
    .io_s(FullAdder_2062_io_s),
    .io_co(FullAdder_2062_io_co)
  );
  FullAdder FullAdder_2063 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2063_io_a),
    .io_b(FullAdder_2063_io_b),
    .io_ci(FullAdder_2063_io_ci),
    .io_s(FullAdder_2063_io_s),
    .io_co(FullAdder_2063_io_co)
  );
  FullAdder FullAdder_2064 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2064_io_a),
    .io_b(FullAdder_2064_io_b),
    .io_ci(FullAdder_2064_io_ci),
    .io_s(FullAdder_2064_io_s),
    .io_co(FullAdder_2064_io_co)
  );
  FullAdder FullAdder_2065 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2065_io_a),
    .io_b(FullAdder_2065_io_b),
    .io_ci(FullAdder_2065_io_ci),
    .io_s(FullAdder_2065_io_s),
    .io_co(FullAdder_2065_io_co)
  );
  FullAdder FullAdder_2066 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2066_io_a),
    .io_b(FullAdder_2066_io_b),
    .io_ci(FullAdder_2066_io_ci),
    .io_s(FullAdder_2066_io_s),
    .io_co(FullAdder_2066_io_co)
  );
  FullAdder FullAdder_2067 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2067_io_a),
    .io_b(FullAdder_2067_io_b),
    .io_ci(FullAdder_2067_io_ci),
    .io_s(FullAdder_2067_io_s),
    .io_co(FullAdder_2067_io_co)
  );
  FullAdder FullAdder_2068 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2068_io_a),
    .io_b(FullAdder_2068_io_b),
    .io_ci(FullAdder_2068_io_ci),
    .io_s(FullAdder_2068_io_s),
    .io_co(FullAdder_2068_io_co)
  );
  FullAdder FullAdder_2069 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2069_io_a),
    .io_b(FullAdder_2069_io_b),
    .io_ci(FullAdder_2069_io_ci),
    .io_s(FullAdder_2069_io_s),
    .io_co(FullAdder_2069_io_co)
  );
  FullAdder FullAdder_2070 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2070_io_a),
    .io_b(FullAdder_2070_io_b),
    .io_ci(FullAdder_2070_io_ci),
    .io_s(FullAdder_2070_io_s),
    .io_co(FullAdder_2070_io_co)
  );
  FullAdder FullAdder_2071 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2071_io_a),
    .io_b(FullAdder_2071_io_b),
    .io_ci(FullAdder_2071_io_ci),
    .io_s(FullAdder_2071_io_s),
    .io_co(FullAdder_2071_io_co)
  );
  FullAdder FullAdder_2072 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2072_io_a),
    .io_b(FullAdder_2072_io_b),
    .io_ci(FullAdder_2072_io_ci),
    .io_s(FullAdder_2072_io_s),
    .io_co(FullAdder_2072_io_co)
  );
  FullAdder FullAdder_2073 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2073_io_a),
    .io_b(FullAdder_2073_io_b),
    .io_ci(FullAdder_2073_io_ci),
    .io_s(FullAdder_2073_io_s),
    .io_co(FullAdder_2073_io_co)
  );
  FullAdder FullAdder_2074 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2074_io_a),
    .io_b(FullAdder_2074_io_b),
    .io_ci(FullAdder_2074_io_ci),
    .io_s(FullAdder_2074_io_s),
    .io_co(FullAdder_2074_io_co)
  );
  FullAdder FullAdder_2075 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2075_io_a),
    .io_b(FullAdder_2075_io_b),
    .io_ci(FullAdder_2075_io_ci),
    .io_s(FullAdder_2075_io_s),
    .io_co(FullAdder_2075_io_co)
  );
  FullAdder FullAdder_2076 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2076_io_a),
    .io_b(FullAdder_2076_io_b),
    .io_ci(FullAdder_2076_io_ci),
    .io_s(FullAdder_2076_io_s),
    .io_co(FullAdder_2076_io_co)
  );
  FullAdder FullAdder_2077 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2077_io_a),
    .io_b(FullAdder_2077_io_b),
    .io_ci(FullAdder_2077_io_ci),
    .io_s(FullAdder_2077_io_s),
    .io_co(FullAdder_2077_io_co)
  );
  FullAdder FullAdder_2078 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2078_io_a),
    .io_b(FullAdder_2078_io_b),
    .io_ci(FullAdder_2078_io_ci),
    .io_s(FullAdder_2078_io_s),
    .io_co(FullAdder_2078_io_co)
  );
  FullAdder FullAdder_2079 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2079_io_a),
    .io_b(FullAdder_2079_io_b),
    .io_ci(FullAdder_2079_io_ci),
    .io_s(FullAdder_2079_io_s),
    .io_co(FullAdder_2079_io_co)
  );
  FullAdder FullAdder_2080 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2080_io_a),
    .io_b(FullAdder_2080_io_b),
    .io_ci(FullAdder_2080_io_ci),
    .io_s(FullAdder_2080_io_s),
    .io_co(FullAdder_2080_io_co)
  );
  FullAdder FullAdder_2081 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2081_io_a),
    .io_b(FullAdder_2081_io_b),
    .io_ci(FullAdder_2081_io_ci),
    .io_s(FullAdder_2081_io_s),
    .io_co(FullAdder_2081_io_co)
  );
  FullAdder FullAdder_2082 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2082_io_a),
    .io_b(FullAdder_2082_io_b),
    .io_ci(FullAdder_2082_io_ci),
    .io_s(FullAdder_2082_io_s),
    .io_co(FullAdder_2082_io_co)
  );
  FullAdder FullAdder_2083 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2083_io_a),
    .io_b(FullAdder_2083_io_b),
    .io_ci(FullAdder_2083_io_ci),
    .io_s(FullAdder_2083_io_s),
    .io_co(FullAdder_2083_io_co)
  );
  FullAdder FullAdder_2084 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2084_io_a),
    .io_b(FullAdder_2084_io_b),
    .io_ci(FullAdder_2084_io_ci),
    .io_s(FullAdder_2084_io_s),
    .io_co(FullAdder_2084_io_co)
  );
  FullAdder FullAdder_2085 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2085_io_a),
    .io_b(FullAdder_2085_io_b),
    .io_ci(FullAdder_2085_io_ci),
    .io_s(FullAdder_2085_io_s),
    .io_co(FullAdder_2085_io_co)
  );
  FullAdder FullAdder_2086 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2086_io_a),
    .io_b(FullAdder_2086_io_b),
    .io_ci(FullAdder_2086_io_ci),
    .io_s(FullAdder_2086_io_s),
    .io_co(FullAdder_2086_io_co)
  );
  FullAdder FullAdder_2087 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2087_io_a),
    .io_b(FullAdder_2087_io_b),
    .io_ci(FullAdder_2087_io_ci),
    .io_s(FullAdder_2087_io_s),
    .io_co(FullAdder_2087_io_co)
  );
  FullAdder FullAdder_2088 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2088_io_a),
    .io_b(FullAdder_2088_io_b),
    .io_ci(FullAdder_2088_io_ci),
    .io_s(FullAdder_2088_io_s),
    .io_co(FullAdder_2088_io_co)
  );
  FullAdder FullAdder_2089 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2089_io_a),
    .io_b(FullAdder_2089_io_b),
    .io_ci(FullAdder_2089_io_ci),
    .io_s(FullAdder_2089_io_s),
    .io_co(FullAdder_2089_io_co)
  );
  HalfAdder HalfAdder_54 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_54_io_a),
    .io_b(HalfAdder_54_io_b),
    .io_s(HalfAdder_54_io_s),
    .io_co(HalfAdder_54_io_co)
  );
  FullAdder FullAdder_2090 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2090_io_a),
    .io_b(FullAdder_2090_io_b),
    .io_ci(FullAdder_2090_io_ci),
    .io_s(FullAdder_2090_io_s),
    .io_co(FullAdder_2090_io_co)
  );
  FullAdder FullAdder_2091 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2091_io_a),
    .io_b(FullAdder_2091_io_b),
    .io_ci(FullAdder_2091_io_ci),
    .io_s(FullAdder_2091_io_s),
    .io_co(FullAdder_2091_io_co)
  );
  FullAdder FullAdder_2092 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2092_io_a),
    .io_b(FullAdder_2092_io_b),
    .io_ci(FullAdder_2092_io_ci),
    .io_s(FullAdder_2092_io_s),
    .io_co(FullAdder_2092_io_co)
  );
  FullAdder FullAdder_2093 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2093_io_a),
    .io_b(FullAdder_2093_io_b),
    .io_ci(FullAdder_2093_io_ci),
    .io_s(FullAdder_2093_io_s),
    .io_co(FullAdder_2093_io_co)
  );
  FullAdder FullAdder_2094 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2094_io_a),
    .io_b(FullAdder_2094_io_b),
    .io_ci(FullAdder_2094_io_ci),
    .io_s(FullAdder_2094_io_s),
    .io_co(FullAdder_2094_io_co)
  );
  FullAdder FullAdder_2095 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2095_io_a),
    .io_b(FullAdder_2095_io_b),
    .io_ci(FullAdder_2095_io_ci),
    .io_s(FullAdder_2095_io_s),
    .io_co(FullAdder_2095_io_co)
  );
  FullAdder FullAdder_2096 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2096_io_a),
    .io_b(FullAdder_2096_io_b),
    .io_ci(FullAdder_2096_io_ci),
    .io_s(FullAdder_2096_io_s),
    .io_co(FullAdder_2096_io_co)
  );
  FullAdder FullAdder_2097 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2097_io_a),
    .io_b(FullAdder_2097_io_b),
    .io_ci(FullAdder_2097_io_ci),
    .io_s(FullAdder_2097_io_s),
    .io_co(FullAdder_2097_io_co)
  );
  FullAdder FullAdder_2098 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2098_io_a),
    .io_b(FullAdder_2098_io_b),
    .io_ci(FullAdder_2098_io_ci),
    .io_s(FullAdder_2098_io_s),
    .io_co(FullAdder_2098_io_co)
  );
  FullAdder FullAdder_2099 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2099_io_a),
    .io_b(FullAdder_2099_io_b),
    .io_ci(FullAdder_2099_io_ci),
    .io_s(FullAdder_2099_io_s),
    .io_co(FullAdder_2099_io_co)
  );
  FullAdder FullAdder_2100 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2100_io_a),
    .io_b(FullAdder_2100_io_b),
    .io_ci(FullAdder_2100_io_ci),
    .io_s(FullAdder_2100_io_s),
    .io_co(FullAdder_2100_io_co)
  );
  FullAdder FullAdder_2101 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2101_io_a),
    .io_b(FullAdder_2101_io_b),
    .io_ci(FullAdder_2101_io_ci),
    .io_s(FullAdder_2101_io_s),
    .io_co(FullAdder_2101_io_co)
  );
  FullAdder FullAdder_2102 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2102_io_a),
    .io_b(FullAdder_2102_io_b),
    .io_ci(FullAdder_2102_io_ci),
    .io_s(FullAdder_2102_io_s),
    .io_co(FullAdder_2102_io_co)
  );
  FullAdder FullAdder_2103 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2103_io_a),
    .io_b(FullAdder_2103_io_b),
    .io_ci(FullAdder_2103_io_ci),
    .io_s(FullAdder_2103_io_s),
    .io_co(FullAdder_2103_io_co)
  );
  FullAdder FullAdder_2104 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2104_io_a),
    .io_b(FullAdder_2104_io_b),
    .io_ci(FullAdder_2104_io_ci),
    .io_s(FullAdder_2104_io_s),
    .io_co(FullAdder_2104_io_co)
  );
  FullAdder FullAdder_2105 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2105_io_a),
    .io_b(FullAdder_2105_io_b),
    .io_ci(FullAdder_2105_io_ci),
    .io_s(FullAdder_2105_io_s),
    .io_co(FullAdder_2105_io_co)
  );
  FullAdder FullAdder_2106 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2106_io_a),
    .io_b(FullAdder_2106_io_b),
    .io_ci(FullAdder_2106_io_ci),
    .io_s(FullAdder_2106_io_s),
    .io_co(FullAdder_2106_io_co)
  );
  FullAdder FullAdder_2107 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2107_io_a),
    .io_b(FullAdder_2107_io_b),
    .io_ci(FullAdder_2107_io_ci),
    .io_s(FullAdder_2107_io_s),
    .io_co(FullAdder_2107_io_co)
  );
  FullAdder FullAdder_2108 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2108_io_a),
    .io_b(FullAdder_2108_io_b),
    .io_ci(FullAdder_2108_io_ci),
    .io_s(FullAdder_2108_io_s),
    .io_co(FullAdder_2108_io_co)
  );
  FullAdder FullAdder_2109 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2109_io_a),
    .io_b(FullAdder_2109_io_b),
    .io_ci(FullAdder_2109_io_ci),
    .io_s(FullAdder_2109_io_s),
    .io_co(FullAdder_2109_io_co)
  );
  FullAdder FullAdder_2110 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2110_io_a),
    .io_b(FullAdder_2110_io_b),
    .io_ci(FullAdder_2110_io_ci),
    .io_s(FullAdder_2110_io_s),
    .io_co(FullAdder_2110_io_co)
  );
  FullAdder FullAdder_2111 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2111_io_a),
    .io_b(FullAdder_2111_io_b),
    .io_ci(FullAdder_2111_io_ci),
    .io_s(FullAdder_2111_io_s),
    .io_co(FullAdder_2111_io_co)
  );
  FullAdder FullAdder_2112 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2112_io_a),
    .io_b(FullAdder_2112_io_b),
    .io_ci(FullAdder_2112_io_ci),
    .io_s(FullAdder_2112_io_s),
    .io_co(FullAdder_2112_io_co)
  );
  FullAdder FullAdder_2113 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2113_io_a),
    .io_b(FullAdder_2113_io_b),
    .io_ci(FullAdder_2113_io_ci),
    .io_s(FullAdder_2113_io_s),
    .io_co(FullAdder_2113_io_co)
  );
  FullAdder FullAdder_2114 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2114_io_a),
    .io_b(FullAdder_2114_io_b),
    .io_ci(FullAdder_2114_io_ci),
    .io_s(FullAdder_2114_io_s),
    .io_co(FullAdder_2114_io_co)
  );
  FullAdder FullAdder_2115 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2115_io_a),
    .io_b(FullAdder_2115_io_b),
    .io_ci(FullAdder_2115_io_ci),
    .io_s(FullAdder_2115_io_s),
    .io_co(FullAdder_2115_io_co)
  );
  FullAdder FullAdder_2116 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2116_io_a),
    .io_b(FullAdder_2116_io_b),
    .io_ci(FullAdder_2116_io_ci),
    .io_s(FullAdder_2116_io_s),
    .io_co(FullAdder_2116_io_co)
  );
  HalfAdder HalfAdder_55 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_55_io_a),
    .io_b(HalfAdder_55_io_b),
    .io_s(HalfAdder_55_io_s),
    .io_co(HalfAdder_55_io_co)
  );
  FullAdder FullAdder_2117 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2117_io_a),
    .io_b(FullAdder_2117_io_b),
    .io_ci(FullAdder_2117_io_ci),
    .io_s(FullAdder_2117_io_s),
    .io_co(FullAdder_2117_io_co)
  );
  FullAdder FullAdder_2118 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2118_io_a),
    .io_b(FullAdder_2118_io_b),
    .io_ci(FullAdder_2118_io_ci),
    .io_s(FullAdder_2118_io_s),
    .io_co(FullAdder_2118_io_co)
  );
  FullAdder FullAdder_2119 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2119_io_a),
    .io_b(FullAdder_2119_io_b),
    .io_ci(FullAdder_2119_io_ci),
    .io_s(FullAdder_2119_io_s),
    .io_co(FullAdder_2119_io_co)
  );
  FullAdder FullAdder_2120 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2120_io_a),
    .io_b(FullAdder_2120_io_b),
    .io_ci(FullAdder_2120_io_ci),
    .io_s(FullAdder_2120_io_s),
    .io_co(FullAdder_2120_io_co)
  );
  FullAdder FullAdder_2121 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2121_io_a),
    .io_b(FullAdder_2121_io_b),
    .io_ci(FullAdder_2121_io_ci),
    .io_s(FullAdder_2121_io_s),
    .io_co(FullAdder_2121_io_co)
  );
  FullAdder FullAdder_2122 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2122_io_a),
    .io_b(FullAdder_2122_io_b),
    .io_ci(FullAdder_2122_io_ci),
    .io_s(FullAdder_2122_io_s),
    .io_co(FullAdder_2122_io_co)
  );
  FullAdder FullAdder_2123 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2123_io_a),
    .io_b(FullAdder_2123_io_b),
    .io_ci(FullAdder_2123_io_ci),
    .io_s(FullAdder_2123_io_s),
    .io_co(FullAdder_2123_io_co)
  );
  FullAdder FullAdder_2124 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2124_io_a),
    .io_b(FullAdder_2124_io_b),
    .io_ci(FullAdder_2124_io_ci),
    .io_s(FullAdder_2124_io_s),
    .io_co(FullAdder_2124_io_co)
  );
  FullAdder FullAdder_2125 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2125_io_a),
    .io_b(FullAdder_2125_io_b),
    .io_ci(FullAdder_2125_io_ci),
    .io_s(FullAdder_2125_io_s),
    .io_co(FullAdder_2125_io_co)
  );
  FullAdder FullAdder_2126 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2126_io_a),
    .io_b(FullAdder_2126_io_b),
    .io_ci(FullAdder_2126_io_ci),
    .io_s(FullAdder_2126_io_s),
    .io_co(FullAdder_2126_io_co)
  );
  FullAdder FullAdder_2127 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2127_io_a),
    .io_b(FullAdder_2127_io_b),
    .io_ci(FullAdder_2127_io_ci),
    .io_s(FullAdder_2127_io_s),
    .io_co(FullAdder_2127_io_co)
  );
  FullAdder FullAdder_2128 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2128_io_a),
    .io_b(FullAdder_2128_io_b),
    .io_ci(FullAdder_2128_io_ci),
    .io_s(FullAdder_2128_io_s),
    .io_co(FullAdder_2128_io_co)
  );
  FullAdder FullAdder_2129 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2129_io_a),
    .io_b(FullAdder_2129_io_b),
    .io_ci(FullAdder_2129_io_ci),
    .io_s(FullAdder_2129_io_s),
    .io_co(FullAdder_2129_io_co)
  );
  FullAdder FullAdder_2130 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2130_io_a),
    .io_b(FullAdder_2130_io_b),
    .io_ci(FullAdder_2130_io_ci),
    .io_s(FullAdder_2130_io_s),
    .io_co(FullAdder_2130_io_co)
  );
  FullAdder FullAdder_2131 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2131_io_a),
    .io_b(FullAdder_2131_io_b),
    .io_ci(FullAdder_2131_io_ci),
    .io_s(FullAdder_2131_io_s),
    .io_co(FullAdder_2131_io_co)
  );
  FullAdder FullAdder_2132 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2132_io_a),
    .io_b(FullAdder_2132_io_b),
    .io_ci(FullAdder_2132_io_ci),
    .io_s(FullAdder_2132_io_s),
    .io_co(FullAdder_2132_io_co)
  );
  FullAdder FullAdder_2133 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2133_io_a),
    .io_b(FullAdder_2133_io_b),
    .io_ci(FullAdder_2133_io_ci),
    .io_s(FullAdder_2133_io_s),
    .io_co(FullAdder_2133_io_co)
  );
  HalfAdder HalfAdder_56 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_56_io_a),
    .io_b(HalfAdder_56_io_b),
    .io_s(HalfAdder_56_io_s),
    .io_co(HalfAdder_56_io_co)
  );
  FullAdder FullAdder_2134 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2134_io_a),
    .io_b(FullAdder_2134_io_b),
    .io_ci(FullAdder_2134_io_ci),
    .io_s(FullAdder_2134_io_s),
    .io_co(FullAdder_2134_io_co)
  );
  FullAdder FullAdder_2135 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2135_io_a),
    .io_b(FullAdder_2135_io_b),
    .io_ci(FullAdder_2135_io_ci),
    .io_s(FullAdder_2135_io_s),
    .io_co(FullAdder_2135_io_co)
  );
  FullAdder FullAdder_2136 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2136_io_a),
    .io_b(FullAdder_2136_io_b),
    .io_ci(FullAdder_2136_io_ci),
    .io_s(FullAdder_2136_io_s),
    .io_co(FullAdder_2136_io_co)
  );
  FullAdder FullAdder_2137 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2137_io_a),
    .io_b(FullAdder_2137_io_b),
    .io_ci(FullAdder_2137_io_ci),
    .io_s(FullAdder_2137_io_s),
    .io_co(FullAdder_2137_io_co)
  );
  FullAdder FullAdder_2138 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2138_io_a),
    .io_b(FullAdder_2138_io_b),
    .io_ci(FullAdder_2138_io_ci),
    .io_s(FullAdder_2138_io_s),
    .io_co(FullAdder_2138_io_co)
  );
  FullAdder FullAdder_2139 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2139_io_a),
    .io_b(FullAdder_2139_io_b),
    .io_ci(FullAdder_2139_io_ci),
    .io_s(FullAdder_2139_io_s),
    .io_co(FullAdder_2139_io_co)
  );
  FullAdder FullAdder_2140 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2140_io_a),
    .io_b(FullAdder_2140_io_b),
    .io_ci(FullAdder_2140_io_ci),
    .io_s(FullAdder_2140_io_s),
    .io_co(FullAdder_2140_io_co)
  );
  FullAdder FullAdder_2141 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2141_io_a),
    .io_b(FullAdder_2141_io_b),
    .io_ci(FullAdder_2141_io_ci),
    .io_s(FullAdder_2141_io_s),
    .io_co(FullAdder_2141_io_co)
  );
  FullAdder FullAdder_2142 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2142_io_a),
    .io_b(FullAdder_2142_io_b),
    .io_ci(FullAdder_2142_io_ci),
    .io_s(FullAdder_2142_io_s),
    .io_co(FullAdder_2142_io_co)
  );
  FullAdder FullAdder_2143 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2143_io_a),
    .io_b(FullAdder_2143_io_b),
    .io_ci(FullAdder_2143_io_ci),
    .io_s(FullAdder_2143_io_s),
    .io_co(FullAdder_2143_io_co)
  );
  FullAdder FullAdder_2144 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2144_io_a),
    .io_b(FullAdder_2144_io_b),
    .io_ci(FullAdder_2144_io_ci),
    .io_s(FullAdder_2144_io_s),
    .io_co(FullAdder_2144_io_co)
  );
  FullAdder FullAdder_2145 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2145_io_a),
    .io_b(FullAdder_2145_io_b),
    .io_ci(FullAdder_2145_io_ci),
    .io_s(FullAdder_2145_io_s),
    .io_co(FullAdder_2145_io_co)
  );
  FullAdder FullAdder_2146 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2146_io_a),
    .io_b(FullAdder_2146_io_b),
    .io_ci(FullAdder_2146_io_ci),
    .io_s(FullAdder_2146_io_s),
    .io_co(FullAdder_2146_io_co)
  );
  FullAdder FullAdder_2147 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2147_io_a),
    .io_b(FullAdder_2147_io_b),
    .io_ci(FullAdder_2147_io_ci),
    .io_s(FullAdder_2147_io_s),
    .io_co(FullAdder_2147_io_co)
  );
  FullAdder FullAdder_2148 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2148_io_a),
    .io_b(FullAdder_2148_io_b),
    .io_ci(FullAdder_2148_io_ci),
    .io_s(FullAdder_2148_io_s),
    .io_co(FullAdder_2148_io_co)
  );
  FullAdder FullAdder_2149 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2149_io_a),
    .io_b(FullAdder_2149_io_b),
    .io_ci(FullAdder_2149_io_ci),
    .io_s(FullAdder_2149_io_s),
    .io_co(FullAdder_2149_io_co)
  );
  FullAdder FullAdder_2150 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2150_io_a),
    .io_b(FullAdder_2150_io_b),
    .io_ci(FullAdder_2150_io_ci),
    .io_s(FullAdder_2150_io_s),
    .io_co(FullAdder_2150_io_co)
  );
  FullAdder FullAdder_2151 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2151_io_a),
    .io_b(FullAdder_2151_io_b),
    .io_ci(FullAdder_2151_io_ci),
    .io_s(FullAdder_2151_io_s),
    .io_co(FullAdder_2151_io_co)
  );
  FullAdder FullAdder_2152 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2152_io_a),
    .io_b(FullAdder_2152_io_b),
    .io_ci(FullAdder_2152_io_ci),
    .io_s(FullAdder_2152_io_s),
    .io_co(FullAdder_2152_io_co)
  );
  FullAdder FullAdder_2153 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2153_io_a),
    .io_b(FullAdder_2153_io_b),
    .io_ci(FullAdder_2153_io_ci),
    .io_s(FullAdder_2153_io_s),
    .io_co(FullAdder_2153_io_co)
  );
  FullAdder FullAdder_2154 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2154_io_a),
    .io_b(FullAdder_2154_io_b),
    .io_ci(FullAdder_2154_io_ci),
    .io_s(FullAdder_2154_io_s),
    .io_co(FullAdder_2154_io_co)
  );
  FullAdder FullAdder_2155 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2155_io_a),
    .io_b(FullAdder_2155_io_b),
    .io_ci(FullAdder_2155_io_ci),
    .io_s(FullAdder_2155_io_s),
    .io_co(FullAdder_2155_io_co)
  );
  FullAdder FullAdder_2156 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2156_io_a),
    .io_b(FullAdder_2156_io_b),
    .io_ci(FullAdder_2156_io_ci),
    .io_s(FullAdder_2156_io_s),
    .io_co(FullAdder_2156_io_co)
  );
  FullAdder FullAdder_2157 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2157_io_a),
    .io_b(FullAdder_2157_io_b),
    .io_ci(FullAdder_2157_io_ci),
    .io_s(FullAdder_2157_io_s),
    .io_co(FullAdder_2157_io_co)
  );
  FullAdder FullAdder_2158 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2158_io_a),
    .io_b(FullAdder_2158_io_b),
    .io_ci(FullAdder_2158_io_ci),
    .io_s(FullAdder_2158_io_s),
    .io_co(FullAdder_2158_io_co)
  );
  FullAdder FullAdder_2159 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2159_io_a),
    .io_b(FullAdder_2159_io_b),
    .io_ci(FullAdder_2159_io_ci),
    .io_s(FullAdder_2159_io_s),
    .io_co(FullAdder_2159_io_co)
  );
  FullAdder FullAdder_2160 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2160_io_a),
    .io_b(FullAdder_2160_io_b),
    .io_ci(FullAdder_2160_io_ci),
    .io_s(FullAdder_2160_io_s),
    .io_co(FullAdder_2160_io_co)
  );
  FullAdder FullAdder_2161 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2161_io_a),
    .io_b(FullAdder_2161_io_b),
    .io_ci(FullAdder_2161_io_ci),
    .io_s(FullAdder_2161_io_s),
    .io_co(FullAdder_2161_io_co)
  );
  FullAdder FullAdder_2162 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2162_io_a),
    .io_b(FullAdder_2162_io_b),
    .io_ci(FullAdder_2162_io_ci),
    .io_s(FullAdder_2162_io_s),
    .io_co(FullAdder_2162_io_co)
  );
  FullAdder FullAdder_2163 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2163_io_a),
    .io_b(FullAdder_2163_io_b),
    .io_ci(FullAdder_2163_io_ci),
    .io_s(FullAdder_2163_io_s),
    .io_co(FullAdder_2163_io_co)
  );
  HalfAdder HalfAdder_57 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_57_io_a),
    .io_b(HalfAdder_57_io_b),
    .io_s(HalfAdder_57_io_s),
    .io_co(HalfAdder_57_io_co)
  );
  FullAdder FullAdder_2164 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2164_io_a),
    .io_b(FullAdder_2164_io_b),
    .io_ci(FullAdder_2164_io_ci),
    .io_s(FullAdder_2164_io_s),
    .io_co(FullAdder_2164_io_co)
  );
  FullAdder FullAdder_2165 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2165_io_a),
    .io_b(FullAdder_2165_io_b),
    .io_ci(FullAdder_2165_io_ci),
    .io_s(FullAdder_2165_io_s),
    .io_co(FullAdder_2165_io_co)
  );
  FullAdder FullAdder_2166 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2166_io_a),
    .io_b(FullAdder_2166_io_b),
    .io_ci(FullAdder_2166_io_ci),
    .io_s(FullAdder_2166_io_s),
    .io_co(FullAdder_2166_io_co)
  );
  FullAdder FullAdder_2167 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2167_io_a),
    .io_b(FullAdder_2167_io_b),
    .io_ci(FullAdder_2167_io_ci),
    .io_s(FullAdder_2167_io_s),
    .io_co(FullAdder_2167_io_co)
  );
  FullAdder FullAdder_2168 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2168_io_a),
    .io_b(FullAdder_2168_io_b),
    .io_ci(FullAdder_2168_io_ci),
    .io_s(FullAdder_2168_io_s),
    .io_co(FullAdder_2168_io_co)
  );
  FullAdder FullAdder_2169 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2169_io_a),
    .io_b(FullAdder_2169_io_b),
    .io_ci(FullAdder_2169_io_ci),
    .io_s(FullAdder_2169_io_s),
    .io_co(FullAdder_2169_io_co)
  );
  FullAdder FullAdder_2170 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2170_io_a),
    .io_b(FullAdder_2170_io_b),
    .io_ci(FullAdder_2170_io_ci),
    .io_s(FullAdder_2170_io_s),
    .io_co(FullAdder_2170_io_co)
  );
  FullAdder FullAdder_2171 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2171_io_a),
    .io_b(FullAdder_2171_io_b),
    .io_ci(FullAdder_2171_io_ci),
    .io_s(FullAdder_2171_io_s),
    .io_co(FullAdder_2171_io_co)
  );
  FullAdder FullAdder_2172 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2172_io_a),
    .io_b(FullAdder_2172_io_b),
    .io_ci(FullAdder_2172_io_ci),
    .io_s(FullAdder_2172_io_s),
    .io_co(FullAdder_2172_io_co)
  );
  FullAdder FullAdder_2173 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2173_io_a),
    .io_b(FullAdder_2173_io_b),
    .io_ci(FullAdder_2173_io_ci),
    .io_s(FullAdder_2173_io_s),
    .io_co(FullAdder_2173_io_co)
  );
  FullAdder FullAdder_2174 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2174_io_a),
    .io_b(FullAdder_2174_io_b),
    .io_ci(FullAdder_2174_io_ci),
    .io_s(FullAdder_2174_io_s),
    .io_co(FullAdder_2174_io_co)
  );
  FullAdder FullAdder_2175 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2175_io_a),
    .io_b(FullAdder_2175_io_b),
    .io_ci(FullAdder_2175_io_ci),
    .io_s(FullAdder_2175_io_s),
    .io_co(FullAdder_2175_io_co)
  );
  FullAdder FullAdder_2176 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2176_io_a),
    .io_b(FullAdder_2176_io_b),
    .io_ci(FullAdder_2176_io_ci),
    .io_s(FullAdder_2176_io_s),
    .io_co(FullAdder_2176_io_co)
  );
  FullAdder FullAdder_2177 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2177_io_a),
    .io_b(FullAdder_2177_io_b),
    .io_ci(FullAdder_2177_io_ci),
    .io_s(FullAdder_2177_io_s),
    .io_co(FullAdder_2177_io_co)
  );
  FullAdder FullAdder_2178 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2178_io_a),
    .io_b(FullAdder_2178_io_b),
    .io_ci(FullAdder_2178_io_ci),
    .io_s(FullAdder_2178_io_s),
    .io_co(FullAdder_2178_io_co)
  );
  HalfAdder HalfAdder_58 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_58_io_a),
    .io_b(HalfAdder_58_io_b),
    .io_s(HalfAdder_58_io_s),
    .io_co(HalfAdder_58_io_co)
  );
  FullAdder FullAdder_2179 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2179_io_a),
    .io_b(FullAdder_2179_io_b),
    .io_ci(FullAdder_2179_io_ci),
    .io_s(FullAdder_2179_io_s),
    .io_co(FullAdder_2179_io_co)
  );
  FullAdder FullAdder_2180 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2180_io_a),
    .io_b(FullAdder_2180_io_b),
    .io_ci(FullAdder_2180_io_ci),
    .io_s(FullAdder_2180_io_s),
    .io_co(FullAdder_2180_io_co)
  );
  FullAdder FullAdder_2181 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2181_io_a),
    .io_b(FullAdder_2181_io_b),
    .io_ci(FullAdder_2181_io_ci),
    .io_s(FullAdder_2181_io_s),
    .io_co(FullAdder_2181_io_co)
  );
  HalfAdder HalfAdder_59 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_59_io_a),
    .io_b(HalfAdder_59_io_b),
    .io_s(HalfAdder_59_io_s),
    .io_co(HalfAdder_59_io_co)
  );
  FullAdder FullAdder_2182 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2182_io_a),
    .io_b(FullAdder_2182_io_b),
    .io_ci(FullAdder_2182_io_ci),
    .io_s(FullAdder_2182_io_s),
    .io_co(FullAdder_2182_io_co)
  );
  FullAdder FullAdder_2183 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2183_io_a),
    .io_b(FullAdder_2183_io_b),
    .io_ci(FullAdder_2183_io_ci),
    .io_s(FullAdder_2183_io_s),
    .io_co(FullAdder_2183_io_co)
  );
  FullAdder FullAdder_2184 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2184_io_a),
    .io_b(FullAdder_2184_io_b),
    .io_ci(FullAdder_2184_io_ci),
    .io_s(FullAdder_2184_io_s),
    .io_co(FullAdder_2184_io_co)
  );
  FullAdder FullAdder_2185 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2185_io_a),
    .io_b(FullAdder_2185_io_b),
    .io_ci(FullAdder_2185_io_ci),
    .io_s(FullAdder_2185_io_s),
    .io_co(FullAdder_2185_io_co)
  );
  FullAdder FullAdder_2186 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2186_io_a),
    .io_b(FullAdder_2186_io_b),
    .io_ci(FullAdder_2186_io_ci),
    .io_s(FullAdder_2186_io_s),
    .io_co(FullAdder_2186_io_co)
  );
  FullAdder FullAdder_2187 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2187_io_a),
    .io_b(FullAdder_2187_io_b),
    .io_ci(FullAdder_2187_io_ci),
    .io_s(FullAdder_2187_io_s),
    .io_co(FullAdder_2187_io_co)
  );
  FullAdder FullAdder_2188 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2188_io_a),
    .io_b(FullAdder_2188_io_b),
    .io_ci(FullAdder_2188_io_ci),
    .io_s(FullAdder_2188_io_s),
    .io_co(FullAdder_2188_io_co)
  );
  FullAdder FullAdder_2189 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2189_io_a),
    .io_b(FullAdder_2189_io_b),
    .io_ci(FullAdder_2189_io_ci),
    .io_s(FullAdder_2189_io_s),
    .io_co(FullAdder_2189_io_co)
  );
  FullAdder FullAdder_2190 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2190_io_a),
    .io_b(FullAdder_2190_io_b),
    .io_ci(FullAdder_2190_io_ci),
    .io_s(FullAdder_2190_io_s),
    .io_co(FullAdder_2190_io_co)
  );
  FullAdder FullAdder_2191 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2191_io_a),
    .io_b(FullAdder_2191_io_b),
    .io_ci(FullAdder_2191_io_ci),
    .io_s(FullAdder_2191_io_s),
    .io_co(FullAdder_2191_io_co)
  );
  FullAdder FullAdder_2192 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2192_io_a),
    .io_b(FullAdder_2192_io_b),
    .io_ci(FullAdder_2192_io_ci),
    .io_s(FullAdder_2192_io_s),
    .io_co(FullAdder_2192_io_co)
  );
  FullAdder FullAdder_2193 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2193_io_a),
    .io_b(FullAdder_2193_io_b),
    .io_ci(FullAdder_2193_io_ci),
    .io_s(FullAdder_2193_io_s),
    .io_co(FullAdder_2193_io_co)
  );
  HalfAdder HalfAdder_60 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_60_io_a),
    .io_b(HalfAdder_60_io_b),
    .io_s(HalfAdder_60_io_s),
    .io_co(HalfAdder_60_io_co)
  );
  HalfAdder HalfAdder_61 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_61_io_a),
    .io_b(HalfAdder_61_io_b),
    .io_s(HalfAdder_61_io_s),
    .io_co(HalfAdder_61_io_co)
  );
  FullAdder FullAdder_2194 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2194_io_a),
    .io_b(FullAdder_2194_io_b),
    .io_ci(FullAdder_2194_io_ci),
    .io_s(FullAdder_2194_io_s),
    .io_co(FullAdder_2194_io_co)
  );
  FullAdder FullAdder_2195 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2195_io_a),
    .io_b(FullAdder_2195_io_b),
    .io_ci(FullAdder_2195_io_ci),
    .io_s(FullAdder_2195_io_s),
    .io_co(FullAdder_2195_io_co)
  );
  FullAdder FullAdder_2196 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2196_io_a),
    .io_b(FullAdder_2196_io_b),
    .io_ci(FullAdder_2196_io_ci),
    .io_s(FullAdder_2196_io_s),
    .io_co(FullAdder_2196_io_co)
  );
  FullAdder FullAdder_2197 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2197_io_a),
    .io_b(FullAdder_2197_io_b),
    .io_ci(FullAdder_2197_io_ci),
    .io_s(FullAdder_2197_io_s),
    .io_co(FullAdder_2197_io_co)
  );
  FullAdder FullAdder_2198 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2198_io_a),
    .io_b(FullAdder_2198_io_b),
    .io_ci(FullAdder_2198_io_ci),
    .io_s(FullAdder_2198_io_s),
    .io_co(FullAdder_2198_io_co)
  );
  HalfAdder HalfAdder_62 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_62_io_a),
    .io_b(HalfAdder_62_io_b),
    .io_s(HalfAdder_62_io_s),
    .io_co(HalfAdder_62_io_co)
  );
  FullAdder FullAdder_2199 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2199_io_a),
    .io_b(FullAdder_2199_io_b),
    .io_ci(FullAdder_2199_io_ci),
    .io_s(FullAdder_2199_io_s),
    .io_co(FullAdder_2199_io_co)
  );
  HalfAdder HalfAdder_63 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_63_io_a),
    .io_b(HalfAdder_63_io_b),
    .io_s(HalfAdder_63_io_s),
    .io_co(HalfAdder_63_io_co)
  );
  FullAdder FullAdder_2200 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2200_io_a),
    .io_b(FullAdder_2200_io_b),
    .io_ci(FullAdder_2200_io_ci),
    .io_s(FullAdder_2200_io_s),
    .io_co(FullAdder_2200_io_co)
  );
  HalfAdder HalfAdder_64 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_64_io_a),
    .io_b(HalfAdder_64_io_b),
    .io_s(HalfAdder_64_io_s),
    .io_co(HalfAdder_64_io_co)
  );
  FullAdder FullAdder_2201 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2201_io_a),
    .io_b(FullAdder_2201_io_b),
    .io_ci(FullAdder_2201_io_ci),
    .io_s(FullAdder_2201_io_s),
    .io_co(FullAdder_2201_io_co)
  );
  HalfAdder HalfAdder_65 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_65_io_a),
    .io_b(HalfAdder_65_io_b),
    .io_s(HalfAdder_65_io_s),
    .io_co(HalfAdder_65_io_co)
  );
  HalfAdder HalfAdder_66 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_66_io_a),
    .io_b(HalfAdder_66_io_b),
    .io_s(HalfAdder_66_io_s),
    .io_co(HalfAdder_66_io_co)
  );
  HalfAdder HalfAdder_67 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_67_io_a),
    .io_b(HalfAdder_67_io_b),
    .io_s(HalfAdder_67_io_s),
    .io_co(HalfAdder_67_io_co)
  );
  HalfAdder HalfAdder_68 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_68_io_a),
    .io_b(HalfAdder_68_io_b),
    .io_s(HalfAdder_68_io_s),
    .io_co(HalfAdder_68_io_co)
  );
  HalfAdder HalfAdder_69 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_69_io_a),
    .io_b(HalfAdder_69_io_b),
    .io_s(HalfAdder_69_io_s),
    .io_co(HalfAdder_69_io_co)
  );
  FullAdder FullAdder_2202 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2202_io_a),
    .io_b(FullAdder_2202_io_b),
    .io_ci(FullAdder_2202_io_ci),
    .io_s(FullAdder_2202_io_s),
    .io_co(FullAdder_2202_io_co)
  );
  FullAdder FullAdder_2203 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2203_io_a),
    .io_b(FullAdder_2203_io_b),
    .io_ci(FullAdder_2203_io_ci),
    .io_s(FullAdder_2203_io_s),
    .io_co(FullAdder_2203_io_co)
  );
  HalfAdder HalfAdder_70 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_70_io_a),
    .io_b(HalfAdder_70_io_b),
    .io_s(HalfAdder_70_io_s),
    .io_co(HalfAdder_70_io_co)
  );
  HalfAdder HalfAdder_71 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_71_io_a),
    .io_b(HalfAdder_71_io_b),
    .io_s(HalfAdder_71_io_s),
    .io_co(HalfAdder_71_io_co)
  );
  FullAdder FullAdder_2204 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2204_io_a),
    .io_b(FullAdder_2204_io_b),
    .io_ci(FullAdder_2204_io_ci),
    .io_s(FullAdder_2204_io_s),
    .io_co(FullAdder_2204_io_co)
  );
  FullAdder FullAdder_2205 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2205_io_a),
    .io_b(FullAdder_2205_io_b),
    .io_ci(FullAdder_2205_io_ci),
    .io_s(FullAdder_2205_io_s),
    .io_co(FullAdder_2205_io_co)
  );
  FullAdder FullAdder_2206 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2206_io_a),
    .io_b(FullAdder_2206_io_b),
    .io_ci(FullAdder_2206_io_ci),
    .io_s(FullAdder_2206_io_s),
    .io_co(FullAdder_2206_io_co)
  );
  FullAdder FullAdder_2207 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2207_io_a),
    .io_b(FullAdder_2207_io_b),
    .io_ci(FullAdder_2207_io_ci),
    .io_s(FullAdder_2207_io_s),
    .io_co(FullAdder_2207_io_co)
  );
  FullAdder FullAdder_2208 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2208_io_a),
    .io_b(FullAdder_2208_io_b),
    .io_ci(FullAdder_2208_io_ci),
    .io_s(FullAdder_2208_io_s),
    .io_co(FullAdder_2208_io_co)
  );
  FullAdder FullAdder_2209 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2209_io_a),
    .io_b(FullAdder_2209_io_b),
    .io_ci(FullAdder_2209_io_ci),
    .io_s(FullAdder_2209_io_s),
    .io_co(FullAdder_2209_io_co)
  );
  FullAdder FullAdder_2210 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2210_io_a),
    .io_b(FullAdder_2210_io_b),
    .io_ci(FullAdder_2210_io_ci),
    .io_s(FullAdder_2210_io_s),
    .io_co(FullAdder_2210_io_co)
  );
  FullAdder FullAdder_2211 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2211_io_a),
    .io_b(FullAdder_2211_io_b),
    .io_ci(FullAdder_2211_io_ci),
    .io_s(FullAdder_2211_io_s),
    .io_co(FullAdder_2211_io_co)
  );
  FullAdder FullAdder_2212 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2212_io_a),
    .io_b(FullAdder_2212_io_b),
    .io_ci(FullAdder_2212_io_ci),
    .io_s(FullAdder_2212_io_s),
    .io_co(FullAdder_2212_io_co)
  );
  FullAdder FullAdder_2213 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2213_io_a),
    .io_b(FullAdder_2213_io_b),
    .io_ci(FullAdder_2213_io_ci),
    .io_s(FullAdder_2213_io_s),
    .io_co(FullAdder_2213_io_co)
  );
  FullAdder FullAdder_2214 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2214_io_a),
    .io_b(FullAdder_2214_io_b),
    .io_ci(FullAdder_2214_io_ci),
    .io_s(FullAdder_2214_io_s),
    .io_co(FullAdder_2214_io_co)
  );
  FullAdder FullAdder_2215 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2215_io_a),
    .io_b(FullAdder_2215_io_b),
    .io_ci(FullAdder_2215_io_ci),
    .io_s(FullAdder_2215_io_s),
    .io_co(FullAdder_2215_io_co)
  );
  FullAdder FullAdder_2216 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2216_io_a),
    .io_b(FullAdder_2216_io_b),
    .io_ci(FullAdder_2216_io_ci),
    .io_s(FullAdder_2216_io_s),
    .io_co(FullAdder_2216_io_co)
  );
  FullAdder FullAdder_2217 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2217_io_a),
    .io_b(FullAdder_2217_io_b),
    .io_ci(FullAdder_2217_io_ci),
    .io_s(FullAdder_2217_io_s),
    .io_co(FullAdder_2217_io_co)
  );
  HalfAdder HalfAdder_72 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_72_io_a),
    .io_b(HalfAdder_72_io_b),
    .io_s(HalfAdder_72_io_s),
    .io_co(HalfAdder_72_io_co)
  );
  FullAdder FullAdder_2218 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2218_io_a),
    .io_b(FullAdder_2218_io_b),
    .io_ci(FullAdder_2218_io_ci),
    .io_s(FullAdder_2218_io_s),
    .io_co(FullAdder_2218_io_co)
  );
  FullAdder FullAdder_2219 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2219_io_a),
    .io_b(FullAdder_2219_io_b),
    .io_ci(FullAdder_2219_io_ci),
    .io_s(FullAdder_2219_io_s),
    .io_co(FullAdder_2219_io_co)
  );
  FullAdder FullAdder_2220 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2220_io_a),
    .io_b(FullAdder_2220_io_b),
    .io_ci(FullAdder_2220_io_ci),
    .io_s(FullAdder_2220_io_s),
    .io_co(FullAdder_2220_io_co)
  );
  FullAdder FullAdder_2221 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2221_io_a),
    .io_b(FullAdder_2221_io_b),
    .io_ci(FullAdder_2221_io_ci),
    .io_s(FullAdder_2221_io_s),
    .io_co(FullAdder_2221_io_co)
  );
  HalfAdder HalfAdder_73 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_73_io_a),
    .io_b(HalfAdder_73_io_b),
    .io_s(HalfAdder_73_io_s),
    .io_co(HalfAdder_73_io_co)
  );
  FullAdder FullAdder_2222 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2222_io_a),
    .io_b(FullAdder_2222_io_b),
    .io_ci(FullAdder_2222_io_ci),
    .io_s(FullAdder_2222_io_s),
    .io_co(FullAdder_2222_io_co)
  );
  FullAdder FullAdder_2223 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2223_io_a),
    .io_b(FullAdder_2223_io_b),
    .io_ci(FullAdder_2223_io_ci),
    .io_s(FullAdder_2223_io_s),
    .io_co(FullAdder_2223_io_co)
  );
  FullAdder FullAdder_2224 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2224_io_a),
    .io_b(FullAdder_2224_io_b),
    .io_ci(FullAdder_2224_io_ci),
    .io_s(FullAdder_2224_io_s),
    .io_co(FullAdder_2224_io_co)
  );
  FullAdder FullAdder_2225 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2225_io_a),
    .io_b(FullAdder_2225_io_b),
    .io_ci(FullAdder_2225_io_ci),
    .io_s(FullAdder_2225_io_s),
    .io_co(FullAdder_2225_io_co)
  );
  FullAdder FullAdder_2226 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2226_io_a),
    .io_b(FullAdder_2226_io_b),
    .io_ci(FullAdder_2226_io_ci),
    .io_s(FullAdder_2226_io_s),
    .io_co(FullAdder_2226_io_co)
  );
  FullAdder FullAdder_2227 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2227_io_a),
    .io_b(FullAdder_2227_io_b),
    .io_ci(FullAdder_2227_io_ci),
    .io_s(FullAdder_2227_io_s),
    .io_co(FullAdder_2227_io_co)
  );
  FullAdder FullAdder_2228 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2228_io_a),
    .io_b(FullAdder_2228_io_b),
    .io_ci(FullAdder_2228_io_ci),
    .io_s(FullAdder_2228_io_s),
    .io_co(FullAdder_2228_io_co)
  );
  FullAdder FullAdder_2229 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2229_io_a),
    .io_b(FullAdder_2229_io_b),
    .io_ci(FullAdder_2229_io_ci),
    .io_s(FullAdder_2229_io_s),
    .io_co(FullAdder_2229_io_co)
  );
  FullAdder FullAdder_2230 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2230_io_a),
    .io_b(FullAdder_2230_io_b),
    .io_ci(FullAdder_2230_io_ci),
    .io_s(FullAdder_2230_io_s),
    .io_co(FullAdder_2230_io_co)
  );
  FullAdder FullAdder_2231 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2231_io_a),
    .io_b(FullAdder_2231_io_b),
    .io_ci(FullAdder_2231_io_ci),
    .io_s(FullAdder_2231_io_s),
    .io_co(FullAdder_2231_io_co)
  );
  FullAdder FullAdder_2232 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2232_io_a),
    .io_b(FullAdder_2232_io_b),
    .io_ci(FullAdder_2232_io_ci),
    .io_s(FullAdder_2232_io_s),
    .io_co(FullAdder_2232_io_co)
  );
  FullAdder FullAdder_2233 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2233_io_a),
    .io_b(FullAdder_2233_io_b),
    .io_ci(FullAdder_2233_io_ci),
    .io_s(FullAdder_2233_io_s),
    .io_co(FullAdder_2233_io_co)
  );
  FullAdder FullAdder_2234 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2234_io_a),
    .io_b(FullAdder_2234_io_b),
    .io_ci(FullAdder_2234_io_ci),
    .io_s(FullAdder_2234_io_s),
    .io_co(FullAdder_2234_io_co)
  );
  FullAdder FullAdder_2235 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2235_io_a),
    .io_b(FullAdder_2235_io_b),
    .io_ci(FullAdder_2235_io_ci),
    .io_s(FullAdder_2235_io_s),
    .io_co(FullAdder_2235_io_co)
  );
  FullAdder FullAdder_2236 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2236_io_a),
    .io_b(FullAdder_2236_io_b),
    .io_ci(FullAdder_2236_io_ci),
    .io_s(FullAdder_2236_io_s),
    .io_co(FullAdder_2236_io_co)
  );
  FullAdder FullAdder_2237 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2237_io_a),
    .io_b(FullAdder_2237_io_b),
    .io_ci(FullAdder_2237_io_ci),
    .io_s(FullAdder_2237_io_s),
    .io_co(FullAdder_2237_io_co)
  );
  FullAdder FullAdder_2238 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2238_io_a),
    .io_b(FullAdder_2238_io_b),
    .io_ci(FullAdder_2238_io_ci),
    .io_s(FullAdder_2238_io_s),
    .io_co(FullAdder_2238_io_co)
  );
  FullAdder FullAdder_2239 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2239_io_a),
    .io_b(FullAdder_2239_io_b),
    .io_ci(FullAdder_2239_io_ci),
    .io_s(FullAdder_2239_io_s),
    .io_co(FullAdder_2239_io_co)
  );
  HalfAdder HalfAdder_74 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_74_io_a),
    .io_b(HalfAdder_74_io_b),
    .io_s(HalfAdder_74_io_s),
    .io_co(HalfAdder_74_io_co)
  );
  FullAdder FullAdder_2240 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2240_io_a),
    .io_b(FullAdder_2240_io_b),
    .io_ci(FullAdder_2240_io_ci),
    .io_s(FullAdder_2240_io_s),
    .io_co(FullAdder_2240_io_co)
  );
  FullAdder FullAdder_2241 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2241_io_a),
    .io_b(FullAdder_2241_io_b),
    .io_ci(FullAdder_2241_io_ci),
    .io_s(FullAdder_2241_io_s),
    .io_co(FullAdder_2241_io_co)
  );
  FullAdder FullAdder_2242 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2242_io_a),
    .io_b(FullAdder_2242_io_b),
    .io_ci(FullAdder_2242_io_ci),
    .io_s(FullAdder_2242_io_s),
    .io_co(FullAdder_2242_io_co)
  );
  FullAdder FullAdder_2243 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2243_io_a),
    .io_b(FullAdder_2243_io_b),
    .io_ci(FullAdder_2243_io_ci),
    .io_s(FullAdder_2243_io_s),
    .io_co(FullAdder_2243_io_co)
  );
  FullAdder FullAdder_2244 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2244_io_a),
    .io_b(FullAdder_2244_io_b),
    .io_ci(FullAdder_2244_io_ci),
    .io_s(FullAdder_2244_io_s),
    .io_co(FullAdder_2244_io_co)
  );
  FullAdder FullAdder_2245 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2245_io_a),
    .io_b(FullAdder_2245_io_b),
    .io_ci(FullAdder_2245_io_ci),
    .io_s(FullAdder_2245_io_s),
    .io_co(FullAdder_2245_io_co)
  );
  FullAdder FullAdder_2246 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2246_io_a),
    .io_b(FullAdder_2246_io_b),
    .io_ci(FullAdder_2246_io_ci),
    .io_s(FullAdder_2246_io_s),
    .io_co(FullAdder_2246_io_co)
  );
  FullAdder FullAdder_2247 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2247_io_a),
    .io_b(FullAdder_2247_io_b),
    .io_ci(FullAdder_2247_io_ci),
    .io_s(FullAdder_2247_io_s),
    .io_co(FullAdder_2247_io_co)
  );
  FullAdder FullAdder_2248 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2248_io_a),
    .io_b(FullAdder_2248_io_b),
    .io_ci(FullAdder_2248_io_ci),
    .io_s(FullAdder_2248_io_s),
    .io_co(FullAdder_2248_io_co)
  );
  FullAdder FullAdder_2249 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2249_io_a),
    .io_b(FullAdder_2249_io_b),
    .io_ci(FullAdder_2249_io_ci),
    .io_s(FullAdder_2249_io_s),
    .io_co(FullAdder_2249_io_co)
  );
  FullAdder FullAdder_2250 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2250_io_a),
    .io_b(FullAdder_2250_io_b),
    .io_ci(FullAdder_2250_io_ci),
    .io_s(FullAdder_2250_io_s),
    .io_co(FullAdder_2250_io_co)
  );
  FullAdder FullAdder_2251 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2251_io_a),
    .io_b(FullAdder_2251_io_b),
    .io_ci(FullAdder_2251_io_ci),
    .io_s(FullAdder_2251_io_s),
    .io_co(FullAdder_2251_io_co)
  );
  FullAdder FullAdder_2252 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2252_io_a),
    .io_b(FullAdder_2252_io_b),
    .io_ci(FullAdder_2252_io_ci),
    .io_s(FullAdder_2252_io_s),
    .io_co(FullAdder_2252_io_co)
  );
  FullAdder FullAdder_2253 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2253_io_a),
    .io_b(FullAdder_2253_io_b),
    .io_ci(FullAdder_2253_io_ci),
    .io_s(FullAdder_2253_io_s),
    .io_co(FullAdder_2253_io_co)
  );
  FullAdder FullAdder_2254 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2254_io_a),
    .io_b(FullAdder_2254_io_b),
    .io_ci(FullAdder_2254_io_ci),
    .io_s(FullAdder_2254_io_s),
    .io_co(FullAdder_2254_io_co)
  );
  FullAdder FullAdder_2255 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2255_io_a),
    .io_b(FullAdder_2255_io_b),
    .io_ci(FullAdder_2255_io_ci),
    .io_s(FullAdder_2255_io_s),
    .io_co(FullAdder_2255_io_co)
  );
  FullAdder FullAdder_2256 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2256_io_a),
    .io_b(FullAdder_2256_io_b),
    .io_ci(FullAdder_2256_io_ci),
    .io_s(FullAdder_2256_io_s),
    .io_co(FullAdder_2256_io_co)
  );
  FullAdder FullAdder_2257 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2257_io_a),
    .io_b(FullAdder_2257_io_b),
    .io_ci(FullAdder_2257_io_ci),
    .io_s(FullAdder_2257_io_s),
    .io_co(FullAdder_2257_io_co)
  );
  FullAdder FullAdder_2258 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2258_io_a),
    .io_b(FullAdder_2258_io_b),
    .io_ci(FullAdder_2258_io_ci),
    .io_s(FullAdder_2258_io_s),
    .io_co(FullAdder_2258_io_co)
  );
  FullAdder FullAdder_2259 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2259_io_a),
    .io_b(FullAdder_2259_io_b),
    .io_ci(FullAdder_2259_io_ci),
    .io_s(FullAdder_2259_io_s),
    .io_co(FullAdder_2259_io_co)
  );
  FullAdder FullAdder_2260 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2260_io_a),
    .io_b(FullAdder_2260_io_b),
    .io_ci(FullAdder_2260_io_ci),
    .io_s(FullAdder_2260_io_s),
    .io_co(FullAdder_2260_io_co)
  );
  FullAdder FullAdder_2261 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2261_io_a),
    .io_b(FullAdder_2261_io_b),
    .io_ci(FullAdder_2261_io_ci),
    .io_s(FullAdder_2261_io_s),
    .io_co(FullAdder_2261_io_co)
  );
  FullAdder FullAdder_2262 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2262_io_a),
    .io_b(FullAdder_2262_io_b),
    .io_ci(FullAdder_2262_io_ci),
    .io_s(FullAdder_2262_io_s),
    .io_co(FullAdder_2262_io_co)
  );
  FullAdder FullAdder_2263 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2263_io_a),
    .io_b(FullAdder_2263_io_b),
    .io_ci(FullAdder_2263_io_ci),
    .io_s(FullAdder_2263_io_s),
    .io_co(FullAdder_2263_io_co)
  );
  FullAdder FullAdder_2264 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2264_io_a),
    .io_b(FullAdder_2264_io_b),
    .io_ci(FullAdder_2264_io_ci),
    .io_s(FullAdder_2264_io_s),
    .io_co(FullAdder_2264_io_co)
  );
  FullAdder FullAdder_2265 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2265_io_a),
    .io_b(FullAdder_2265_io_b),
    .io_ci(FullAdder_2265_io_ci),
    .io_s(FullAdder_2265_io_s),
    .io_co(FullAdder_2265_io_co)
  );
  FullAdder FullAdder_2266 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2266_io_a),
    .io_b(FullAdder_2266_io_b),
    .io_ci(FullAdder_2266_io_ci),
    .io_s(FullAdder_2266_io_s),
    .io_co(FullAdder_2266_io_co)
  );
  FullAdder FullAdder_2267 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2267_io_a),
    .io_b(FullAdder_2267_io_b),
    .io_ci(FullAdder_2267_io_ci),
    .io_s(FullAdder_2267_io_s),
    .io_co(FullAdder_2267_io_co)
  );
  FullAdder FullAdder_2268 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2268_io_a),
    .io_b(FullAdder_2268_io_b),
    .io_ci(FullAdder_2268_io_ci),
    .io_s(FullAdder_2268_io_s),
    .io_co(FullAdder_2268_io_co)
  );
  FullAdder FullAdder_2269 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2269_io_a),
    .io_b(FullAdder_2269_io_b),
    .io_ci(FullAdder_2269_io_ci),
    .io_s(FullAdder_2269_io_s),
    .io_co(FullAdder_2269_io_co)
  );
  FullAdder FullAdder_2270 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2270_io_a),
    .io_b(FullAdder_2270_io_b),
    .io_ci(FullAdder_2270_io_ci),
    .io_s(FullAdder_2270_io_s),
    .io_co(FullAdder_2270_io_co)
  );
  FullAdder FullAdder_2271 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2271_io_a),
    .io_b(FullAdder_2271_io_b),
    .io_ci(FullAdder_2271_io_ci),
    .io_s(FullAdder_2271_io_s),
    .io_co(FullAdder_2271_io_co)
  );
  FullAdder FullAdder_2272 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2272_io_a),
    .io_b(FullAdder_2272_io_b),
    .io_ci(FullAdder_2272_io_ci),
    .io_s(FullAdder_2272_io_s),
    .io_co(FullAdder_2272_io_co)
  );
  FullAdder FullAdder_2273 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2273_io_a),
    .io_b(FullAdder_2273_io_b),
    .io_ci(FullAdder_2273_io_ci),
    .io_s(FullAdder_2273_io_s),
    .io_co(FullAdder_2273_io_co)
  );
  FullAdder FullAdder_2274 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2274_io_a),
    .io_b(FullAdder_2274_io_b),
    .io_ci(FullAdder_2274_io_ci),
    .io_s(FullAdder_2274_io_s),
    .io_co(FullAdder_2274_io_co)
  );
  FullAdder FullAdder_2275 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2275_io_a),
    .io_b(FullAdder_2275_io_b),
    .io_ci(FullAdder_2275_io_ci),
    .io_s(FullAdder_2275_io_s),
    .io_co(FullAdder_2275_io_co)
  );
  FullAdder FullAdder_2276 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2276_io_a),
    .io_b(FullAdder_2276_io_b),
    .io_ci(FullAdder_2276_io_ci),
    .io_s(FullAdder_2276_io_s),
    .io_co(FullAdder_2276_io_co)
  );
  FullAdder FullAdder_2277 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2277_io_a),
    .io_b(FullAdder_2277_io_b),
    .io_ci(FullAdder_2277_io_ci),
    .io_s(FullAdder_2277_io_s),
    .io_co(FullAdder_2277_io_co)
  );
  FullAdder FullAdder_2278 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2278_io_a),
    .io_b(FullAdder_2278_io_b),
    .io_ci(FullAdder_2278_io_ci),
    .io_s(FullAdder_2278_io_s),
    .io_co(FullAdder_2278_io_co)
  );
  FullAdder FullAdder_2279 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2279_io_a),
    .io_b(FullAdder_2279_io_b),
    .io_ci(FullAdder_2279_io_ci),
    .io_s(FullAdder_2279_io_s),
    .io_co(FullAdder_2279_io_co)
  );
  FullAdder FullAdder_2280 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2280_io_a),
    .io_b(FullAdder_2280_io_b),
    .io_ci(FullAdder_2280_io_ci),
    .io_s(FullAdder_2280_io_s),
    .io_co(FullAdder_2280_io_co)
  );
  FullAdder FullAdder_2281 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2281_io_a),
    .io_b(FullAdder_2281_io_b),
    .io_ci(FullAdder_2281_io_ci),
    .io_s(FullAdder_2281_io_s),
    .io_co(FullAdder_2281_io_co)
  );
  FullAdder FullAdder_2282 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2282_io_a),
    .io_b(FullAdder_2282_io_b),
    .io_ci(FullAdder_2282_io_ci),
    .io_s(FullAdder_2282_io_s),
    .io_co(FullAdder_2282_io_co)
  );
  FullAdder FullAdder_2283 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2283_io_a),
    .io_b(FullAdder_2283_io_b),
    .io_ci(FullAdder_2283_io_ci),
    .io_s(FullAdder_2283_io_s),
    .io_co(FullAdder_2283_io_co)
  );
  FullAdder FullAdder_2284 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2284_io_a),
    .io_b(FullAdder_2284_io_b),
    .io_ci(FullAdder_2284_io_ci),
    .io_s(FullAdder_2284_io_s),
    .io_co(FullAdder_2284_io_co)
  );
  FullAdder FullAdder_2285 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2285_io_a),
    .io_b(FullAdder_2285_io_b),
    .io_ci(FullAdder_2285_io_ci),
    .io_s(FullAdder_2285_io_s),
    .io_co(FullAdder_2285_io_co)
  );
  FullAdder FullAdder_2286 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2286_io_a),
    .io_b(FullAdder_2286_io_b),
    .io_ci(FullAdder_2286_io_ci),
    .io_s(FullAdder_2286_io_s),
    .io_co(FullAdder_2286_io_co)
  );
  FullAdder FullAdder_2287 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2287_io_a),
    .io_b(FullAdder_2287_io_b),
    .io_ci(FullAdder_2287_io_ci),
    .io_s(FullAdder_2287_io_s),
    .io_co(FullAdder_2287_io_co)
  );
  FullAdder FullAdder_2288 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2288_io_a),
    .io_b(FullAdder_2288_io_b),
    .io_ci(FullAdder_2288_io_ci),
    .io_s(FullAdder_2288_io_s),
    .io_co(FullAdder_2288_io_co)
  );
  FullAdder FullAdder_2289 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2289_io_a),
    .io_b(FullAdder_2289_io_b),
    .io_ci(FullAdder_2289_io_ci),
    .io_s(FullAdder_2289_io_s),
    .io_co(FullAdder_2289_io_co)
  );
  FullAdder FullAdder_2290 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2290_io_a),
    .io_b(FullAdder_2290_io_b),
    .io_ci(FullAdder_2290_io_ci),
    .io_s(FullAdder_2290_io_s),
    .io_co(FullAdder_2290_io_co)
  );
  FullAdder FullAdder_2291 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2291_io_a),
    .io_b(FullAdder_2291_io_b),
    .io_ci(FullAdder_2291_io_ci),
    .io_s(FullAdder_2291_io_s),
    .io_co(FullAdder_2291_io_co)
  );
  FullAdder FullAdder_2292 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2292_io_a),
    .io_b(FullAdder_2292_io_b),
    .io_ci(FullAdder_2292_io_ci),
    .io_s(FullAdder_2292_io_s),
    .io_co(FullAdder_2292_io_co)
  );
  FullAdder FullAdder_2293 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2293_io_a),
    .io_b(FullAdder_2293_io_b),
    .io_ci(FullAdder_2293_io_ci),
    .io_s(FullAdder_2293_io_s),
    .io_co(FullAdder_2293_io_co)
  );
  FullAdder FullAdder_2294 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2294_io_a),
    .io_b(FullAdder_2294_io_b),
    .io_ci(FullAdder_2294_io_ci),
    .io_s(FullAdder_2294_io_s),
    .io_co(FullAdder_2294_io_co)
  );
  FullAdder FullAdder_2295 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2295_io_a),
    .io_b(FullAdder_2295_io_b),
    .io_ci(FullAdder_2295_io_ci),
    .io_s(FullAdder_2295_io_s),
    .io_co(FullAdder_2295_io_co)
  );
  FullAdder FullAdder_2296 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2296_io_a),
    .io_b(FullAdder_2296_io_b),
    .io_ci(FullAdder_2296_io_ci),
    .io_s(FullAdder_2296_io_s),
    .io_co(FullAdder_2296_io_co)
  );
  FullAdder FullAdder_2297 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2297_io_a),
    .io_b(FullAdder_2297_io_b),
    .io_ci(FullAdder_2297_io_ci),
    .io_s(FullAdder_2297_io_s),
    .io_co(FullAdder_2297_io_co)
  );
  FullAdder FullAdder_2298 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2298_io_a),
    .io_b(FullAdder_2298_io_b),
    .io_ci(FullAdder_2298_io_ci),
    .io_s(FullAdder_2298_io_s),
    .io_co(FullAdder_2298_io_co)
  );
  FullAdder FullAdder_2299 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2299_io_a),
    .io_b(FullAdder_2299_io_b),
    .io_ci(FullAdder_2299_io_ci),
    .io_s(FullAdder_2299_io_s),
    .io_co(FullAdder_2299_io_co)
  );
  FullAdder FullAdder_2300 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2300_io_a),
    .io_b(FullAdder_2300_io_b),
    .io_ci(FullAdder_2300_io_ci),
    .io_s(FullAdder_2300_io_s),
    .io_co(FullAdder_2300_io_co)
  );
  FullAdder FullAdder_2301 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2301_io_a),
    .io_b(FullAdder_2301_io_b),
    .io_ci(FullAdder_2301_io_ci),
    .io_s(FullAdder_2301_io_s),
    .io_co(FullAdder_2301_io_co)
  );
  FullAdder FullAdder_2302 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2302_io_a),
    .io_b(FullAdder_2302_io_b),
    .io_ci(FullAdder_2302_io_ci),
    .io_s(FullAdder_2302_io_s),
    .io_co(FullAdder_2302_io_co)
  );
  FullAdder FullAdder_2303 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2303_io_a),
    .io_b(FullAdder_2303_io_b),
    .io_ci(FullAdder_2303_io_ci),
    .io_s(FullAdder_2303_io_s),
    .io_co(FullAdder_2303_io_co)
  );
  FullAdder FullAdder_2304 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2304_io_a),
    .io_b(FullAdder_2304_io_b),
    .io_ci(FullAdder_2304_io_ci),
    .io_s(FullAdder_2304_io_s),
    .io_co(FullAdder_2304_io_co)
  );
  FullAdder FullAdder_2305 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2305_io_a),
    .io_b(FullAdder_2305_io_b),
    .io_ci(FullAdder_2305_io_ci),
    .io_s(FullAdder_2305_io_s),
    .io_co(FullAdder_2305_io_co)
  );
  FullAdder FullAdder_2306 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2306_io_a),
    .io_b(FullAdder_2306_io_b),
    .io_ci(FullAdder_2306_io_ci),
    .io_s(FullAdder_2306_io_s),
    .io_co(FullAdder_2306_io_co)
  );
  FullAdder FullAdder_2307 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2307_io_a),
    .io_b(FullAdder_2307_io_b),
    .io_ci(FullAdder_2307_io_ci),
    .io_s(FullAdder_2307_io_s),
    .io_co(FullAdder_2307_io_co)
  );
  FullAdder FullAdder_2308 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2308_io_a),
    .io_b(FullAdder_2308_io_b),
    .io_ci(FullAdder_2308_io_ci),
    .io_s(FullAdder_2308_io_s),
    .io_co(FullAdder_2308_io_co)
  );
  FullAdder FullAdder_2309 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2309_io_a),
    .io_b(FullAdder_2309_io_b),
    .io_ci(FullAdder_2309_io_ci),
    .io_s(FullAdder_2309_io_s),
    .io_co(FullAdder_2309_io_co)
  );
  FullAdder FullAdder_2310 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2310_io_a),
    .io_b(FullAdder_2310_io_b),
    .io_ci(FullAdder_2310_io_ci),
    .io_s(FullAdder_2310_io_s),
    .io_co(FullAdder_2310_io_co)
  );
  FullAdder FullAdder_2311 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2311_io_a),
    .io_b(FullAdder_2311_io_b),
    .io_ci(FullAdder_2311_io_ci),
    .io_s(FullAdder_2311_io_s),
    .io_co(FullAdder_2311_io_co)
  );
  FullAdder FullAdder_2312 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2312_io_a),
    .io_b(FullAdder_2312_io_b),
    .io_ci(FullAdder_2312_io_ci),
    .io_s(FullAdder_2312_io_s),
    .io_co(FullAdder_2312_io_co)
  );
  FullAdder FullAdder_2313 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2313_io_a),
    .io_b(FullAdder_2313_io_b),
    .io_ci(FullAdder_2313_io_ci),
    .io_s(FullAdder_2313_io_s),
    .io_co(FullAdder_2313_io_co)
  );
  FullAdder FullAdder_2314 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2314_io_a),
    .io_b(FullAdder_2314_io_b),
    .io_ci(FullAdder_2314_io_ci),
    .io_s(FullAdder_2314_io_s),
    .io_co(FullAdder_2314_io_co)
  );
  FullAdder FullAdder_2315 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2315_io_a),
    .io_b(FullAdder_2315_io_b),
    .io_ci(FullAdder_2315_io_ci),
    .io_s(FullAdder_2315_io_s),
    .io_co(FullAdder_2315_io_co)
  );
  FullAdder FullAdder_2316 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2316_io_a),
    .io_b(FullAdder_2316_io_b),
    .io_ci(FullAdder_2316_io_ci),
    .io_s(FullAdder_2316_io_s),
    .io_co(FullAdder_2316_io_co)
  );
  FullAdder FullAdder_2317 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2317_io_a),
    .io_b(FullAdder_2317_io_b),
    .io_ci(FullAdder_2317_io_ci),
    .io_s(FullAdder_2317_io_s),
    .io_co(FullAdder_2317_io_co)
  );
  FullAdder FullAdder_2318 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2318_io_a),
    .io_b(FullAdder_2318_io_b),
    .io_ci(FullAdder_2318_io_ci),
    .io_s(FullAdder_2318_io_s),
    .io_co(FullAdder_2318_io_co)
  );
  FullAdder FullAdder_2319 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2319_io_a),
    .io_b(FullAdder_2319_io_b),
    .io_ci(FullAdder_2319_io_ci),
    .io_s(FullAdder_2319_io_s),
    .io_co(FullAdder_2319_io_co)
  );
  FullAdder FullAdder_2320 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2320_io_a),
    .io_b(FullAdder_2320_io_b),
    .io_ci(FullAdder_2320_io_ci),
    .io_s(FullAdder_2320_io_s),
    .io_co(FullAdder_2320_io_co)
  );
  FullAdder FullAdder_2321 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2321_io_a),
    .io_b(FullAdder_2321_io_b),
    .io_ci(FullAdder_2321_io_ci),
    .io_s(FullAdder_2321_io_s),
    .io_co(FullAdder_2321_io_co)
  );
  FullAdder FullAdder_2322 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2322_io_a),
    .io_b(FullAdder_2322_io_b),
    .io_ci(FullAdder_2322_io_ci),
    .io_s(FullAdder_2322_io_s),
    .io_co(FullAdder_2322_io_co)
  );
  FullAdder FullAdder_2323 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2323_io_a),
    .io_b(FullAdder_2323_io_b),
    .io_ci(FullAdder_2323_io_ci),
    .io_s(FullAdder_2323_io_s),
    .io_co(FullAdder_2323_io_co)
  );
  FullAdder FullAdder_2324 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2324_io_a),
    .io_b(FullAdder_2324_io_b),
    .io_ci(FullAdder_2324_io_ci),
    .io_s(FullAdder_2324_io_s),
    .io_co(FullAdder_2324_io_co)
  );
  FullAdder FullAdder_2325 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2325_io_a),
    .io_b(FullAdder_2325_io_b),
    .io_ci(FullAdder_2325_io_ci),
    .io_s(FullAdder_2325_io_s),
    .io_co(FullAdder_2325_io_co)
  );
  FullAdder FullAdder_2326 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2326_io_a),
    .io_b(FullAdder_2326_io_b),
    .io_ci(FullAdder_2326_io_ci),
    .io_s(FullAdder_2326_io_s),
    .io_co(FullAdder_2326_io_co)
  );
  FullAdder FullAdder_2327 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2327_io_a),
    .io_b(FullAdder_2327_io_b),
    .io_ci(FullAdder_2327_io_ci),
    .io_s(FullAdder_2327_io_s),
    .io_co(FullAdder_2327_io_co)
  );
  FullAdder FullAdder_2328 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2328_io_a),
    .io_b(FullAdder_2328_io_b),
    .io_ci(FullAdder_2328_io_ci),
    .io_s(FullAdder_2328_io_s),
    .io_co(FullAdder_2328_io_co)
  );
  FullAdder FullAdder_2329 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2329_io_a),
    .io_b(FullAdder_2329_io_b),
    .io_ci(FullAdder_2329_io_ci),
    .io_s(FullAdder_2329_io_s),
    .io_co(FullAdder_2329_io_co)
  );
  FullAdder FullAdder_2330 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2330_io_a),
    .io_b(FullAdder_2330_io_b),
    .io_ci(FullAdder_2330_io_ci),
    .io_s(FullAdder_2330_io_s),
    .io_co(FullAdder_2330_io_co)
  );
  FullAdder FullAdder_2331 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2331_io_a),
    .io_b(FullAdder_2331_io_b),
    .io_ci(FullAdder_2331_io_ci),
    .io_s(FullAdder_2331_io_s),
    .io_co(FullAdder_2331_io_co)
  );
  FullAdder FullAdder_2332 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2332_io_a),
    .io_b(FullAdder_2332_io_b),
    .io_ci(FullAdder_2332_io_ci),
    .io_s(FullAdder_2332_io_s),
    .io_co(FullAdder_2332_io_co)
  );
  FullAdder FullAdder_2333 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2333_io_a),
    .io_b(FullAdder_2333_io_b),
    .io_ci(FullAdder_2333_io_ci),
    .io_s(FullAdder_2333_io_s),
    .io_co(FullAdder_2333_io_co)
  );
  FullAdder FullAdder_2334 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2334_io_a),
    .io_b(FullAdder_2334_io_b),
    .io_ci(FullAdder_2334_io_ci),
    .io_s(FullAdder_2334_io_s),
    .io_co(FullAdder_2334_io_co)
  );
  FullAdder FullAdder_2335 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2335_io_a),
    .io_b(FullAdder_2335_io_b),
    .io_ci(FullAdder_2335_io_ci),
    .io_s(FullAdder_2335_io_s),
    .io_co(FullAdder_2335_io_co)
  );
  FullAdder FullAdder_2336 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2336_io_a),
    .io_b(FullAdder_2336_io_b),
    .io_ci(FullAdder_2336_io_ci),
    .io_s(FullAdder_2336_io_s),
    .io_co(FullAdder_2336_io_co)
  );
  FullAdder FullAdder_2337 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2337_io_a),
    .io_b(FullAdder_2337_io_b),
    .io_ci(FullAdder_2337_io_ci),
    .io_s(FullAdder_2337_io_s),
    .io_co(FullAdder_2337_io_co)
  );
  FullAdder FullAdder_2338 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2338_io_a),
    .io_b(FullAdder_2338_io_b),
    .io_ci(FullAdder_2338_io_ci),
    .io_s(FullAdder_2338_io_s),
    .io_co(FullAdder_2338_io_co)
  );
  HalfAdder HalfAdder_75 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_75_io_a),
    .io_b(HalfAdder_75_io_b),
    .io_s(HalfAdder_75_io_s),
    .io_co(HalfAdder_75_io_co)
  );
  FullAdder FullAdder_2339 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2339_io_a),
    .io_b(FullAdder_2339_io_b),
    .io_ci(FullAdder_2339_io_ci),
    .io_s(FullAdder_2339_io_s),
    .io_co(FullAdder_2339_io_co)
  );
  FullAdder FullAdder_2340 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2340_io_a),
    .io_b(FullAdder_2340_io_b),
    .io_ci(FullAdder_2340_io_ci),
    .io_s(FullAdder_2340_io_s),
    .io_co(FullAdder_2340_io_co)
  );
  FullAdder FullAdder_2341 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2341_io_a),
    .io_b(FullAdder_2341_io_b),
    .io_ci(FullAdder_2341_io_ci),
    .io_s(FullAdder_2341_io_s),
    .io_co(FullAdder_2341_io_co)
  );
  FullAdder FullAdder_2342 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2342_io_a),
    .io_b(FullAdder_2342_io_b),
    .io_ci(FullAdder_2342_io_ci),
    .io_s(FullAdder_2342_io_s),
    .io_co(FullAdder_2342_io_co)
  );
  FullAdder FullAdder_2343 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2343_io_a),
    .io_b(FullAdder_2343_io_b),
    .io_ci(FullAdder_2343_io_ci),
    .io_s(FullAdder_2343_io_s),
    .io_co(FullAdder_2343_io_co)
  );
  FullAdder FullAdder_2344 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2344_io_a),
    .io_b(FullAdder_2344_io_b),
    .io_ci(FullAdder_2344_io_ci),
    .io_s(FullAdder_2344_io_s),
    .io_co(FullAdder_2344_io_co)
  );
  HalfAdder HalfAdder_76 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_76_io_a),
    .io_b(HalfAdder_76_io_b),
    .io_s(HalfAdder_76_io_s),
    .io_co(HalfAdder_76_io_co)
  );
  FullAdder FullAdder_2345 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2345_io_a),
    .io_b(FullAdder_2345_io_b),
    .io_ci(FullAdder_2345_io_ci),
    .io_s(FullAdder_2345_io_s),
    .io_co(FullAdder_2345_io_co)
  );
  FullAdder FullAdder_2346 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2346_io_a),
    .io_b(FullAdder_2346_io_b),
    .io_ci(FullAdder_2346_io_ci),
    .io_s(FullAdder_2346_io_s),
    .io_co(FullAdder_2346_io_co)
  );
  FullAdder FullAdder_2347 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2347_io_a),
    .io_b(FullAdder_2347_io_b),
    .io_ci(FullAdder_2347_io_ci),
    .io_s(FullAdder_2347_io_s),
    .io_co(FullAdder_2347_io_co)
  );
  FullAdder FullAdder_2348 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2348_io_a),
    .io_b(FullAdder_2348_io_b),
    .io_ci(FullAdder_2348_io_ci),
    .io_s(FullAdder_2348_io_s),
    .io_co(FullAdder_2348_io_co)
  );
  FullAdder FullAdder_2349 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2349_io_a),
    .io_b(FullAdder_2349_io_b),
    .io_ci(FullAdder_2349_io_ci),
    .io_s(FullAdder_2349_io_s),
    .io_co(FullAdder_2349_io_co)
  );
  FullAdder FullAdder_2350 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2350_io_a),
    .io_b(FullAdder_2350_io_b),
    .io_ci(FullAdder_2350_io_ci),
    .io_s(FullAdder_2350_io_s),
    .io_co(FullAdder_2350_io_co)
  );
  FullAdder FullAdder_2351 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2351_io_a),
    .io_b(FullAdder_2351_io_b),
    .io_ci(FullAdder_2351_io_ci),
    .io_s(FullAdder_2351_io_s),
    .io_co(FullAdder_2351_io_co)
  );
  FullAdder FullAdder_2352 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2352_io_a),
    .io_b(FullAdder_2352_io_b),
    .io_ci(FullAdder_2352_io_ci),
    .io_s(FullAdder_2352_io_s),
    .io_co(FullAdder_2352_io_co)
  );
  FullAdder FullAdder_2353 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2353_io_a),
    .io_b(FullAdder_2353_io_b),
    .io_ci(FullAdder_2353_io_ci),
    .io_s(FullAdder_2353_io_s),
    .io_co(FullAdder_2353_io_co)
  );
  FullAdder FullAdder_2354 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2354_io_a),
    .io_b(FullAdder_2354_io_b),
    .io_ci(FullAdder_2354_io_ci),
    .io_s(FullAdder_2354_io_s),
    .io_co(FullAdder_2354_io_co)
  );
  FullAdder FullAdder_2355 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2355_io_a),
    .io_b(FullAdder_2355_io_b),
    .io_ci(FullAdder_2355_io_ci),
    .io_s(FullAdder_2355_io_s),
    .io_co(FullAdder_2355_io_co)
  );
  FullAdder FullAdder_2356 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2356_io_a),
    .io_b(FullAdder_2356_io_b),
    .io_ci(FullAdder_2356_io_ci),
    .io_s(FullAdder_2356_io_s),
    .io_co(FullAdder_2356_io_co)
  );
  FullAdder FullAdder_2357 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2357_io_a),
    .io_b(FullAdder_2357_io_b),
    .io_ci(FullAdder_2357_io_ci),
    .io_s(FullAdder_2357_io_s),
    .io_co(FullAdder_2357_io_co)
  );
  FullAdder FullAdder_2358 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2358_io_a),
    .io_b(FullAdder_2358_io_b),
    .io_ci(FullAdder_2358_io_ci),
    .io_s(FullAdder_2358_io_s),
    .io_co(FullAdder_2358_io_co)
  );
  FullAdder FullAdder_2359 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2359_io_a),
    .io_b(FullAdder_2359_io_b),
    .io_ci(FullAdder_2359_io_ci),
    .io_s(FullAdder_2359_io_s),
    .io_co(FullAdder_2359_io_co)
  );
  FullAdder FullAdder_2360 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2360_io_a),
    .io_b(FullAdder_2360_io_b),
    .io_ci(FullAdder_2360_io_ci),
    .io_s(FullAdder_2360_io_s),
    .io_co(FullAdder_2360_io_co)
  );
  FullAdder FullAdder_2361 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2361_io_a),
    .io_b(FullAdder_2361_io_b),
    .io_ci(FullAdder_2361_io_ci),
    .io_s(FullAdder_2361_io_s),
    .io_co(FullAdder_2361_io_co)
  );
  FullAdder FullAdder_2362 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2362_io_a),
    .io_b(FullAdder_2362_io_b),
    .io_ci(FullAdder_2362_io_ci),
    .io_s(FullAdder_2362_io_s),
    .io_co(FullAdder_2362_io_co)
  );
  FullAdder FullAdder_2363 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2363_io_a),
    .io_b(FullAdder_2363_io_b),
    .io_ci(FullAdder_2363_io_ci),
    .io_s(FullAdder_2363_io_s),
    .io_co(FullAdder_2363_io_co)
  );
  FullAdder FullAdder_2364 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2364_io_a),
    .io_b(FullAdder_2364_io_b),
    .io_ci(FullAdder_2364_io_ci),
    .io_s(FullAdder_2364_io_s),
    .io_co(FullAdder_2364_io_co)
  );
  FullAdder FullAdder_2365 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2365_io_a),
    .io_b(FullAdder_2365_io_b),
    .io_ci(FullAdder_2365_io_ci),
    .io_s(FullAdder_2365_io_s),
    .io_co(FullAdder_2365_io_co)
  );
  FullAdder FullAdder_2366 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2366_io_a),
    .io_b(FullAdder_2366_io_b),
    .io_ci(FullAdder_2366_io_ci),
    .io_s(FullAdder_2366_io_s),
    .io_co(FullAdder_2366_io_co)
  );
  FullAdder FullAdder_2367 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2367_io_a),
    .io_b(FullAdder_2367_io_b),
    .io_ci(FullAdder_2367_io_ci),
    .io_s(FullAdder_2367_io_s),
    .io_co(FullAdder_2367_io_co)
  );
  FullAdder FullAdder_2368 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2368_io_a),
    .io_b(FullAdder_2368_io_b),
    .io_ci(FullAdder_2368_io_ci),
    .io_s(FullAdder_2368_io_s),
    .io_co(FullAdder_2368_io_co)
  );
  FullAdder FullAdder_2369 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2369_io_a),
    .io_b(FullAdder_2369_io_b),
    .io_ci(FullAdder_2369_io_ci),
    .io_s(FullAdder_2369_io_s),
    .io_co(FullAdder_2369_io_co)
  );
  FullAdder FullAdder_2370 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2370_io_a),
    .io_b(FullAdder_2370_io_b),
    .io_ci(FullAdder_2370_io_ci),
    .io_s(FullAdder_2370_io_s),
    .io_co(FullAdder_2370_io_co)
  );
  FullAdder FullAdder_2371 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2371_io_a),
    .io_b(FullAdder_2371_io_b),
    .io_ci(FullAdder_2371_io_ci),
    .io_s(FullAdder_2371_io_s),
    .io_co(FullAdder_2371_io_co)
  );
  FullAdder FullAdder_2372 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2372_io_a),
    .io_b(FullAdder_2372_io_b),
    .io_ci(FullAdder_2372_io_ci),
    .io_s(FullAdder_2372_io_s),
    .io_co(FullAdder_2372_io_co)
  );
  FullAdder FullAdder_2373 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2373_io_a),
    .io_b(FullAdder_2373_io_b),
    .io_ci(FullAdder_2373_io_ci),
    .io_s(FullAdder_2373_io_s),
    .io_co(FullAdder_2373_io_co)
  );
  FullAdder FullAdder_2374 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2374_io_a),
    .io_b(FullAdder_2374_io_b),
    .io_ci(FullAdder_2374_io_ci),
    .io_s(FullAdder_2374_io_s),
    .io_co(FullAdder_2374_io_co)
  );
  FullAdder FullAdder_2375 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2375_io_a),
    .io_b(FullAdder_2375_io_b),
    .io_ci(FullAdder_2375_io_ci),
    .io_s(FullAdder_2375_io_s),
    .io_co(FullAdder_2375_io_co)
  );
  FullAdder FullAdder_2376 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2376_io_a),
    .io_b(FullAdder_2376_io_b),
    .io_ci(FullAdder_2376_io_ci),
    .io_s(FullAdder_2376_io_s),
    .io_co(FullAdder_2376_io_co)
  );
  FullAdder FullAdder_2377 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2377_io_a),
    .io_b(FullAdder_2377_io_b),
    .io_ci(FullAdder_2377_io_ci),
    .io_s(FullAdder_2377_io_s),
    .io_co(FullAdder_2377_io_co)
  );
  FullAdder FullAdder_2378 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2378_io_a),
    .io_b(FullAdder_2378_io_b),
    .io_ci(FullAdder_2378_io_ci),
    .io_s(FullAdder_2378_io_s),
    .io_co(FullAdder_2378_io_co)
  );
  FullAdder FullAdder_2379 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2379_io_a),
    .io_b(FullAdder_2379_io_b),
    .io_ci(FullAdder_2379_io_ci),
    .io_s(FullAdder_2379_io_s),
    .io_co(FullAdder_2379_io_co)
  );
  FullAdder FullAdder_2380 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2380_io_a),
    .io_b(FullAdder_2380_io_b),
    .io_ci(FullAdder_2380_io_ci),
    .io_s(FullAdder_2380_io_s),
    .io_co(FullAdder_2380_io_co)
  );
  FullAdder FullAdder_2381 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2381_io_a),
    .io_b(FullAdder_2381_io_b),
    .io_ci(FullAdder_2381_io_ci),
    .io_s(FullAdder_2381_io_s),
    .io_co(FullAdder_2381_io_co)
  );
  FullAdder FullAdder_2382 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2382_io_a),
    .io_b(FullAdder_2382_io_b),
    .io_ci(FullAdder_2382_io_ci),
    .io_s(FullAdder_2382_io_s),
    .io_co(FullAdder_2382_io_co)
  );
  FullAdder FullAdder_2383 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2383_io_a),
    .io_b(FullAdder_2383_io_b),
    .io_ci(FullAdder_2383_io_ci),
    .io_s(FullAdder_2383_io_s),
    .io_co(FullAdder_2383_io_co)
  );
  FullAdder FullAdder_2384 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2384_io_a),
    .io_b(FullAdder_2384_io_b),
    .io_ci(FullAdder_2384_io_ci),
    .io_s(FullAdder_2384_io_s),
    .io_co(FullAdder_2384_io_co)
  );
  FullAdder FullAdder_2385 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2385_io_a),
    .io_b(FullAdder_2385_io_b),
    .io_ci(FullAdder_2385_io_ci),
    .io_s(FullAdder_2385_io_s),
    .io_co(FullAdder_2385_io_co)
  );
  HalfAdder HalfAdder_77 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_77_io_a),
    .io_b(HalfAdder_77_io_b),
    .io_s(HalfAdder_77_io_s),
    .io_co(HalfAdder_77_io_co)
  );
  FullAdder FullAdder_2386 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2386_io_a),
    .io_b(FullAdder_2386_io_b),
    .io_ci(FullAdder_2386_io_ci),
    .io_s(FullAdder_2386_io_s),
    .io_co(FullAdder_2386_io_co)
  );
  FullAdder FullAdder_2387 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2387_io_a),
    .io_b(FullAdder_2387_io_b),
    .io_ci(FullAdder_2387_io_ci),
    .io_s(FullAdder_2387_io_s),
    .io_co(FullAdder_2387_io_co)
  );
  FullAdder FullAdder_2388 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2388_io_a),
    .io_b(FullAdder_2388_io_b),
    .io_ci(FullAdder_2388_io_ci),
    .io_s(FullAdder_2388_io_s),
    .io_co(FullAdder_2388_io_co)
  );
  FullAdder FullAdder_2389 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2389_io_a),
    .io_b(FullAdder_2389_io_b),
    .io_ci(FullAdder_2389_io_ci),
    .io_s(FullAdder_2389_io_s),
    .io_co(FullAdder_2389_io_co)
  );
  FullAdder FullAdder_2390 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2390_io_a),
    .io_b(FullAdder_2390_io_b),
    .io_ci(FullAdder_2390_io_ci),
    .io_s(FullAdder_2390_io_s),
    .io_co(FullAdder_2390_io_co)
  );
  FullAdder FullAdder_2391 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2391_io_a),
    .io_b(FullAdder_2391_io_b),
    .io_ci(FullAdder_2391_io_ci),
    .io_s(FullAdder_2391_io_s),
    .io_co(FullAdder_2391_io_co)
  );
  FullAdder FullAdder_2392 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2392_io_a),
    .io_b(FullAdder_2392_io_b),
    .io_ci(FullAdder_2392_io_ci),
    .io_s(FullAdder_2392_io_s),
    .io_co(FullAdder_2392_io_co)
  );
  FullAdder FullAdder_2393 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2393_io_a),
    .io_b(FullAdder_2393_io_b),
    .io_ci(FullAdder_2393_io_ci),
    .io_s(FullAdder_2393_io_s),
    .io_co(FullAdder_2393_io_co)
  );
  FullAdder FullAdder_2394 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2394_io_a),
    .io_b(FullAdder_2394_io_b),
    .io_ci(FullAdder_2394_io_ci),
    .io_s(FullAdder_2394_io_s),
    .io_co(FullAdder_2394_io_co)
  );
  FullAdder FullAdder_2395 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2395_io_a),
    .io_b(FullAdder_2395_io_b),
    .io_ci(FullAdder_2395_io_ci),
    .io_s(FullAdder_2395_io_s),
    .io_co(FullAdder_2395_io_co)
  );
  FullAdder FullAdder_2396 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2396_io_a),
    .io_b(FullAdder_2396_io_b),
    .io_ci(FullAdder_2396_io_ci),
    .io_s(FullAdder_2396_io_s),
    .io_co(FullAdder_2396_io_co)
  );
  FullAdder FullAdder_2397 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2397_io_a),
    .io_b(FullAdder_2397_io_b),
    .io_ci(FullAdder_2397_io_ci),
    .io_s(FullAdder_2397_io_s),
    .io_co(FullAdder_2397_io_co)
  );
  FullAdder FullAdder_2398 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2398_io_a),
    .io_b(FullAdder_2398_io_b),
    .io_ci(FullAdder_2398_io_ci),
    .io_s(FullAdder_2398_io_s),
    .io_co(FullAdder_2398_io_co)
  );
  FullAdder FullAdder_2399 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2399_io_a),
    .io_b(FullAdder_2399_io_b),
    .io_ci(FullAdder_2399_io_ci),
    .io_s(FullAdder_2399_io_s),
    .io_co(FullAdder_2399_io_co)
  );
  FullAdder FullAdder_2400 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2400_io_a),
    .io_b(FullAdder_2400_io_b),
    .io_ci(FullAdder_2400_io_ci),
    .io_s(FullAdder_2400_io_s),
    .io_co(FullAdder_2400_io_co)
  );
  FullAdder FullAdder_2401 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2401_io_a),
    .io_b(FullAdder_2401_io_b),
    .io_ci(FullAdder_2401_io_ci),
    .io_s(FullAdder_2401_io_s),
    .io_co(FullAdder_2401_io_co)
  );
  FullAdder FullAdder_2402 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2402_io_a),
    .io_b(FullAdder_2402_io_b),
    .io_ci(FullAdder_2402_io_ci),
    .io_s(FullAdder_2402_io_s),
    .io_co(FullAdder_2402_io_co)
  );
  FullAdder FullAdder_2403 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2403_io_a),
    .io_b(FullAdder_2403_io_b),
    .io_ci(FullAdder_2403_io_ci),
    .io_s(FullAdder_2403_io_s),
    .io_co(FullAdder_2403_io_co)
  );
  FullAdder FullAdder_2404 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2404_io_a),
    .io_b(FullAdder_2404_io_b),
    .io_ci(FullAdder_2404_io_ci),
    .io_s(FullAdder_2404_io_s),
    .io_co(FullAdder_2404_io_co)
  );
  FullAdder FullAdder_2405 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2405_io_a),
    .io_b(FullAdder_2405_io_b),
    .io_ci(FullAdder_2405_io_ci),
    .io_s(FullAdder_2405_io_s),
    .io_co(FullAdder_2405_io_co)
  );
  FullAdder FullAdder_2406 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2406_io_a),
    .io_b(FullAdder_2406_io_b),
    .io_ci(FullAdder_2406_io_ci),
    .io_s(FullAdder_2406_io_s),
    .io_co(FullAdder_2406_io_co)
  );
  FullAdder FullAdder_2407 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2407_io_a),
    .io_b(FullAdder_2407_io_b),
    .io_ci(FullAdder_2407_io_ci),
    .io_s(FullAdder_2407_io_s),
    .io_co(FullAdder_2407_io_co)
  );
  FullAdder FullAdder_2408 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2408_io_a),
    .io_b(FullAdder_2408_io_b),
    .io_ci(FullAdder_2408_io_ci),
    .io_s(FullAdder_2408_io_s),
    .io_co(FullAdder_2408_io_co)
  );
  FullAdder FullAdder_2409 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2409_io_a),
    .io_b(FullAdder_2409_io_b),
    .io_ci(FullAdder_2409_io_ci),
    .io_s(FullAdder_2409_io_s),
    .io_co(FullAdder_2409_io_co)
  );
  FullAdder FullAdder_2410 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2410_io_a),
    .io_b(FullAdder_2410_io_b),
    .io_ci(FullAdder_2410_io_ci),
    .io_s(FullAdder_2410_io_s),
    .io_co(FullAdder_2410_io_co)
  );
  FullAdder FullAdder_2411 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2411_io_a),
    .io_b(FullAdder_2411_io_b),
    .io_ci(FullAdder_2411_io_ci),
    .io_s(FullAdder_2411_io_s),
    .io_co(FullAdder_2411_io_co)
  );
  FullAdder FullAdder_2412 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2412_io_a),
    .io_b(FullAdder_2412_io_b),
    .io_ci(FullAdder_2412_io_ci),
    .io_s(FullAdder_2412_io_s),
    .io_co(FullAdder_2412_io_co)
  );
  FullAdder FullAdder_2413 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2413_io_a),
    .io_b(FullAdder_2413_io_b),
    .io_ci(FullAdder_2413_io_ci),
    .io_s(FullAdder_2413_io_s),
    .io_co(FullAdder_2413_io_co)
  );
  FullAdder FullAdder_2414 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2414_io_a),
    .io_b(FullAdder_2414_io_b),
    .io_ci(FullAdder_2414_io_ci),
    .io_s(FullAdder_2414_io_s),
    .io_co(FullAdder_2414_io_co)
  );
  FullAdder FullAdder_2415 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2415_io_a),
    .io_b(FullAdder_2415_io_b),
    .io_ci(FullAdder_2415_io_ci),
    .io_s(FullAdder_2415_io_s),
    .io_co(FullAdder_2415_io_co)
  );
  FullAdder FullAdder_2416 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2416_io_a),
    .io_b(FullAdder_2416_io_b),
    .io_ci(FullAdder_2416_io_ci),
    .io_s(FullAdder_2416_io_s),
    .io_co(FullAdder_2416_io_co)
  );
  FullAdder FullAdder_2417 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2417_io_a),
    .io_b(FullAdder_2417_io_b),
    .io_ci(FullAdder_2417_io_ci),
    .io_s(FullAdder_2417_io_s),
    .io_co(FullAdder_2417_io_co)
  );
  FullAdder FullAdder_2418 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2418_io_a),
    .io_b(FullAdder_2418_io_b),
    .io_ci(FullAdder_2418_io_ci),
    .io_s(FullAdder_2418_io_s),
    .io_co(FullAdder_2418_io_co)
  );
  FullAdder FullAdder_2419 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2419_io_a),
    .io_b(FullAdder_2419_io_b),
    .io_ci(FullAdder_2419_io_ci),
    .io_s(FullAdder_2419_io_s),
    .io_co(FullAdder_2419_io_co)
  );
  FullAdder FullAdder_2420 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2420_io_a),
    .io_b(FullAdder_2420_io_b),
    .io_ci(FullAdder_2420_io_ci),
    .io_s(FullAdder_2420_io_s),
    .io_co(FullAdder_2420_io_co)
  );
  FullAdder FullAdder_2421 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2421_io_a),
    .io_b(FullAdder_2421_io_b),
    .io_ci(FullAdder_2421_io_ci),
    .io_s(FullAdder_2421_io_s),
    .io_co(FullAdder_2421_io_co)
  );
  FullAdder FullAdder_2422 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2422_io_a),
    .io_b(FullAdder_2422_io_b),
    .io_ci(FullAdder_2422_io_ci),
    .io_s(FullAdder_2422_io_s),
    .io_co(FullAdder_2422_io_co)
  );
  FullAdder FullAdder_2423 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2423_io_a),
    .io_b(FullAdder_2423_io_b),
    .io_ci(FullAdder_2423_io_ci),
    .io_s(FullAdder_2423_io_s),
    .io_co(FullAdder_2423_io_co)
  );
  FullAdder FullAdder_2424 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2424_io_a),
    .io_b(FullAdder_2424_io_b),
    .io_ci(FullAdder_2424_io_ci),
    .io_s(FullAdder_2424_io_s),
    .io_co(FullAdder_2424_io_co)
  );
  FullAdder FullAdder_2425 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2425_io_a),
    .io_b(FullAdder_2425_io_b),
    .io_ci(FullAdder_2425_io_ci),
    .io_s(FullAdder_2425_io_s),
    .io_co(FullAdder_2425_io_co)
  );
  FullAdder FullAdder_2426 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2426_io_a),
    .io_b(FullAdder_2426_io_b),
    .io_ci(FullAdder_2426_io_ci),
    .io_s(FullAdder_2426_io_s),
    .io_co(FullAdder_2426_io_co)
  );
  FullAdder FullAdder_2427 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2427_io_a),
    .io_b(FullAdder_2427_io_b),
    .io_ci(FullAdder_2427_io_ci),
    .io_s(FullAdder_2427_io_s),
    .io_co(FullAdder_2427_io_co)
  );
  FullAdder FullAdder_2428 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2428_io_a),
    .io_b(FullAdder_2428_io_b),
    .io_ci(FullAdder_2428_io_ci),
    .io_s(FullAdder_2428_io_s),
    .io_co(FullAdder_2428_io_co)
  );
  FullAdder FullAdder_2429 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2429_io_a),
    .io_b(FullAdder_2429_io_b),
    .io_ci(FullAdder_2429_io_ci),
    .io_s(FullAdder_2429_io_s),
    .io_co(FullAdder_2429_io_co)
  );
  FullAdder FullAdder_2430 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2430_io_a),
    .io_b(FullAdder_2430_io_b),
    .io_ci(FullAdder_2430_io_ci),
    .io_s(FullAdder_2430_io_s),
    .io_co(FullAdder_2430_io_co)
  );
  FullAdder FullAdder_2431 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2431_io_a),
    .io_b(FullAdder_2431_io_b),
    .io_ci(FullAdder_2431_io_ci),
    .io_s(FullAdder_2431_io_s),
    .io_co(FullAdder_2431_io_co)
  );
  FullAdder FullAdder_2432 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2432_io_a),
    .io_b(FullAdder_2432_io_b),
    .io_ci(FullAdder_2432_io_ci),
    .io_s(FullAdder_2432_io_s),
    .io_co(FullAdder_2432_io_co)
  );
  FullAdder FullAdder_2433 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2433_io_a),
    .io_b(FullAdder_2433_io_b),
    .io_ci(FullAdder_2433_io_ci),
    .io_s(FullAdder_2433_io_s),
    .io_co(FullAdder_2433_io_co)
  );
  FullAdder FullAdder_2434 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2434_io_a),
    .io_b(FullAdder_2434_io_b),
    .io_ci(FullAdder_2434_io_ci),
    .io_s(FullAdder_2434_io_s),
    .io_co(FullAdder_2434_io_co)
  );
  FullAdder FullAdder_2435 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2435_io_a),
    .io_b(FullAdder_2435_io_b),
    .io_ci(FullAdder_2435_io_ci),
    .io_s(FullAdder_2435_io_s),
    .io_co(FullAdder_2435_io_co)
  );
  FullAdder FullAdder_2436 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2436_io_a),
    .io_b(FullAdder_2436_io_b),
    .io_ci(FullAdder_2436_io_ci),
    .io_s(FullAdder_2436_io_s),
    .io_co(FullAdder_2436_io_co)
  );
  FullAdder FullAdder_2437 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2437_io_a),
    .io_b(FullAdder_2437_io_b),
    .io_ci(FullAdder_2437_io_ci),
    .io_s(FullAdder_2437_io_s),
    .io_co(FullAdder_2437_io_co)
  );
  FullAdder FullAdder_2438 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2438_io_a),
    .io_b(FullAdder_2438_io_b),
    .io_ci(FullAdder_2438_io_ci),
    .io_s(FullAdder_2438_io_s),
    .io_co(FullAdder_2438_io_co)
  );
  FullAdder FullAdder_2439 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2439_io_a),
    .io_b(FullAdder_2439_io_b),
    .io_ci(FullAdder_2439_io_ci),
    .io_s(FullAdder_2439_io_s),
    .io_co(FullAdder_2439_io_co)
  );
  FullAdder FullAdder_2440 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2440_io_a),
    .io_b(FullAdder_2440_io_b),
    .io_ci(FullAdder_2440_io_ci),
    .io_s(FullAdder_2440_io_s),
    .io_co(FullAdder_2440_io_co)
  );
  FullAdder FullAdder_2441 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2441_io_a),
    .io_b(FullAdder_2441_io_b),
    .io_ci(FullAdder_2441_io_ci),
    .io_s(FullAdder_2441_io_s),
    .io_co(FullAdder_2441_io_co)
  );
  FullAdder FullAdder_2442 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2442_io_a),
    .io_b(FullAdder_2442_io_b),
    .io_ci(FullAdder_2442_io_ci),
    .io_s(FullAdder_2442_io_s),
    .io_co(FullAdder_2442_io_co)
  );
  FullAdder FullAdder_2443 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2443_io_a),
    .io_b(FullAdder_2443_io_b),
    .io_ci(FullAdder_2443_io_ci),
    .io_s(FullAdder_2443_io_s),
    .io_co(FullAdder_2443_io_co)
  );
  FullAdder FullAdder_2444 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2444_io_a),
    .io_b(FullAdder_2444_io_b),
    .io_ci(FullAdder_2444_io_ci),
    .io_s(FullAdder_2444_io_s),
    .io_co(FullAdder_2444_io_co)
  );
  FullAdder FullAdder_2445 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2445_io_a),
    .io_b(FullAdder_2445_io_b),
    .io_ci(FullAdder_2445_io_ci),
    .io_s(FullAdder_2445_io_s),
    .io_co(FullAdder_2445_io_co)
  );
  FullAdder FullAdder_2446 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2446_io_a),
    .io_b(FullAdder_2446_io_b),
    .io_ci(FullAdder_2446_io_ci),
    .io_s(FullAdder_2446_io_s),
    .io_co(FullAdder_2446_io_co)
  );
  FullAdder FullAdder_2447 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2447_io_a),
    .io_b(FullAdder_2447_io_b),
    .io_ci(FullAdder_2447_io_ci),
    .io_s(FullAdder_2447_io_s),
    .io_co(FullAdder_2447_io_co)
  );
  FullAdder FullAdder_2448 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2448_io_a),
    .io_b(FullAdder_2448_io_b),
    .io_ci(FullAdder_2448_io_ci),
    .io_s(FullAdder_2448_io_s),
    .io_co(FullAdder_2448_io_co)
  );
  FullAdder FullAdder_2449 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2449_io_a),
    .io_b(FullAdder_2449_io_b),
    .io_ci(FullAdder_2449_io_ci),
    .io_s(FullAdder_2449_io_s),
    .io_co(FullAdder_2449_io_co)
  );
  FullAdder FullAdder_2450 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2450_io_a),
    .io_b(FullAdder_2450_io_b),
    .io_ci(FullAdder_2450_io_ci),
    .io_s(FullAdder_2450_io_s),
    .io_co(FullAdder_2450_io_co)
  );
  FullAdder FullAdder_2451 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2451_io_a),
    .io_b(FullAdder_2451_io_b),
    .io_ci(FullAdder_2451_io_ci),
    .io_s(FullAdder_2451_io_s),
    .io_co(FullAdder_2451_io_co)
  );
  FullAdder FullAdder_2452 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2452_io_a),
    .io_b(FullAdder_2452_io_b),
    .io_ci(FullAdder_2452_io_ci),
    .io_s(FullAdder_2452_io_s),
    .io_co(FullAdder_2452_io_co)
  );
  FullAdder FullAdder_2453 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2453_io_a),
    .io_b(FullAdder_2453_io_b),
    .io_ci(FullAdder_2453_io_ci),
    .io_s(FullAdder_2453_io_s),
    .io_co(FullAdder_2453_io_co)
  );
  FullAdder FullAdder_2454 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2454_io_a),
    .io_b(FullAdder_2454_io_b),
    .io_ci(FullAdder_2454_io_ci),
    .io_s(FullAdder_2454_io_s),
    .io_co(FullAdder_2454_io_co)
  );
  FullAdder FullAdder_2455 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2455_io_a),
    .io_b(FullAdder_2455_io_b),
    .io_ci(FullAdder_2455_io_ci),
    .io_s(FullAdder_2455_io_s),
    .io_co(FullAdder_2455_io_co)
  );
  FullAdder FullAdder_2456 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2456_io_a),
    .io_b(FullAdder_2456_io_b),
    .io_ci(FullAdder_2456_io_ci),
    .io_s(FullAdder_2456_io_s),
    .io_co(FullAdder_2456_io_co)
  );
  FullAdder FullAdder_2457 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2457_io_a),
    .io_b(FullAdder_2457_io_b),
    .io_ci(FullAdder_2457_io_ci),
    .io_s(FullAdder_2457_io_s),
    .io_co(FullAdder_2457_io_co)
  );
  FullAdder FullAdder_2458 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2458_io_a),
    .io_b(FullAdder_2458_io_b),
    .io_ci(FullAdder_2458_io_ci),
    .io_s(FullAdder_2458_io_s),
    .io_co(FullAdder_2458_io_co)
  );
  FullAdder FullAdder_2459 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2459_io_a),
    .io_b(FullAdder_2459_io_b),
    .io_ci(FullAdder_2459_io_ci),
    .io_s(FullAdder_2459_io_s),
    .io_co(FullAdder_2459_io_co)
  );
  FullAdder FullAdder_2460 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2460_io_a),
    .io_b(FullAdder_2460_io_b),
    .io_ci(FullAdder_2460_io_ci),
    .io_s(FullAdder_2460_io_s),
    .io_co(FullAdder_2460_io_co)
  );
  FullAdder FullAdder_2461 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2461_io_a),
    .io_b(FullAdder_2461_io_b),
    .io_ci(FullAdder_2461_io_ci),
    .io_s(FullAdder_2461_io_s),
    .io_co(FullAdder_2461_io_co)
  );
  FullAdder FullAdder_2462 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2462_io_a),
    .io_b(FullAdder_2462_io_b),
    .io_ci(FullAdder_2462_io_ci),
    .io_s(FullAdder_2462_io_s),
    .io_co(FullAdder_2462_io_co)
  );
  FullAdder FullAdder_2463 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2463_io_a),
    .io_b(FullAdder_2463_io_b),
    .io_ci(FullAdder_2463_io_ci),
    .io_s(FullAdder_2463_io_s),
    .io_co(FullAdder_2463_io_co)
  );
  FullAdder FullAdder_2464 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2464_io_a),
    .io_b(FullAdder_2464_io_b),
    .io_ci(FullAdder_2464_io_ci),
    .io_s(FullAdder_2464_io_s),
    .io_co(FullAdder_2464_io_co)
  );
  FullAdder FullAdder_2465 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2465_io_a),
    .io_b(FullAdder_2465_io_b),
    .io_ci(FullAdder_2465_io_ci),
    .io_s(FullAdder_2465_io_s),
    .io_co(FullAdder_2465_io_co)
  );
  FullAdder FullAdder_2466 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2466_io_a),
    .io_b(FullAdder_2466_io_b),
    .io_ci(FullAdder_2466_io_ci),
    .io_s(FullAdder_2466_io_s),
    .io_co(FullAdder_2466_io_co)
  );
  FullAdder FullAdder_2467 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2467_io_a),
    .io_b(FullAdder_2467_io_b),
    .io_ci(FullAdder_2467_io_ci),
    .io_s(FullAdder_2467_io_s),
    .io_co(FullAdder_2467_io_co)
  );
  FullAdder FullAdder_2468 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2468_io_a),
    .io_b(FullAdder_2468_io_b),
    .io_ci(FullAdder_2468_io_ci),
    .io_s(FullAdder_2468_io_s),
    .io_co(FullAdder_2468_io_co)
  );
  FullAdder FullAdder_2469 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2469_io_a),
    .io_b(FullAdder_2469_io_b),
    .io_ci(FullAdder_2469_io_ci),
    .io_s(FullAdder_2469_io_s),
    .io_co(FullAdder_2469_io_co)
  );
  FullAdder FullAdder_2470 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2470_io_a),
    .io_b(FullAdder_2470_io_b),
    .io_ci(FullAdder_2470_io_ci),
    .io_s(FullAdder_2470_io_s),
    .io_co(FullAdder_2470_io_co)
  );
  FullAdder FullAdder_2471 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2471_io_a),
    .io_b(FullAdder_2471_io_b),
    .io_ci(FullAdder_2471_io_ci),
    .io_s(FullAdder_2471_io_s),
    .io_co(FullAdder_2471_io_co)
  );
  FullAdder FullAdder_2472 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2472_io_a),
    .io_b(FullAdder_2472_io_b),
    .io_ci(FullAdder_2472_io_ci),
    .io_s(FullAdder_2472_io_s),
    .io_co(FullAdder_2472_io_co)
  );
  FullAdder FullAdder_2473 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2473_io_a),
    .io_b(FullAdder_2473_io_b),
    .io_ci(FullAdder_2473_io_ci),
    .io_s(FullAdder_2473_io_s),
    .io_co(FullAdder_2473_io_co)
  );
  FullAdder FullAdder_2474 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2474_io_a),
    .io_b(FullAdder_2474_io_b),
    .io_ci(FullAdder_2474_io_ci),
    .io_s(FullAdder_2474_io_s),
    .io_co(FullAdder_2474_io_co)
  );
  FullAdder FullAdder_2475 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2475_io_a),
    .io_b(FullAdder_2475_io_b),
    .io_ci(FullAdder_2475_io_ci),
    .io_s(FullAdder_2475_io_s),
    .io_co(FullAdder_2475_io_co)
  );
  FullAdder FullAdder_2476 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2476_io_a),
    .io_b(FullAdder_2476_io_b),
    .io_ci(FullAdder_2476_io_ci),
    .io_s(FullAdder_2476_io_s),
    .io_co(FullAdder_2476_io_co)
  );
  FullAdder FullAdder_2477 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2477_io_a),
    .io_b(FullAdder_2477_io_b),
    .io_ci(FullAdder_2477_io_ci),
    .io_s(FullAdder_2477_io_s),
    .io_co(FullAdder_2477_io_co)
  );
  FullAdder FullAdder_2478 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2478_io_a),
    .io_b(FullAdder_2478_io_b),
    .io_ci(FullAdder_2478_io_ci),
    .io_s(FullAdder_2478_io_s),
    .io_co(FullAdder_2478_io_co)
  );
  FullAdder FullAdder_2479 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2479_io_a),
    .io_b(FullAdder_2479_io_b),
    .io_ci(FullAdder_2479_io_ci),
    .io_s(FullAdder_2479_io_s),
    .io_co(FullAdder_2479_io_co)
  );
  FullAdder FullAdder_2480 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2480_io_a),
    .io_b(FullAdder_2480_io_b),
    .io_ci(FullAdder_2480_io_ci),
    .io_s(FullAdder_2480_io_s),
    .io_co(FullAdder_2480_io_co)
  );
  FullAdder FullAdder_2481 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2481_io_a),
    .io_b(FullAdder_2481_io_b),
    .io_ci(FullAdder_2481_io_ci),
    .io_s(FullAdder_2481_io_s),
    .io_co(FullAdder_2481_io_co)
  );
  FullAdder FullAdder_2482 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2482_io_a),
    .io_b(FullAdder_2482_io_b),
    .io_ci(FullAdder_2482_io_ci),
    .io_s(FullAdder_2482_io_s),
    .io_co(FullAdder_2482_io_co)
  );
  FullAdder FullAdder_2483 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2483_io_a),
    .io_b(FullAdder_2483_io_b),
    .io_ci(FullAdder_2483_io_ci),
    .io_s(FullAdder_2483_io_s),
    .io_co(FullAdder_2483_io_co)
  );
  FullAdder FullAdder_2484 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2484_io_a),
    .io_b(FullAdder_2484_io_b),
    .io_ci(FullAdder_2484_io_ci),
    .io_s(FullAdder_2484_io_s),
    .io_co(FullAdder_2484_io_co)
  );
  FullAdder FullAdder_2485 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2485_io_a),
    .io_b(FullAdder_2485_io_b),
    .io_ci(FullAdder_2485_io_ci),
    .io_s(FullAdder_2485_io_s),
    .io_co(FullAdder_2485_io_co)
  );
  FullAdder FullAdder_2486 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2486_io_a),
    .io_b(FullAdder_2486_io_b),
    .io_ci(FullAdder_2486_io_ci),
    .io_s(FullAdder_2486_io_s),
    .io_co(FullAdder_2486_io_co)
  );
  FullAdder FullAdder_2487 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2487_io_a),
    .io_b(FullAdder_2487_io_b),
    .io_ci(FullAdder_2487_io_ci),
    .io_s(FullAdder_2487_io_s),
    .io_co(FullAdder_2487_io_co)
  );
  FullAdder FullAdder_2488 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2488_io_a),
    .io_b(FullAdder_2488_io_b),
    .io_ci(FullAdder_2488_io_ci),
    .io_s(FullAdder_2488_io_s),
    .io_co(FullAdder_2488_io_co)
  );
  FullAdder FullAdder_2489 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2489_io_a),
    .io_b(FullAdder_2489_io_b),
    .io_ci(FullAdder_2489_io_ci),
    .io_s(FullAdder_2489_io_s),
    .io_co(FullAdder_2489_io_co)
  );
  FullAdder FullAdder_2490 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2490_io_a),
    .io_b(FullAdder_2490_io_b),
    .io_ci(FullAdder_2490_io_ci),
    .io_s(FullAdder_2490_io_s),
    .io_co(FullAdder_2490_io_co)
  );
  FullAdder FullAdder_2491 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2491_io_a),
    .io_b(FullAdder_2491_io_b),
    .io_ci(FullAdder_2491_io_ci),
    .io_s(FullAdder_2491_io_s),
    .io_co(FullAdder_2491_io_co)
  );
  FullAdder FullAdder_2492 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2492_io_a),
    .io_b(FullAdder_2492_io_b),
    .io_ci(FullAdder_2492_io_ci),
    .io_s(FullAdder_2492_io_s),
    .io_co(FullAdder_2492_io_co)
  );
  FullAdder FullAdder_2493 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2493_io_a),
    .io_b(FullAdder_2493_io_b),
    .io_ci(FullAdder_2493_io_ci),
    .io_s(FullAdder_2493_io_s),
    .io_co(FullAdder_2493_io_co)
  );
  FullAdder FullAdder_2494 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2494_io_a),
    .io_b(FullAdder_2494_io_b),
    .io_ci(FullAdder_2494_io_ci),
    .io_s(FullAdder_2494_io_s),
    .io_co(FullAdder_2494_io_co)
  );
  FullAdder FullAdder_2495 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2495_io_a),
    .io_b(FullAdder_2495_io_b),
    .io_ci(FullAdder_2495_io_ci),
    .io_s(FullAdder_2495_io_s),
    .io_co(FullAdder_2495_io_co)
  );
  FullAdder FullAdder_2496 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2496_io_a),
    .io_b(FullAdder_2496_io_b),
    .io_ci(FullAdder_2496_io_ci),
    .io_s(FullAdder_2496_io_s),
    .io_co(FullAdder_2496_io_co)
  );
  FullAdder FullAdder_2497 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2497_io_a),
    .io_b(FullAdder_2497_io_b),
    .io_ci(FullAdder_2497_io_ci),
    .io_s(FullAdder_2497_io_s),
    .io_co(FullAdder_2497_io_co)
  );
  FullAdder FullAdder_2498 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2498_io_a),
    .io_b(FullAdder_2498_io_b),
    .io_ci(FullAdder_2498_io_ci),
    .io_s(FullAdder_2498_io_s),
    .io_co(FullAdder_2498_io_co)
  );
  FullAdder FullAdder_2499 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2499_io_a),
    .io_b(FullAdder_2499_io_b),
    .io_ci(FullAdder_2499_io_ci),
    .io_s(FullAdder_2499_io_s),
    .io_co(FullAdder_2499_io_co)
  );
  FullAdder FullAdder_2500 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2500_io_a),
    .io_b(FullAdder_2500_io_b),
    .io_ci(FullAdder_2500_io_ci),
    .io_s(FullAdder_2500_io_s),
    .io_co(FullAdder_2500_io_co)
  );
  FullAdder FullAdder_2501 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2501_io_a),
    .io_b(FullAdder_2501_io_b),
    .io_ci(FullAdder_2501_io_ci),
    .io_s(FullAdder_2501_io_s),
    .io_co(FullAdder_2501_io_co)
  );
  FullAdder FullAdder_2502 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2502_io_a),
    .io_b(FullAdder_2502_io_b),
    .io_ci(FullAdder_2502_io_ci),
    .io_s(FullAdder_2502_io_s),
    .io_co(FullAdder_2502_io_co)
  );
  FullAdder FullAdder_2503 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2503_io_a),
    .io_b(FullAdder_2503_io_b),
    .io_ci(FullAdder_2503_io_ci),
    .io_s(FullAdder_2503_io_s),
    .io_co(FullAdder_2503_io_co)
  );
  FullAdder FullAdder_2504 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2504_io_a),
    .io_b(FullAdder_2504_io_b),
    .io_ci(FullAdder_2504_io_ci),
    .io_s(FullAdder_2504_io_s),
    .io_co(FullAdder_2504_io_co)
  );
  FullAdder FullAdder_2505 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2505_io_a),
    .io_b(FullAdder_2505_io_b),
    .io_ci(FullAdder_2505_io_ci),
    .io_s(FullAdder_2505_io_s),
    .io_co(FullAdder_2505_io_co)
  );
  HalfAdder HalfAdder_78 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_78_io_a),
    .io_b(HalfAdder_78_io_b),
    .io_s(HalfAdder_78_io_s),
    .io_co(HalfAdder_78_io_co)
  );
  FullAdder FullAdder_2506 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2506_io_a),
    .io_b(FullAdder_2506_io_b),
    .io_ci(FullAdder_2506_io_ci),
    .io_s(FullAdder_2506_io_s),
    .io_co(FullAdder_2506_io_co)
  );
  FullAdder FullAdder_2507 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2507_io_a),
    .io_b(FullAdder_2507_io_b),
    .io_ci(FullAdder_2507_io_ci),
    .io_s(FullAdder_2507_io_s),
    .io_co(FullAdder_2507_io_co)
  );
  FullAdder FullAdder_2508 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2508_io_a),
    .io_b(FullAdder_2508_io_b),
    .io_ci(FullAdder_2508_io_ci),
    .io_s(FullAdder_2508_io_s),
    .io_co(FullAdder_2508_io_co)
  );
  FullAdder FullAdder_2509 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2509_io_a),
    .io_b(FullAdder_2509_io_b),
    .io_ci(FullAdder_2509_io_ci),
    .io_s(FullAdder_2509_io_s),
    .io_co(FullAdder_2509_io_co)
  );
  FullAdder FullAdder_2510 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2510_io_a),
    .io_b(FullAdder_2510_io_b),
    .io_ci(FullAdder_2510_io_ci),
    .io_s(FullAdder_2510_io_s),
    .io_co(FullAdder_2510_io_co)
  );
  FullAdder FullAdder_2511 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2511_io_a),
    .io_b(FullAdder_2511_io_b),
    .io_ci(FullAdder_2511_io_ci),
    .io_s(FullAdder_2511_io_s),
    .io_co(FullAdder_2511_io_co)
  );
  FullAdder FullAdder_2512 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2512_io_a),
    .io_b(FullAdder_2512_io_b),
    .io_ci(FullAdder_2512_io_ci),
    .io_s(FullAdder_2512_io_s),
    .io_co(FullAdder_2512_io_co)
  );
  FullAdder FullAdder_2513 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2513_io_a),
    .io_b(FullAdder_2513_io_b),
    .io_ci(FullAdder_2513_io_ci),
    .io_s(FullAdder_2513_io_s),
    .io_co(FullAdder_2513_io_co)
  );
  FullAdder FullAdder_2514 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2514_io_a),
    .io_b(FullAdder_2514_io_b),
    .io_ci(FullAdder_2514_io_ci),
    .io_s(FullAdder_2514_io_s),
    .io_co(FullAdder_2514_io_co)
  );
  FullAdder FullAdder_2515 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2515_io_a),
    .io_b(FullAdder_2515_io_b),
    .io_ci(FullAdder_2515_io_ci),
    .io_s(FullAdder_2515_io_s),
    .io_co(FullAdder_2515_io_co)
  );
  FullAdder FullAdder_2516 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2516_io_a),
    .io_b(FullAdder_2516_io_b),
    .io_ci(FullAdder_2516_io_ci),
    .io_s(FullAdder_2516_io_s),
    .io_co(FullAdder_2516_io_co)
  );
  FullAdder FullAdder_2517 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2517_io_a),
    .io_b(FullAdder_2517_io_b),
    .io_ci(FullAdder_2517_io_ci),
    .io_s(FullAdder_2517_io_s),
    .io_co(FullAdder_2517_io_co)
  );
  FullAdder FullAdder_2518 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2518_io_a),
    .io_b(FullAdder_2518_io_b),
    .io_ci(FullAdder_2518_io_ci),
    .io_s(FullAdder_2518_io_s),
    .io_co(FullAdder_2518_io_co)
  );
  FullAdder FullAdder_2519 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2519_io_a),
    .io_b(FullAdder_2519_io_b),
    .io_ci(FullAdder_2519_io_ci),
    .io_s(FullAdder_2519_io_s),
    .io_co(FullAdder_2519_io_co)
  );
  FullAdder FullAdder_2520 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2520_io_a),
    .io_b(FullAdder_2520_io_b),
    .io_ci(FullAdder_2520_io_ci),
    .io_s(FullAdder_2520_io_s),
    .io_co(FullAdder_2520_io_co)
  );
  FullAdder FullAdder_2521 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2521_io_a),
    .io_b(FullAdder_2521_io_b),
    .io_ci(FullAdder_2521_io_ci),
    .io_s(FullAdder_2521_io_s),
    .io_co(FullAdder_2521_io_co)
  );
  FullAdder FullAdder_2522 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2522_io_a),
    .io_b(FullAdder_2522_io_b),
    .io_ci(FullAdder_2522_io_ci),
    .io_s(FullAdder_2522_io_s),
    .io_co(FullAdder_2522_io_co)
  );
  FullAdder FullAdder_2523 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2523_io_a),
    .io_b(FullAdder_2523_io_b),
    .io_ci(FullAdder_2523_io_ci),
    .io_s(FullAdder_2523_io_s),
    .io_co(FullAdder_2523_io_co)
  );
  FullAdder FullAdder_2524 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2524_io_a),
    .io_b(FullAdder_2524_io_b),
    .io_ci(FullAdder_2524_io_ci),
    .io_s(FullAdder_2524_io_s),
    .io_co(FullAdder_2524_io_co)
  );
  FullAdder FullAdder_2525 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2525_io_a),
    .io_b(FullAdder_2525_io_b),
    .io_ci(FullAdder_2525_io_ci),
    .io_s(FullAdder_2525_io_s),
    .io_co(FullAdder_2525_io_co)
  );
  FullAdder FullAdder_2526 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2526_io_a),
    .io_b(FullAdder_2526_io_b),
    .io_ci(FullAdder_2526_io_ci),
    .io_s(FullAdder_2526_io_s),
    .io_co(FullAdder_2526_io_co)
  );
  FullAdder FullAdder_2527 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2527_io_a),
    .io_b(FullAdder_2527_io_b),
    .io_ci(FullAdder_2527_io_ci),
    .io_s(FullAdder_2527_io_s),
    .io_co(FullAdder_2527_io_co)
  );
  FullAdder FullAdder_2528 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2528_io_a),
    .io_b(FullAdder_2528_io_b),
    .io_ci(FullAdder_2528_io_ci),
    .io_s(FullAdder_2528_io_s),
    .io_co(FullAdder_2528_io_co)
  );
  FullAdder FullAdder_2529 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2529_io_a),
    .io_b(FullAdder_2529_io_b),
    .io_ci(FullAdder_2529_io_ci),
    .io_s(FullAdder_2529_io_s),
    .io_co(FullAdder_2529_io_co)
  );
  FullAdder FullAdder_2530 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2530_io_a),
    .io_b(FullAdder_2530_io_b),
    .io_ci(FullAdder_2530_io_ci),
    .io_s(FullAdder_2530_io_s),
    .io_co(FullAdder_2530_io_co)
  );
  FullAdder FullAdder_2531 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2531_io_a),
    .io_b(FullAdder_2531_io_b),
    .io_ci(FullAdder_2531_io_ci),
    .io_s(FullAdder_2531_io_s),
    .io_co(FullAdder_2531_io_co)
  );
  FullAdder FullAdder_2532 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2532_io_a),
    .io_b(FullAdder_2532_io_b),
    .io_ci(FullAdder_2532_io_ci),
    .io_s(FullAdder_2532_io_s),
    .io_co(FullAdder_2532_io_co)
  );
  FullAdder FullAdder_2533 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2533_io_a),
    .io_b(FullAdder_2533_io_b),
    .io_ci(FullAdder_2533_io_ci),
    .io_s(FullAdder_2533_io_s),
    .io_co(FullAdder_2533_io_co)
  );
  FullAdder FullAdder_2534 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2534_io_a),
    .io_b(FullAdder_2534_io_b),
    .io_ci(FullAdder_2534_io_ci),
    .io_s(FullAdder_2534_io_s),
    .io_co(FullAdder_2534_io_co)
  );
  FullAdder FullAdder_2535 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2535_io_a),
    .io_b(FullAdder_2535_io_b),
    .io_ci(FullAdder_2535_io_ci),
    .io_s(FullAdder_2535_io_s),
    .io_co(FullAdder_2535_io_co)
  );
  FullAdder FullAdder_2536 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2536_io_a),
    .io_b(FullAdder_2536_io_b),
    .io_ci(FullAdder_2536_io_ci),
    .io_s(FullAdder_2536_io_s),
    .io_co(FullAdder_2536_io_co)
  );
  FullAdder FullAdder_2537 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2537_io_a),
    .io_b(FullAdder_2537_io_b),
    .io_ci(FullAdder_2537_io_ci),
    .io_s(FullAdder_2537_io_s),
    .io_co(FullAdder_2537_io_co)
  );
  FullAdder FullAdder_2538 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2538_io_a),
    .io_b(FullAdder_2538_io_b),
    .io_ci(FullAdder_2538_io_ci),
    .io_s(FullAdder_2538_io_s),
    .io_co(FullAdder_2538_io_co)
  );
  FullAdder FullAdder_2539 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2539_io_a),
    .io_b(FullAdder_2539_io_b),
    .io_ci(FullAdder_2539_io_ci),
    .io_s(FullAdder_2539_io_s),
    .io_co(FullAdder_2539_io_co)
  );
  FullAdder FullAdder_2540 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2540_io_a),
    .io_b(FullAdder_2540_io_b),
    .io_ci(FullAdder_2540_io_ci),
    .io_s(FullAdder_2540_io_s),
    .io_co(FullAdder_2540_io_co)
  );
  FullAdder FullAdder_2541 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2541_io_a),
    .io_b(FullAdder_2541_io_b),
    .io_ci(FullAdder_2541_io_ci),
    .io_s(FullAdder_2541_io_s),
    .io_co(FullAdder_2541_io_co)
  );
  FullAdder FullAdder_2542 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2542_io_a),
    .io_b(FullAdder_2542_io_b),
    .io_ci(FullAdder_2542_io_ci),
    .io_s(FullAdder_2542_io_s),
    .io_co(FullAdder_2542_io_co)
  );
  FullAdder FullAdder_2543 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2543_io_a),
    .io_b(FullAdder_2543_io_b),
    .io_ci(FullAdder_2543_io_ci),
    .io_s(FullAdder_2543_io_s),
    .io_co(FullAdder_2543_io_co)
  );
  FullAdder FullAdder_2544 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2544_io_a),
    .io_b(FullAdder_2544_io_b),
    .io_ci(FullAdder_2544_io_ci),
    .io_s(FullAdder_2544_io_s),
    .io_co(FullAdder_2544_io_co)
  );
  FullAdder FullAdder_2545 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2545_io_a),
    .io_b(FullAdder_2545_io_b),
    .io_ci(FullAdder_2545_io_ci),
    .io_s(FullAdder_2545_io_s),
    .io_co(FullAdder_2545_io_co)
  );
  FullAdder FullAdder_2546 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2546_io_a),
    .io_b(FullAdder_2546_io_b),
    .io_ci(FullAdder_2546_io_ci),
    .io_s(FullAdder_2546_io_s),
    .io_co(FullAdder_2546_io_co)
  );
  FullAdder FullAdder_2547 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2547_io_a),
    .io_b(FullAdder_2547_io_b),
    .io_ci(FullAdder_2547_io_ci),
    .io_s(FullAdder_2547_io_s),
    .io_co(FullAdder_2547_io_co)
  );
  FullAdder FullAdder_2548 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2548_io_a),
    .io_b(FullAdder_2548_io_b),
    .io_ci(FullAdder_2548_io_ci),
    .io_s(FullAdder_2548_io_s),
    .io_co(FullAdder_2548_io_co)
  );
  FullAdder FullAdder_2549 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2549_io_a),
    .io_b(FullAdder_2549_io_b),
    .io_ci(FullAdder_2549_io_ci),
    .io_s(FullAdder_2549_io_s),
    .io_co(FullAdder_2549_io_co)
  );
  HalfAdder HalfAdder_79 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_79_io_a),
    .io_b(HalfAdder_79_io_b),
    .io_s(HalfAdder_79_io_s),
    .io_co(HalfAdder_79_io_co)
  );
  FullAdder FullAdder_2550 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2550_io_a),
    .io_b(FullAdder_2550_io_b),
    .io_ci(FullAdder_2550_io_ci),
    .io_s(FullAdder_2550_io_s),
    .io_co(FullAdder_2550_io_co)
  );
  FullAdder FullAdder_2551 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2551_io_a),
    .io_b(FullAdder_2551_io_b),
    .io_ci(FullAdder_2551_io_ci),
    .io_s(FullAdder_2551_io_s),
    .io_co(FullAdder_2551_io_co)
  );
  FullAdder FullAdder_2552 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2552_io_a),
    .io_b(FullAdder_2552_io_b),
    .io_ci(FullAdder_2552_io_ci),
    .io_s(FullAdder_2552_io_s),
    .io_co(FullAdder_2552_io_co)
  );
  FullAdder FullAdder_2553 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2553_io_a),
    .io_b(FullAdder_2553_io_b),
    .io_ci(FullAdder_2553_io_ci),
    .io_s(FullAdder_2553_io_s),
    .io_co(FullAdder_2553_io_co)
  );
  FullAdder FullAdder_2554 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2554_io_a),
    .io_b(FullAdder_2554_io_b),
    .io_ci(FullAdder_2554_io_ci),
    .io_s(FullAdder_2554_io_s),
    .io_co(FullAdder_2554_io_co)
  );
  FullAdder FullAdder_2555 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2555_io_a),
    .io_b(FullAdder_2555_io_b),
    .io_ci(FullAdder_2555_io_ci),
    .io_s(FullAdder_2555_io_s),
    .io_co(FullAdder_2555_io_co)
  );
  FullAdder FullAdder_2556 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2556_io_a),
    .io_b(FullAdder_2556_io_b),
    .io_ci(FullAdder_2556_io_ci),
    .io_s(FullAdder_2556_io_s),
    .io_co(FullAdder_2556_io_co)
  );
  FullAdder FullAdder_2557 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2557_io_a),
    .io_b(FullAdder_2557_io_b),
    .io_ci(FullAdder_2557_io_ci),
    .io_s(FullAdder_2557_io_s),
    .io_co(FullAdder_2557_io_co)
  );
  FullAdder FullAdder_2558 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2558_io_a),
    .io_b(FullAdder_2558_io_b),
    .io_ci(FullAdder_2558_io_ci),
    .io_s(FullAdder_2558_io_s),
    .io_co(FullAdder_2558_io_co)
  );
  FullAdder FullAdder_2559 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2559_io_a),
    .io_b(FullAdder_2559_io_b),
    .io_ci(FullAdder_2559_io_ci),
    .io_s(FullAdder_2559_io_s),
    .io_co(FullAdder_2559_io_co)
  );
  FullAdder FullAdder_2560 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2560_io_a),
    .io_b(FullAdder_2560_io_b),
    .io_ci(FullAdder_2560_io_ci),
    .io_s(FullAdder_2560_io_s),
    .io_co(FullAdder_2560_io_co)
  );
  FullAdder FullAdder_2561 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2561_io_a),
    .io_b(FullAdder_2561_io_b),
    .io_ci(FullAdder_2561_io_ci),
    .io_s(FullAdder_2561_io_s),
    .io_co(FullAdder_2561_io_co)
  );
  FullAdder FullAdder_2562 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2562_io_a),
    .io_b(FullAdder_2562_io_b),
    .io_ci(FullAdder_2562_io_ci),
    .io_s(FullAdder_2562_io_s),
    .io_co(FullAdder_2562_io_co)
  );
  FullAdder FullAdder_2563 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2563_io_a),
    .io_b(FullAdder_2563_io_b),
    .io_ci(FullAdder_2563_io_ci),
    .io_s(FullAdder_2563_io_s),
    .io_co(FullAdder_2563_io_co)
  );
  FullAdder FullAdder_2564 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2564_io_a),
    .io_b(FullAdder_2564_io_b),
    .io_ci(FullAdder_2564_io_ci),
    .io_s(FullAdder_2564_io_s),
    .io_co(FullAdder_2564_io_co)
  );
  FullAdder FullAdder_2565 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2565_io_a),
    .io_b(FullAdder_2565_io_b),
    .io_ci(FullAdder_2565_io_ci),
    .io_s(FullAdder_2565_io_s),
    .io_co(FullAdder_2565_io_co)
  );
  FullAdder FullAdder_2566 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2566_io_a),
    .io_b(FullAdder_2566_io_b),
    .io_ci(FullAdder_2566_io_ci),
    .io_s(FullAdder_2566_io_s),
    .io_co(FullAdder_2566_io_co)
  );
  FullAdder FullAdder_2567 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2567_io_a),
    .io_b(FullAdder_2567_io_b),
    .io_ci(FullAdder_2567_io_ci),
    .io_s(FullAdder_2567_io_s),
    .io_co(FullAdder_2567_io_co)
  );
  FullAdder FullAdder_2568 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2568_io_a),
    .io_b(FullAdder_2568_io_b),
    .io_ci(FullAdder_2568_io_ci),
    .io_s(FullAdder_2568_io_s),
    .io_co(FullAdder_2568_io_co)
  );
  FullAdder FullAdder_2569 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2569_io_a),
    .io_b(FullAdder_2569_io_b),
    .io_ci(FullAdder_2569_io_ci),
    .io_s(FullAdder_2569_io_s),
    .io_co(FullAdder_2569_io_co)
  );
  FullAdder FullAdder_2570 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2570_io_a),
    .io_b(FullAdder_2570_io_b),
    .io_ci(FullAdder_2570_io_ci),
    .io_s(FullAdder_2570_io_s),
    .io_co(FullAdder_2570_io_co)
  );
  FullAdder FullAdder_2571 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2571_io_a),
    .io_b(FullAdder_2571_io_b),
    .io_ci(FullAdder_2571_io_ci),
    .io_s(FullAdder_2571_io_s),
    .io_co(FullAdder_2571_io_co)
  );
  FullAdder FullAdder_2572 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2572_io_a),
    .io_b(FullAdder_2572_io_b),
    .io_ci(FullAdder_2572_io_ci),
    .io_s(FullAdder_2572_io_s),
    .io_co(FullAdder_2572_io_co)
  );
  FullAdder FullAdder_2573 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2573_io_a),
    .io_b(FullAdder_2573_io_b),
    .io_ci(FullAdder_2573_io_ci),
    .io_s(FullAdder_2573_io_s),
    .io_co(FullAdder_2573_io_co)
  );
  FullAdder FullAdder_2574 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2574_io_a),
    .io_b(FullAdder_2574_io_b),
    .io_ci(FullAdder_2574_io_ci),
    .io_s(FullAdder_2574_io_s),
    .io_co(FullAdder_2574_io_co)
  );
  FullAdder FullAdder_2575 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2575_io_a),
    .io_b(FullAdder_2575_io_b),
    .io_ci(FullAdder_2575_io_ci),
    .io_s(FullAdder_2575_io_s),
    .io_co(FullAdder_2575_io_co)
  );
  FullAdder FullAdder_2576 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2576_io_a),
    .io_b(FullAdder_2576_io_b),
    .io_ci(FullAdder_2576_io_ci),
    .io_s(FullAdder_2576_io_s),
    .io_co(FullAdder_2576_io_co)
  );
  FullAdder FullAdder_2577 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2577_io_a),
    .io_b(FullAdder_2577_io_b),
    .io_ci(FullAdder_2577_io_ci),
    .io_s(FullAdder_2577_io_s),
    .io_co(FullAdder_2577_io_co)
  );
  FullAdder FullAdder_2578 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2578_io_a),
    .io_b(FullAdder_2578_io_b),
    .io_ci(FullAdder_2578_io_ci),
    .io_s(FullAdder_2578_io_s),
    .io_co(FullAdder_2578_io_co)
  );
  FullAdder FullAdder_2579 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2579_io_a),
    .io_b(FullAdder_2579_io_b),
    .io_ci(FullAdder_2579_io_ci),
    .io_s(FullAdder_2579_io_s),
    .io_co(FullAdder_2579_io_co)
  );
  FullAdder FullAdder_2580 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2580_io_a),
    .io_b(FullAdder_2580_io_b),
    .io_ci(FullAdder_2580_io_ci),
    .io_s(FullAdder_2580_io_s),
    .io_co(FullAdder_2580_io_co)
  );
  FullAdder FullAdder_2581 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2581_io_a),
    .io_b(FullAdder_2581_io_b),
    .io_ci(FullAdder_2581_io_ci),
    .io_s(FullAdder_2581_io_s),
    .io_co(FullAdder_2581_io_co)
  );
  FullAdder FullAdder_2582 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2582_io_a),
    .io_b(FullAdder_2582_io_b),
    .io_ci(FullAdder_2582_io_ci),
    .io_s(FullAdder_2582_io_s),
    .io_co(FullAdder_2582_io_co)
  );
  FullAdder FullAdder_2583 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2583_io_a),
    .io_b(FullAdder_2583_io_b),
    .io_ci(FullAdder_2583_io_ci),
    .io_s(FullAdder_2583_io_s),
    .io_co(FullAdder_2583_io_co)
  );
  FullAdder FullAdder_2584 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2584_io_a),
    .io_b(FullAdder_2584_io_b),
    .io_ci(FullAdder_2584_io_ci),
    .io_s(FullAdder_2584_io_s),
    .io_co(FullAdder_2584_io_co)
  );
  FullAdder FullAdder_2585 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2585_io_a),
    .io_b(FullAdder_2585_io_b),
    .io_ci(FullAdder_2585_io_ci),
    .io_s(FullAdder_2585_io_s),
    .io_co(FullAdder_2585_io_co)
  );
  FullAdder FullAdder_2586 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2586_io_a),
    .io_b(FullAdder_2586_io_b),
    .io_ci(FullAdder_2586_io_ci),
    .io_s(FullAdder_2586_io_s),
    .io_co(FullAdder_2586_io_co)
  );
  FullAdder FullAdder_2587 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2587_io_a),
    .io_b(FullAdder_2587_io_b),
    .io_ci(FullAdder_2587_io_ci),
    .io_s(FullAdder_2587_io_s),
    .io_co(FullAdder_2587_io_co)
  );
  FullAdder FullAdder_2588 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2588_io_a),
    .io_b(FullAdder_2588_io_b),
    .io_ci(FullAdder_2588_io_ci),
    .io_s(FullAdder_2588_io_s),
    .io_co(FullAdder_2588_io_co)
  );
  FullAdder FullAdder_2589 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2589_io_a),
    .io_b(FullAdder_2589_io_b),
    .io_ci(FullAdder_2589_io_ci),
    .io_s(FullAdder_2589_io_s),
    .io_co(FullAdder_2589_io_co)
  );
  FullAdder FullAdder_2590 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2590_io_a),
    .io_b(FullAdder_2590_io_b),
    .io_ci(FullAdder_2590_io_ci),
    .io_s(FullAdder_2590_io_s),
    .io_co(FullAdder_2590_io_co)
  );
  FullAdder FullAdder_2591 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2591_io_a),
    .io_b(FullAdder_2591_io_b),
    .io_ci(FullAdder_2591_io_ci),
    .io_s(FullAdder_2591_io_s),
    .io_co(FullAdder_2591_io_co)
  );
  FullAdder FullAdder_2592 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2592_io_a),
    .io_b(FullAdder_2592_io_b),
    .io_ci(FullAdder_2592_io_ci),
    .io_s(FullAdder_2592_io_s),
    .io_co(FullAdder_2592_io_co)
  );
  FullAdder FullAdder_2593 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2593_io_a),
    .io_b(FullAdder_2593_io_b),
    .io_ci(FullAdder_2593_io_ci),
    .io_s(FullAdder_2593_io_s),
    .io_co(FullAdder_2593_io_co)
  );
  FullAdder FullAdder_2594 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2594_io_a),
    .io_b(FullAdder_2594_io_b),
    .io_ci(FullAdder_2594_io_ci),
    .io_s(FullAdder_2594_io_s),
    .io_co(FullAdder_2594_io_co)
  );
  FullAdder FullAdder_2595 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2595_io_a),
    .io_b(FullAdder_2595_io_b),
    .io_ci(FullAdder_2595_io_ci),
    .io_s(FullAdder_2595_io_s),
    .io_co(FullAdder_2595_io_co)
  );
  FullAdder FullAdder_2596 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2596_io_a),
    .io_b(FullAdder_2596_io_b),
    .io_ci(FullAdder_2596_io_ci),
    .io_s(FullAdder_2596_io_s),
    .io_co(FullAdder_2596_io_co)
  );
  FullAdder FullAdder_2597 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2597_io_a),
    .io_b(FullAdder_2597_io_b),
    .io_ci(FullAdder_2597_io_ci),
    .io_s(FullAdder_2597_io_s),
    .io_co(FullAdder_2597_io_co)
  );
  FullAdder FullAdder_2598 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2598_io_a),
    .io_b(FullAdder_2598_io_b),
    .io_ci(FullAdder_2598_io_ci),
    .io_s(FullAdder_2598_io_s),
    .io_co(FullAdder_2598_io_co)
  );
  FullAdder FullAdder_2599 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2599_io_a),
    .io_b(FullAdder_2599_io_b),
    .io_ci(FullAdder_2599_io_ci),
    .io_s(FullAdder_2599_io_s),
    .io_co(FullAdder_2599_io_co)
  );
  FullAdder FullAdder_2600 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2600_io_a),
    .io_b(FullAdder_2600_io_b),
    .io_ci(FullAdder_2600_io_ci),
    .io_s(FullAdder_2600_io_s),
    .io_co(FullAdder_2600_io_co)
  );
  FullAdder FullAdder_2601 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2601_io_a),
    .io_b(FullAdder_2601_io_b),
    .io_ci(FullAdder_2601_io_ci),
    .io_s(FullAdder_2601_io_s),
    .io_co(FullAdder_2601_io_co)
  );
  FullAdder FullAdder_2602 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2602_io_a),
    .io_b(FullAdder_2602_io_b),
    .io_ci(FullAdder_2602_io_ci),
    .io_s(FullAdder_2602_io_s),
    .io_co(FullAdder_2602_io_co)
  );
  FullAdder FullAdder_2603 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2603_io_a),
    .io_b(FullAdder_2603_io_b),
    .io_ci(FullAdder_2603_io_ci),
    .io_s(FullAdder_2603_io_s),
    .io_co(FullAdder_2603_io_co)
  );
  HalfAdder HalfAdder_80 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_80_io_a),
    .io_b(HalfAdder_80_io_b),
    .io_s(HalfAdder_80_io_s),
    .io_co(HalfAdder_80_io_co)
  );
  FullAdder FullAdder_2604 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2604_io_a),
    .io_b(FullAdder_2604_io_b),
    .io_ci(FullAdder_2604_io_ci),
    .io_s(FullAdder_2604_io_s),
    .io_co(FullAdder_2604_io_co)
  );
  FullAdder FullAdder_2605 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2605_io_a),
    .io_b(FullAdder_2605_io_b),
    .io_ci(FullAdder_2605_io_ci),
    .io_s(FullAdder_2605_io_s),
    .io_co(FullAdder_2605_io_co)
  );
  FullAdder FullAdder_2606 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2606_io_a),
    .io_b(FullAdder_2606_io_b),
    .io_ci(FullAdder_2606_io_ci),
    .io_s(FullAdder_2606_io_s),
    .io_co(FullAdder_2606_io_co)
  );
  FullAdder FullAdder_2607 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2607_io_a),
    .io_b(FullAdder_2607_io_b),
    .io_ci(FullAdder_2607_io_ci),
    .io_s(FullAdder_2607_io_s),
    .io_co(FullAdder_2607_io_co)
  );
  FullAdder FullAdder_2608 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2608_io_a),
    .io_b(FullAdder_2608_io_b),
    .io_ci(FullAdder_2608_io_ci),
    .io_s(FullAdder_2608_io_s),
    .io_co(FullAdder_2608_io_co)
  );
  FullAdder FullAdder_2609 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2609_io_a),
    .io_b(FullAdder_2609_io_b),
    .io_ci(FullAdder_2609_io_ci),
    .io_s(FullAdder_2609_io_s),
    .io_co(FullAdder_2609_io_co)
  );
  FullAdder FullAdder_2610 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2610_io_a),
    .io_b(FullAdder_2610_io_b),
    .io_ci(FullAdder_2610_io_ci),
    .io_s(FullAdder_2610_io_s),
    .io_co(FullAdder_2610_io_co)
  );
  FullAdder FullAdder_2611 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2611_io_a),
    .io_b(FullAdder_2611_io_b),
    .io_ci(FullAdder_2611_io_ci),
    .io_s(FullAdder_2611_io_s),
    .io_co(FullAdder_2611_io_co)
  );
  FullAdder FullAdder_2612 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2612_io_a),
    .io_b(FullAdder_2612_io_b),
    .io_ci(FullAdder_2612_io_ci),
    .io_s(FullAdder_2612_io_s),
    .io_co(FullAdder_2612_io_co)
  );
  FullAdder FullAdder_2613 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2613_io_a),
    .io_b(FullAdder_2613_io_b),
    .io_ci(FullAdder_2613_io_ci),
    .io_s(FullAdder_2613_io_s),
    .io_co(FullAdder_2613_io_co)
  );
  FullAdder FullAdder_2614 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2614_io_a),
    .io_b(FullAdder_2614_io_b),
    .io_ci(FullAdder_2614_io_ci),
    .io_s(FullAdder_2614_io_s),
    .io_co(FullAdder_2614_io_co)
  );
  FullAdder FullAdder_2615 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2615_io_a),
    .io_b(FullAdder_2615_io_b),
    .io_ci(FullAdder_2615_io_ci),
    .io_s(FullAdder_2615_io_s),
    .io_co(FullAdder_2615_io_co)
  );
  FullAdder FullAdder_2616 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2616_io_a),
    .io_b(FullAdder_2616_io_b),
    .io_ci(FullAdder_2616_io_ci),
    .io_s(FullAdder_2616_io_s),
    .io_co(FullAdder_2616_io_co)
  );
  FullAdder FullAdder_2617 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2617_io_a),
    .io_b(FullAdder_2617_io_b),
    .io_ci(FullAdder_2617_io_ci),
    .io_s(FullAdder_2617_io_s),
    .io_co(FullAdder_2617_io_co)
  );
  FullAdder FullAdder_2618 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2618_io_a),
    .io_b(FullAdder_2618_io_b),
    .io_ci(FullAdder_2618_io_ci),
    .io_s(FullAdder_2618_io_s),
    .io_co(FullAdder_2618_io_co)
  );
  FullAdder FullAdder_2619 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2619_io_a),
    .io_b(FullAdder_2619_io_b),
    .io_ci(FullAdder_2619_io_ci),
    .io_s(FullAdder_2619_io_s),
    .io_co(FullAdder_2619_io_co)
  );
  FullAdder FullAdder_2620 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2620_io_a),
    .io_b(FullAdder_2620_io_b),
    .io_ci(FullAdder_2620_io_ci),
    .io_s(FullAdder_2620_io_s),
    .io_co(FullAdder_2620_io_co)
  );
  FullAdder FullAdder_2621 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2621_io_a),
    .io_b(FullAdder_2621_io_b),
    .io_ci(FullAdder_2621_io_ci),
    .io_s(FullAdder_2621_io_s),
    .io_co(FullAdder_2621_io_co)
  );
  FullAdder FullAdder_2622 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2622_io_a),
    .io_b(FullAdder_2622_io_b),
    .io_ci(FullAdder_2622_io_ci),
    .io_s(FullAdder_2622_io_s),
    .io_co(FullAdder_2622_io_co)
  );
  FullAdder FullAdder_2623 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2623_io_a),
    .io_b(FullAdder_2623_io_b),
    .io_ci(FullAdder_2623_io_ci),
    .io_s(FullAdder_2623_io_s),
    .io_co(FullAdder_2623_io_co)
  );
  FullAdder FullAdder_2624 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2624_io_a),
    .io_b(FullAdder_2624_io_b),
    .io_ci(FullAdder_2624_io_ci),
    .io_s(FullAdder_2624_io_s),
    .io_co(FullAdder_2624_io_co)
  );
  FullAdder FullAdder_2625 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2625_io_a),
    .io_b(FullAdder_2625_io_b),
    .io_ci(FullAdder_2625_io_ci),
    .io_s(FullAdder_2625_io_s),
    .io_co(FullAdder_2625_io_co)
  );
  FullAdder FullAdder_2626 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2626_io_a),
    .io_b(FullAdder_2626_io_b),
    .io_ci(FullAdder_2626_io_ci),
    .io_s(FullAdder_2626_io_s),
    .io_co(FullAdder_2626_io_co)
  );
  FullAdder FullAdder_2627 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2627_io_a),
    .io_b(FullAdder_2627_io_b),
    .io_ci(FullAdder_2627_io_ci),
    .io_s(FullAdder_2627_io_s),
    .io_co(FullAdder_2627_io_co)
  );
  FullAdder FullAdder_2628 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2628_io_a),
    .io_b(FullAdder_2628_io_b),
    .io_ci(FullAdder_2628_io_ci),
    .io_s(FullAdder_2628_io_s),
    .io_co(FullAdder_2628_io_co)
  );
  FullAdder FullAdder_2629 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2629_io_a),
    .io_b(FullAdder_2629_io_b),
    .io_ci(FullAdder_2629_io_ci),
    .io_s(FullAdder_2629_io_s),
    .io_co(FullAdder_2629_io_co)
  );
  FullAdder FullAdder_2630 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2630_io_a),
    .io_b(FullAdder_2630_io_b),
    .io_ci(FullAdder_2630_io_ci),
    .io_s(FullAdder_2630_io_s),
    .io_co(FullAdder_2630_io_co)
  );
  FullAdder FullAdder_2631 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2631_io_a),
    .io_b(FullAdder_2631_io_b),
    .io_ci(FullAdder_2631_io_ci),
    .io_s(FullAdder_2631_io_s),
    .io_co(FullAdder_2631_io_co)
  );
  FullAdder FullAdder_2632 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2632_io_a),
    .io_b(FullAdder_2632_io_b),
    .io_ci(FullAdder_2632_io_ci),
    .io_s(FullAdder_2632_io_s),
    .io_co(FullAdder_2632_io_co)
  );
  FullAdder FullAdder_2633 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2633_io_a),
    .io_b(FullAdder_2633_io_b),
    .io_ci(FullAdder_2633_io_ci),
    .io_s(FullAdder_2633_io_s),
    .io_co(FullAdder_2633_io_co)
  );
  FullAdder FullAdder_2634 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2634_io_a),
    .io_b(FullAdder_2634_io_b),
    .io_ci(FullAdder_2634_io_ci),
    .io_s(FullAdder_2634_io_s),
    .io_co(FullAdder_2634_io_co)
  );
  FullAdder FullAdder_2635 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2635_io_a),
    .io_b(FullAdder_2635_io_b),
    .io_ci(FullAdder_2635_io_ci),
    .io_s(FullAdder_2635_io_s),
    .io_co(FullAdder_2635_io_co)
  );
  FullAdder FullAdder_2636 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2636_io_a),
    .io_b(FullAdder_2636_io_b),
    .io_ci(FullAdder_2636_io_ci),
    .io_s(FullAdder_2636_io_s),
    .io_co(FullAdder_2636_io_co)
  );
  FullAdder FullAdder_2637 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2637_io_a),
    .io_b(FullAdder_2637_io_b),
    .io_ci(FullAdder_2637_io_ci),
    .io_s(FullAdder_2637_io_s),
    .io_co(FullAdder_2637_io_co)
  );
  FullAdder FullAdder_2638 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2638_io_a),
    .io_b(FullAdder_2638_io_b),
    .io_ci(FullAdder_2638_io_ci),
    .io_s(FullAdder_2638_io_s),
    .io_co(FullAdder_2638_io_co)
  );
  FullAdder FullAdder_2639 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2639_io_a),
    .io_b(FullAdder_2639_io_b),
    .io_ci(FullAdder_2639_io_ci),
    .io_s(FullAdder_2639_io_s),
    .io_co(FullAdder_2639_io_co)
  );
  FullAdder FullAdder_2640 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2640_io_a),
    .io_b(FullAdder_2640_io_b),
    .io_ci(FullAdder_2640_io_ci),
    .io_s(FullAdder_2640_io_s),
    .io_co(FullAdder_2640_io_co)
  );
  FullAdder FullAdder_2641 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2641_io_a),
    .io_b(FullAdder_2641_io_b),
    .io_ci(FullAdder_2641_io_ci),
    .io_s(FullAdder_2641_io_s),
    .io_co(FullAdder_2641_io_co)
  );
  FullAdder FullAdder_2642 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2642_io_a),
    .io_b(FullAdder_2642_io_b),
    .io_ci(FullAdder_2642_io_ci),
    .io_s(FullAdder_2642_io_s),
    .io_co(FullAdder_2642_io_co)
  );
  FullAdder FullAdder_2643 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2643_io_a),
    .io_b(FullAdder_2643_io_b),
    .io_ci(FullAdder_2643_io_ci),
    .io_s(FullAdder_2643_io_s),
    .io_co(FullAdder_2643_io_co)
  );
  FullAdder FullAdder_2644 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2644_io_a),
    .io_b(FullAdder_2644_io_b),
    .io_ci(FullAdder_2644_io_ci),
    .io_s(FullAdder_2644_io_s),
    .io_co(FullAdder_2644_io_co)
  );
  HalfAdder HalfAdder_81 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_81_io_a),
    .io_b(HalfAdder_81_io_b),
    .io_s(HalfAdder_81_io_s),
    .io_co(HalfAdder_81_io_co)
  );
  FullAdder FullAdder_2645 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2645_io_a),
    .io_b(FullAdder_2645_io_b),
    .io_ci(FullAdder_2645_io_ci),
    .io_s(FullAdder_2645_io_s),
    .io_co(FullAdder_2645_io_co)
  );
  FullAdder FullAdder_2646 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2646_io_a),
    .io_b(FullAdder_2646_io_b),
    .io_ci(FullAdder_2646_io_ci),
    .io_s(FullAdder_2646_io_s),
    .io_co(FullAdder_2646_io_co)
  );
  FullAdder FullAdder_2647 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2647_io_a),
    .io_b(FullAdder_2647_io_b),
    .io_ci(FullAdder_2647_io_ci),
    .io_s(FullAdder_2647_io_s),
    .io_co(FullAdder_2647_io_co)
  );
  FullAdder FullAdder_2648 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2648_io_a),
    .io_b(FullAdder_2648_io_b),
    .io_ci(FullAdder_2648_io_ci),
    .io_s(FullAdder_2648_io_s),
    .io_co(FullAdder_2648_io_co)
  );
  FullAdder FullAdder_2649 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2649_io_a),
    .io_b(FullAdder_2649_io_b),
    .io_ci(FullAdder_2649_io_ci),
    .io_s(FullAdder_2649_io_s),
    .io_co(FullAdder_2649_io_co)
  );
  FullAdder FullAdder_2650 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2650_io_a),
    .io_b(FullAdder_2650_io_b),
    .io_ci(FullAdder_2650_io_ci),
    .io_s(FullAdder_2650_io_s),
    .io_co(FullAdder_2650_io_co)
  );
  FullAdder FullAdder_2651 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2651_io_a),
    .io_b(FullAdder_2651_io_b),
    .io_ci(FullAdder_2651_io_ci),
    .io_s(FullAdder_2651_io_s),
    .io_co(FullAdder_2651_io_co)
  );
  FullAdder FullAdder_2652 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2652_io_a),
    .io_b(FullAdder_2652_io_b),
    .io_ci(FullAdder_2652_io_ci),
    .io_s(FullAdder_2652_io_s),
    .io_co(FullAdder_2652_io_co)
  );
  FullAdder FullAdder_2653 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2653_io_a),
    .io_b(FullAdder_2653_io_b),
    .io_ci(FullAdder_2653_io_ci),
    .io_s(FullAdder_2653_io_s),
    .io_co(FullAdder_2653_io_co)
  );
  FullAdder FullAdder_2654 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2654_io_a),
    .io_b(FullAdder_2654_io_b),
    .io_ci(FullAdder_2654_io_ci),
    .io_s(FullAdder_2654_io_s),
    .io_co(FullAdder_2654_io_co)
  );
  FullAdder FullAdder_2655 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2655_io_a),
    .io_b(FullAdder_2655_io_b),
    .io_ci(FullAdder_2655_io_ci),
    .io_s(FullAdder_2655_io_s),
    .io_co(FullAdder_2655_io_co)
  );
  FullAdder FullAdder_2656 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2656_io_a),
    .io_b(FullAdder_2656_io_b),
    .io_ci(FullAdder_2656_io_ci),
    .io_s(FullAdder_2656_io_s),
    .io_co(FullAdder_2656_io_co)
  );
  FullAdder FullAdder_2657 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2657_io_a),
    .io_b(FullAdder_2657_io_b),
    .io_ci(FullAdder_2657_io_ci),
    .io_s(FullAdder_2657_io_s),
    .io_co(FullAdder_2657_io_co)
  );
  FullAdder FullAdder_2658 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2658_io_a),
    .io_b(FullAdder_2658_io_b),
    .io_ci(FullAdder_2658_io_ci),
    .io_s(FullAdder_2658_io_s),
    .io_co(FullAdder_2658_io_co)
  );
  FullAdder FullAdder_2659 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2659_io_a),
    .io_b(FullAdder_2659_io_b),
    .io_ci(FullAdder_2659_io_ci),
    .io_s(FullAdder_2659_io_s),
    .io_co(FullAdder_2659_io_co)
  );
  FullAdder FullAdder_2660 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2660_io_a),
    .io_b(FullAdder_2660_io_b),
    .io_ci(FullAdder_2660_io_ci),
    .io_s(FullAdder_2660_io_s),
    .io_co(FullAdder_2660_io_co)
  );
  FullAdder FullAdder_2661 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2661_io_a),
    .io_b(FullAdder_2661_io_b),
    .io_ci(FullAdder_2661_io_ci),
    .io_s(FullAdder_2661_io_s),
    .io_co(FullAdder_2661_io_co)
  );
  FullAdder FullAdder_2662 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2662_io_a),
    .io_b(FullAdder_2662_io_b),
    .io_ci(FullAdder_2662_io_ci),
    .io_s(FullAdder_2662_io_s),
    .io_co(FullAdder_2662_io_co)
  );
  FullAdder FullAdder_2663 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2663_io_a),
    .io_b(FullAdder_2663_io_b),
    .io_ci(FullAdder_2663_io_ci),
    .io_s(FullAdder_2663_io_s),
    .io_co(FullAdder_2663_io_co)
  );
  FullAdder FullAdder_2664 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2664_io_a),
    .io_b(FullAdder_2664_io_b),
    .io_ci(FullAdder_2664_io_ci),
    .io_s(FullAdder_2664_io_s),
    .io_co(FullAdder_2664_io_co)
  );
  FullAdder FullAdder_2665 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2665_io_a),
    .io_b(FullAdder_2665_io_b),
    .io_ci(FullAdder_2665_io_ci),
    .io_s(FullAdder_2665_io_s),
    .io_co(FullAdder_2665_io_co)
  );
  FullAdder FullAdder_2666 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2666_io_a),
    .io_b(FullAdder_2666_io_b),
    .io_ci(FullAdder_2666_io_ci),
    .io_s(FullAdder_2666_io_s),
    .io_co(FullAdder_2666_io_co)
  );
  FullAdder FullAdder_2667 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2667_io_a),
    .io_b(FullAdder_2667_io_b),
    .io_ci(FullAdder_2667_io_ci),
    .io_s(FullAdder_2667_io_s),
    .io_co(FullAdder_2667_io_co)
  );
  FullAdder FullAdder_2668 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2668_io_a),
    .io_b(FullAdder_2668_io_b),
    .io_ci(FullAdder_2668_io_ci),
    .io_s(FullAdder_2668_io_s),
    .io_co(FullAdder_2668_io_co)
  );
  FullAdder FullAdder_2669 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2669_io_a),
    .io_b(FullAdder_2669_io_b),
    .io_ci(FullAdder_2669_io_ci),
    .io_s(FullAdder_2669_io_s),
    .io_co(FullAdder_2669_io_co)
  );
  FullAdder FullAdder_2670 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2670_io_a),
    .io_b(FullAdder_2670_io_b),
    .io_ci(FullAdder_2670_io_ci),
    .io_s(FullAdder_2670_io_s),
    .io_co(FullAdder_2670_io_co)
  );
  FullAdder FullAdder_2671 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2671_io_a),
    .io_b(FullAdder_2671_io_b),
    .io_ci(FullAdder_2671_io_ci),
    .io_s(FullAdder_2671_io_s),
    .io_co(FullAdder_2671_io_co)
  );
  FullAdder FullAdder_2672 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2672_io_a),
    .io_b(FullAdder_2672_io_b),
    .io_ci(FullAdder_2672_io_ci),
    .io_s(FullAdder_2672_io_s),
    .io_co(FullAdder_2672_io_co)
  );
  FullAdder FullAdder_2673 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2673_io_a),
    .io_b(FullAdder_2673_io_b),
    .io_ci(FullAdder_2673_io_ci),
    .io_s(FullAdder_2673_io_s),
    .io_co(FullAdder_2673_io_co)
  );
  FullAdder FullAdder_2674 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2674_io_a),
    .io_b(FullAdder_2674_io_b),
    .io_ci(FullAdder_2674_io_ci),
    .io_s(FullAdder_2674_io_s),
    .io_co(FullAdder_2674_io_co)
  );
  FullAdder FullAdder_2675 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2675_io_a),
    .io_b(FullAdder_2675_io_b),
    .io_ci(FullAdder_2675_io_ci),
    .io_s(FullAdder_2675_io_s),
    .io_co(FullAdder_2675_io_co)
  );
  FullAdder FullAdder_2676 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2676_io_a),
    .io_b(FullAdder_2676_io_b),
    .io_ci(FullAdder_2676_io_ci),
    .io_s(FullAdder_2676_io_s),
    .io_co(FullAdder_2676_io_co)
  );
  FullAdder FullAdder_2677 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2677_io_a),
    .io_b(FullAdder_2677_io_b),
    .io_ci(FullAdder_2677_io_ci),
    .io_s(FullAdder_2677_io_s),
    .io_co(FullAdder_2677_io_co)
  );
  FullAdder FullAdder_2678 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2678_io_a),
    .io_b(FullAdder_2678_io_b),
    .io_ci(FullAdder_2678_io_ci),
    .io_s(FullAdder_2678_io_s),
    .io_co(FullAdder_2678_io_co)
  );
  FullAdder FullAdder_2679 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2679_io_a),
    .io_b(FullAdder_2679_io_b),
    .io_ci(FullAdder_2679_io_ci),
    .io_s(FullAdder_2679_io_s),
    .io_co(FullAdder_2679_io_co)
  );
  FullAdder FullAdder_2680 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2680_io_a),
    .io_b(FullAdder_2680_io_b),
    .io_ci(FullAdder_2680_io_ci),
    .io_s(FullAdder_2680_io_s),
    .io_co(FullAdder_2680_io_co)
  );
  FullAdder FullAdder_2681 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2681_io_a),
    .io_b(FullAdder_2681_io_b),
    .io_ci(FullAdder_2681_io_ci),
    .io_s(FullAdder_2681_io_s),
    .io_co(FullAdder_2681_io_co)
  );
  FullAdder FullAdder_2682 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2682_io_a),
    .io_b(FullAdder_2682_io_b),
    .io_ci(FullAdder_2682_io_ci),
    .io_s(FullAdder_2682_io_s),
    .io_co(FullAdder_2682_io_co)
  );
  FullAdder FullAdder_2683 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2683_io_a),
    .io_b(FullAdder_2683_io_b),
    .io_ci(FullAdder_2683_io_ci),
    .io_s(FullAdder_2683_io_s),
    .io_co(FullAdder_2683_io_co)
  );
  FullAdder FullAdder_2684 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2684_io_a),
    .io_b(FullAdder_2684_io_b),
    .io_ci(FullAdder_2684_io_ci),
    .io_s(FullAdder_2684_io_s),
    .io_co(FullAdder_2684_io_co)
  );
  FullAdder FullAdder_2685 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2685_io_a),
    .io_b(FullAdder_2685_io_b),
    .io_ci(FullAdder_2685_io_ci),
    .io_s(FullAdder_2685_io_s),
    .io_co(FullAdder_2685_io_co)
  );
  FullAdder FullAdder_2686 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2686_io_a),
    .io_b(FullAdder_2686_io_b),
    .io_ci(FullAdder_2686_io_ci),
    .io_s(FullAdder_2686_io_s),
    .io_co(FullAdder_2686_io_co)
  );
  FullAdder FullAdder_2687 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2687_io_a),
    .io_b(FullAdder_2687_io_b),
    .io_ci(FullAdder_2687_io_ci),
    .io_s(FullAdder_2687_io_s),
    .io_co(FullAdder_2687_io_co)
  );
  FullAdder FullAdder_2688 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2688_io_a),
    .io_b(FullAdder_2688_io_b),
    .io_ci(FullAdder_2688_io_ci),
    .io_s(FullAdder_2688_io_s),
    .io_co(FullAdder_2688_io_co)
  );
  FullAdder FullAdder_2689 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2689_io_a),
    .io_b(FullAdder_2689_io_b),
    .io_ci(FullAdder_2689_io_ci),
    .io_s(FullAdder_2689_io_s),
    .io_co(FullAdder_2689_io_co)
  );
  FullAdder FullAdder_2690 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2690_io_a),
    .io_b(FullAdder_2690_io_b),
    .io_ci(FullAdder_2690_io_ci),
    .io_s(FullAdder_2690_io_s),
    .io_co(FullAdder_2690_io_co)
  );
  FullAdder FullAdder_2691 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2691_io_a),
    .io_b(FullAdder_2691_io_b),
    .io_ci(FullAdder_2691_io_ci),
    .io_s(FullAdder_2691_io_s),
    .io_co(FullAdder_2691_io_co)
  );
  HalfAdder HalfAdder_82 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_82_io_a),
    .io_b(HalfAdder_82_io_b),
    .io_s(HalfAdder_82_io_s),
    .io_co(HalfAdder_82_io_co)
  );
  FullAdder FullAdder_2692 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2692_io_a),
    .io_b(FullAdder_2692_io_b),
    .io_ci(FullAdder_2692_io_ci),
    .io_s(FullAdder_2692_io_s),
    .io_co(FullAdder_2692_io_co)
  );
  FullAdder FullAdder_2693 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2693_io_a),
    .io_b(FullAdder_2693_io_b),
    .io_ci(FullAdder_2693_io_ci),
    .io_s(FullAdder_2693_io_s),
    .io_co(FullAdder_2693_io_co)
  );
  FullAdder FullAdder_2694 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2694_io_a),
    .io_b(FullAdder_2694_io_b),
    .io_ci(FullAdder_2694_io_ci),
    .io_s(FullAdder_2694_io_s),
    .io_co(FullAdder_2694_io_co)
  );
  FullAdder FullAdder_2695 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2695_io_a),
    .io_b(FullAdder_2695_io_b),
    .io_ci(FullAdder_2695_io_ci),
    .io_s(FullAdder_2695_io_s),
    .io_co(FullAdder_2695_io_co)
  );
  FullAdder FullAdder_2696 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2696_io_a),
    .io_b(FullAdder_2696_io_b),
    .io_ci(FullAdder_2696_io_ci),
    .io_s(FullAdder_2696_io_s),
    .io_co(FullAdder_2696_io_co)
  );
  HalfAdder HalfAdder_83 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_83_io_a),
    .io_b(HalfAdder_83_io_b),
    .io_s(HalfAdder_83_io_s),
    .io_co(HalfAdder_83_io_co)
  );
  FullAdder FullAdder_2697 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2697_io_a),
    .io_b(FullAdder_2697_io_b),
    .io_ci(FullAdder_2697_io_ci),
    .io_s(FullAdder_2697_io_s),
    .io_co(FullAdder_2697_io_co)
  );
  FullAdder FullAdder_2698 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2698_io_a),
    .io_b(FullAdder_2698_io_b),
    .io_ci(FullAdder_2698_io_ci),
    .io_s(FullAdder_2698_io_s),
    .io_co(FullAdder_2698_io_co)
  );
  FullAdder FullAdder_2699 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2699_io_a),
    .io_b(FullAdder_2699_io_b),
    .io_ci(FullAdder_2699_io_ci),
    .io_s(FullAdder_2699_io_s),
    .io_co(FullAdder_2699_io_co)
  );
  FullAdder FullAdder_2700 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2700_io_a),
    .io_b(FullAdder_2700_io_b),
    .io_ci(FullAdder_2700_io_ci),
    .io_s(FullAdder_2700_io_s),
    .io_co(FullAdder_2700_io_co)
  );
  FullAdder FullAdder_2701 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2701_io_a),
    .io_b(FullAdder_2701_io_b),
    .io_ci(FullAdder_2701_io_ci),
    .io_s(FullAdder_2701_io_s),
    .io_co(FullAdder_2701_io_co)
  );
  FullAdder FullAdder_2702 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2702_io_a),
    .io_b(FullAdder_2702_io_b),
    .io_ci(FullAdder_2702_io_ci),
    .io_s(FullAdder_2702_io_s),
    .io_co(FullAdder_2702_io_co)
  );
  FullAdder FullAdder_2703 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2703_io_a),
    .io_b(FullAdder_2703_io_b),
    .io_ci(FullAdder_2703_io_ci),
    .io_s(FullAdder_2703_io_s),
    .io_co(FullAdder_2703_io_co)
  );
  FullAdder FullAdder_2704 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2704_io_a),
    .io_b(FullAdder_2704_io_b),
    .io_ci(FullAdder_2704_io_ci),
    .io_s(FullAdder_2704_io_s),
    .io_co(FullAdder_2704_io_co)
  );
  FullAdder FullAdder_2705 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2705_io_a),
    .io_b(FullAdder_2705_io_b),
    .io_ci(FullAdder_2705_io_ci),
    .io_s(FullAdder_2705_io_s),
    .io_co(FullAdder_2705_io_co)
  );
  FullAdder FullAdder_2706 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2706_io_a),
    .io_b(FullAdder_2706_io_b),
    .io_ci(FullAdder_2706_io_ci),
    .io_s(FullAdder_2706_io_s),
    .io_co(FullAdder_2706_io_co)
  );
  FullAdder FullAdder_2707 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2707_io_a),
    .io_b(FullAdder_2707_io_b),
    .io_ci(FullAdder_2707_io_ci),
    .io_s(FullAdder_2707_io_s),
    .io_co(FullAdder_2707_io_co)
  );
  FullAdder FullAdder_2708 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2708_io_a),
    .io_b(FullAdder_2708_io_b),
    .io_ci(FullAdder_2708_io_ci),
    .io_s(FullAdder_2708_io_s),
    .io_co(FullAdder_2708_io_co)
  );
  FullAdder FullAdder_2709 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2709_io_a),
    .io_b(FullAdder_2709_io_b),
    .io_ci(FullAdder_2709_io_ci),
    .io_s(FullAdder_2709_io_s),
    .io_co(FullAdder_2709_io_co)
  );
  FullAdder FullAdder_2710 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2710_io_a),
    .io_b(FullAdder_2710_io_b),
    .io_ci(FullAdder_2710_io_ci),
    .io_s(FullAdder_2710_io_s),
    .io_co(FullAdder_2710_io_co)
  );
  FullAdder FullAdder_2711 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2711_io_a),
    .io_b(FullAdder_2711_io_b),
    .io_ci(FullAdder_2711_io_ci),
    .io_s(FullAdder_2711_io_s),
    .io_co(FullAdder_2711_io_co)
  );
  FullAdder FullAdder_2712 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2712_io_a),
    .io_b(FullAdder_2712_io_b),
    .io_ci(FullAdder_2712_io_ci),
    .io_s(FullAdder_2712_io_s),
    .io_co(FullAdder_2712_io_co)
  );
  FullAdder FullAdder_2713 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2713_io_a),
    .io_b(FullAdder_2713_io_b),
    .io_ci(FullAdder_2713_io_ci),
    .io_s(FullAdder_2713_io_s),
    .io_co(FullAdder_2713_io_co)
  );
  FullAdder FullAdder_2714 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2714_io_a),
    .io_b(FullAdder_2714_io_b),
    .io_ci(FullAdder_2714_io_ci),
    .io_s(FullAdder_2714_io_s),
    .io_co(FullAdder_2714_io_co)
  );
  FullAdder FullAdder_2715 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2715_io_a),
    .io_b(FullAdder_2715_io_b),
    .io_ci(FullAdder_2715_io_ci),
    .io_s(FullAdder_2715_io_s),
    .io_co(FullAdder_2715_io_co)
  );
  FullAdder FullAdder_2716 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2716_io_a),
    .io_b(FullAdder_2716_io_b),
    .io_ci(FullAdder_2716_io_ci),
    .io_s(FullAdder_2716_io_s),
    .io_co(FullAdder_2716_io_co)
  );
  FullAdder FullAdder_2717 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2717_io_a),
    .io_b(FullAdder_2717_io_b),
    .io_ci(FullAdder_2717_io_ci),
    .io_s(FullAdder_2717_io_s),
    .io_co(FullAdder_2717_io_co)
  );
  FullAdder FullAdder_2718 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2718_io_a),
    .io_b(FullAdder_2718_io_b),
    .io_ci(FullAdder_2718_io_ci),
    .io_s(FullAdder_2718_io_s),
    .io_co(FullAdder_2718_io_co)
  );
  FullAdder FullAdder_2719 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2719_io_a),
    .io_b(FullAdder_2719_io_b),
    .io_ci(FullAdder_2719_io_ci),
    .io_s(FullAdder_2719_io_s),
    .io_co(FullAdder_2719_io_co)
  );
  FullAdder FullAdder_2720 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2720_io_a),
    .io_b(FullAdder_2720_io_b),
    .io_ci(FullAdder_2720_io_ci),
    .io_s(FullAdder_2720_io_s),
    .io_co(FullAdder_2720_io_co)
  );
  FullAdder FullAdder_2721 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2721_io_a),
    .io_b(FullAdder_2721_io_b),
    .io_ci(FullAdder_2721_io_ci),
    .io_s(FullAdder_2721_io_s),
    .io_co(FullAdder_2721_io_co)
  );
  FullAdder FullAdder_2722 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2722_io_a),
    .io_b(FullAdder_2722_io_b),
    .io_ci(FullAdder_2722_io_ci),
    .io_s(FullAdder_2722_io_s),
    .io_co(FullAdder_2722_io_co)
  );
  FullAdder FullAdder_2723 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2723_io_a),
    .io_b(FullAdder_2723_io_b),
    .io_ci(FullAdder_2723_io_ci),
    .io_s(FullAdder_2723_io_s),
    .io_co(FullAdder_2723_io_co)
  );
  FullAdder FullAdder_2724 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2724_io_a),
    .io_b(FullAdder_2724_io_b),
    .io_ci(FullAdder_2724_io_ci),
    .io_s(FullAdder_2724_io_s),
    .io_co(FullAdder_2724_io_co)
  );
  HalfAdder HalfAdder_84 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_84_io_a),
    .io_b(HalfAdder_84_io_b),
    .io_s(HalfAdder_84_io_s),
    .io_co(HalfAdder_84_io_co)
  );
  FullAdder FullAdder_2725 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2725_io_a),
    .io_b(FullAdder_2725_io_b),
    .io_ci(FullAdder_2725_io_ci),
    .io_s(FullAdder_2725_io_s),
    .io_co(FullAdder_2725_io_co)
  );
  FullAdder FullAdder_2726 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2726_io_a),
    .io_b(FullAdder_2726_io_b),
    .io_ci(FullAdder_2726_io_ci),
    .io_s(FullAdder_2726_io_s),
    .io_co(FullAdder_2726_io_co)
  );
  FullAdder FullAdder_2727 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2727_io_a),
    .io_b(FullAdder_2727_io_b),
    .io_ci(FullAdder_2727_io_ci),
    .io_s(FullAdder_2727_io_s),
    .io_co(FullAdder_2727_io_co)
  );
  FullAdder FullAdder_2728 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2728_io_a),
    .io_b(FullAdder_2728_io_b),
    .io_ci(FullAdder_2728_io_ci),
    .io_s(FullAdder_2728_io_s),
    .io_co(FullAdder_2728_io_co)
  );
  FullAdder FullAdder_2729 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2729_io_a),
    .io_b(FullAdder_2729_io_b),
    .io_ci(FullAdder_2729_io_ci),
    .io_s(FullAdder_2729_io_s),
    .io_co(FullAdder_2729_io_co)
  );
  FullAdder FullAdder_2730 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2730_io_a),
    .io_b(FullAdder_2730_io_b),
    .io_ci(FullAdder_2730_io_ci),
    .io_s(FullAdder_2730_io_s),
    .io_co(FullAdder_2730_io_co)
  );
  FullAdder FullAdder_2731 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2731_io_a),
    .io_b(FullAdder_2731_io_b),
    .io_ci(FullAdder_2731_io_ci),
    .io_s(FullAdder_2731_io_s),
    .io_co(FullAdder_2731_io_co)
  );
  FullAdder FullAdder_2732 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2732_io_a),
    .io_b(FullAdder_2732_io_b),
    .io_ci(FullAdder_2732_io_ci),
    .io_s(FullAdder_2732_io_s),
    .io_co(FullAdder_2732_io_co)
  );
  FullAdder FullAdder_2733 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2733_io_a),
    .io_b(FullAdder_2733_io_b),
    .io_ci(FullAdder_2733_io_ci),
    .io_s(FullAdder_2733_io_s),
    .io_co(FullAdder_2733_io_co)
  );
  FullAdder FullAdder_2734 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2734_io_a),
    .io_b(FullAdder_2734_io_b),
    .io_ci(FullAdder_2734_io_ci),
    .io_s(FullAdder_2734_io_s),
    .io_co(FullAdder_2734_io_co)
  );
  FullAdder FullAdder_2735 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2735_io_a),
    .io_b(FullAdder_2735_io_b),
    .io_ci(FullAdder_2735_io_ci),
    .io_s(FullAdder_2735_io_s),
    .io_co(FullAdder_2735_io_co)
  );
  FullAdder FullAdder_2736 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2736_io_a),
    .io_b(FullAdder_2736_io_b),
    .io_ci(FullAdder_2736_io_ci),
    .io_s(FullAdder_2736_io_s),
    .io_co(FullAdder_2736_io_co)
  );
  FullAdder FullAdder_2737 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2737_io_a),
    .io_b(FullAdder_2737_io_b),
    .io_ci(FullAdder_2737_io_ci),
    .io_s(FullAdder_2737_io_s),
    .io_co(FullAdder_2737_io_co)
  );
  FullAdder FullAdder_2738 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2738_io_a),
    .io_b(FullAdder_2738_io_b),
    .io_ci(FullAdder_2738_io_ci),
    .io_s(FullAdder_2738_io_s),
    .io_co(FullAdder_2738_io_co)
  );
  FullAdder FullAdder_2739 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2739_io_a),
    .io_b(FullAdder_2739_io_b),
    .io_ci(FullAdder_2739_io_ci),
    .io_s(FullAdder_2739_io_s),
    .io_co(FullAdder_2739_io_co)
  );
  FullAdder FullAdder_2740 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2740_io_a),
    .io_b(FullAdder_2740_io_b),
    .io_ci(FullAdder_2740_io_ci),
    .io_s(FullAdder_2740_io_s),
    .io_co(FullAdder_2740_io_co)
  );
  FullAdder FullAdder_2741 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2741_io_a),
    .io_b(FullAdder_2741_io_b),
    .io_ci(FullAdder_2741_io_ci),
    .io_s(FullAdder_2741_io_s),
    .io_co(FullAdder_2741_io_co)
  );
  FullAdder FullAdder_2742 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2742_io_a),
    .io_b(FullAdder_2742_io_b),
    .io_ci(FullAdder_2742_io_ci),
    .io_s(FullAdder_2742_io_s),
    .io_co(FullAdder_2742_io_co)
  );
  FullAdder FullAdder_2743 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2743_io_a),
    .io_b(FullAdder_2743_io_b),
    .io_ci(FullAdder_2743_io_ci),
    .io_s(FullAdder_2743_io_s),
    .io_co(FullAdder_2743_io_co)
  );
  FullAdder FullAdder_2744 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2744_io_a),
    .io_b(FullAdder_2744_io_b),
    .io_ci(FullAdder_2744_io_ci),
    .io_s(FullAdder_2744_io_s),
    .io_co(FullAdder_2744_io_co)
  );
  FullAdder FullAdder_2745 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2745_io_a),
    .io_b(FullAdder_2745_io_b),
    .io_ci(FullAdder_2745_io_ci),
    .io_s(FullAdder_2745_io_s),
    .io_co(FullAdder_2745_io_co)
  );
  FullAdder FullAdder_2746 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2746_io_a),
    .io_b(FullAdder_2746_io_b),
    .io_ci(FullAdder_2746_io_ci),
    .io_s(FullAdder_2746_io_s),
    .io_co(FullAdder_2746_io_co)
  );
  FullAdder FullAdder_2747 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2747_io_a),
    .io_b(FullAdder_2747_io_b),
    .io_ci(FullAdder_2747_io_ci),
    .io_s(FullAdder_2747_io_s),
    .io_co(FullAdder_2747_io_co)
  );
  FullAdder FullAdder_2748 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2748_io_a),
    .io_b(FullAdder_2748_io_b),
    .io_ci(FullAdder_2748_io_ci),
    .io_s(FullAdder_2748_io_s),
    .io_co(FullAdder_2748_io_co)
  );
  FullAdder FullAdder_2749 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2749_io_a),
    .io_b(FullAdder_2749_io_b),
    .io_ci(FullAdder_2749_io_ci),
    .io_s(FullAdder_2749_io_s),
    .io_co(FullAdder_2749_io_co)
  );
  FullAdder FullAdder_2750 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2750_io_a),
    .io_b(FullAdder_2750_io_b),
    .io_ci(FullAdder_2750_io_ci),
    .io_s(FullAdder_2750_io_s),
    .io_co(FullAdder_2750_io_co)
  );
  HalfAdder HalfAdder_85 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_85_io_a),
    .io_b(HalfAdder_85_io_b),
    .io_s(HalfAdder_85_io_s),
    .io_co(HalfAdder_85_io_co)
  );
  FullAdder FullAdder_2751 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2751_io_a),
    .io_b(FullAdder_2751_io_b),
    .io_ci(FullAdder_2751_io_ci),
    .io_s(FullAdder_2751_io_s),
    .io_co(FullAdder_2751_io_co)
  );
  FullAdder FullAdder_2752 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2752_io_a),
    .io_b(FullAdder_2752_io_b),
    .io_ci(FullAdder_2752_io_ci),
    .io_s(FullAdder_2752_io_s),
    .io_co(FullAdder_2752_io_co)
  );
  FullAdder FullAdder_2753 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2753_io_a),
    .io_b(FullAdder_2753_io_b),
    .io_ci(FullAdder_2753_io_ci),
    .io_s(FullAdder_2753_io_s),
    .io_co(FullAdder_2753_io_co)
  );
  FullAdder FullAdder_2754 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2754_io_a),
    .io_b(FullAdder_2754_io_b),
    .io_ci(FullAdder_2754_io_ci),
    .io_s(FullAdder_2754_io_s),
    .io_co(FullAdder_2754_io_co)
  );
  FullAdder FullAdder_2755 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2755_io_a),
    .io_b(FullAdder_2755_io_b),
    .io_ci(FullAdder_2755_io_ci),
    .io_s(FullAdder_2755_io_s),
    .io_co(FullAdder_2755_io_co)
  );
  FullAdder FullAdder_2756 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2756_io_a),
    .io_b(FullAdder_2756_io_b),
    .io_ci(FullAdder_2756_io_ci),
    .io_s(FullAdder_2756_io_s),
    .io_co(FullAdder_2756_io_co)
  );
  FullAdder FullAdder_2757 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2757_io_a),
    .io_b(FullAdder_2757_io_b),
    .io_ci(FullAdder_2757_io_ci),
    .io_s(FullAdder_2757_io_s),
    .io_co(FullAdder_2757_io_co)
  );
  FullAdder FullAdder_2758 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2758_io_a),
    .io_b(FullAdder_2758_io_b),
    .io_ci(FullAdder_2758_io_ci),
    .io_s(FullAdder_2758_io_s),
    .io_co(FullAdder_2758_io_co)
  );
  FullAdder FullAdder_2759 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2759_io_a),
    .io_b(FullAdder_2759_io_b),
    .io_ci(FullAdder_2759_io_ci),
    .io_s(FullAdder_2759_io_s),
    .io_co(FullAdder_2759_io_co)
  );
  FullAdder FullAdder_2760 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2760_io_a),
    .io_b(FullAdder_2760_io_b),
    .io_ci(FullAdder_2760_io_ci),
    .io_s(FullAdder_2760_io_s),
    .io_co(FullAdder_2760_io_co)
  );
  FullAdder FullAdder_2761 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2761_io_a),
    .io_b(FullAdder_2761_io_b),
    .io_ci(FullAdder_2761_io_ci),
    .io_s(FullAdder_2761_io_s),
    .io_co(FullAdder_2761_io_co)
  );
  FullAdder FullAdder_2762 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2762_io_a),
    .io_b(FullAdder_2762_io_b),
    .io_ci(FullAdder_2762_io_ci),
    .io_s(FullAdder_2762_io_s),
    .io_co(FullAdder_2762_io_co)
  );
  FullAdder FullAdder_2763 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2763_io_a),
    .io_b(FullAdder_2763_io_b),
    .io_ci(FullAdder_2763_io_ci),
    .io_s(FullAdder_2763_io_s),
    .io_co(FullAdder_2763_io_co)
  );
  FullAdder FullAdder_2764 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2764_io_a),
    .io_b(FullAdder_2764_io_b),
    .io_ci(FullAdder_2764_io_ci),
    .io_s(FullAdder_2764_io_s),
    .io_co(FullAdder_2764_io_co)
  );
  FullAdder FullAdder_2765 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2765_io_a),
    .io_b(FullAdder_2765_io_b),
    .io_ci(FullAdder_2765_io_ci),
    .io_s(FullAdder_2765_io_s),
    .io_co(FullAdder_2765_io_co)
  );
  FullAdder FullAdder_2766 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2766_io_a),
    .io_b(FullAdder_2766_io_b),
    .io_ci(FullAdder_2766_io_ci),
    .io_s(FullAdder_2766_io_s),
    .io_co(FullAdder_2766_io_co)
  );
  FullAdder FullAdder_2767 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2767_io_a),
    .io_b(FullAdder_2767_io_b),
    .io_ci(FullAdder_2767_io_ci),
    .io_s(FullAdder_2767_io_s),
    .io_co(FullAdder_2767_io_co)
  );
  FullAdder FullAdder_2768 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2768_io_a),
    .io_b(FullAdder_2768_io_b),
    .io_ci(FullAdder_2768_io_ci),
    .io_s(FullAdder_2768_io_s),
    .io_co(FullAdder_2768_io_co)
  );
  FullAdder FullAdder_2769 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2769_io_a),
    .io_b(FullAdder_2769_io_b),
    .io_ci(FullAdder_2769_io_ci),
    .io_s(FullAdder_2769_io_s),
    .io_co(FullAdder_2769_io_co)
  );
  HalfAdder HalfAdder_86 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_86_io_a),
    .io_b(HalfAdder_86_io_b),
    .io_s(HalfAdder_86_io_s),
    .io_co(HalfAdder_86_io_co)
  );
  FullAdder FullAdder_2770 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2770_io_a),
    .io_b(FullAdder_2770_io_b),
    .io_ci(FullAdder_2770_io_ci),
    .io_s(FullAdder_2770_io_s),
    .io_co(FullAdder_2770_io_co)
  );
  FullAdder FullAdder_2771 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2771_io_a),
    .io_b(FullAdder_2771_io_b),
    .io_ci(FullAdder_2771_io_ci),
    .io_s(FullAdder_2771_io_s),
    .io_co(FullAdder_2771_io_co)
  );
  FullAdder FullAdder_2772 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2772_io_a),
    .io_b(FullAdder_2772_io_b),
    .io_ci(FullAdder_2772_io_ci),
    .io_s(FullAdder_2772_io_s),
    .io_co(FullAdder_2772_io_co)
  );
  FullAdder FullAdder_2773 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2773_io_a),
    .io_b(FullAdder_2773_io_b),
    .io_ci(FullAdder_2773_io_ci),
    .io_s(FullAdder_2773_io_s),
    .io_co(FullAdder_2773_io_co)
  );
  FullAdder FullAdder_2774 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2774_io_a),
    .io_b(FullAdder_2774_io_b),
    .io_ci(FullAdder_2774_io_ci),
    .io_s(FullAdder_2774_io_s),
    .io_co(FullAdder_2774_io_co)
  );
  FullAdder FullAdder_2775 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2775_io_a),
    .io_b(FullAdder_2775_io_b),
    .io_ci(FullAdder_2775_io_ci),
    .io_s(FullAdder_2775_io_s),
    .io_co(FullAdder_2775_io_co)
  );
  FullAdder FullAdder_2776 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2776_io_a),
    .io_b(FullAdder_2776_io_b),
    .io_ci(FullAdder_2776_io_ci),
    .io_s(FullAdder_2776_io_s),
    .io_co(FullAdder_2776_io_co)
  );
  FullAdder FullAdder_2777 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2777_io_a),
    .io_b(FullAdder_2777_io_b),
    .io_ci(FullAdder_2777_io_ci),
    .io_s(FullAdder_2777_io_s),
    .io_co(FullAdder_2777_io_co)
  );
  FullAdder FullAdder_2778 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2778_io_a),
    .io_b(FullAdder_2778_io_b),
    .io_ci(FullAdder_2778_io_ci),
    .io_s(FullAdder_2778_io_s),
    .io_co(FullAdder_2778_io_co)
  );
  HalfAdder HalfAdder_87 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_87_io_a),
    .io_b(HalfAdder_87_io_b),
    .io_s(HalfAdder_87_io_s),
    .io_co(HalfAdder_87_io_co)
  );
  HalfAdder HalfAdder_88 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_88_io_a),
    .io_b(HalfAdder_88_io_b),
    .io_s(HalfAdder_88_io_s),
    .io_co(HalfAdder_88_io_co)
  );
  FullAdder FullAdder_2779 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2779_io_a),
    .io_b(FullAdder_2779_io_b),
    .io_ci(FullAdder_2779_io_ci),
    .io_s(FullAdder_2779_io_s),
    .io_co(FullAdder_2779_io_co)
  );
  HalfAdder HalfAdder_89 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_89_io_a),
    .io_b(HalfAdder_89_io_b),
    .io_s(HalfAdder_89_io_s),
    .io_co(HalfAdder_89_io_co)
  );
  FullAdder FullAdder_2780 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2780_io_a),
    .io_b(FullAdder_2780_io_b),
    .io_ci(FullAdder_2780_io_ci),
    .io_s(FullAdder_2780_io_s),
    .io_co(FullAdder_2780_io_co)
  );
  FullAdder FullAdder_2781 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2781_io_a),
    .io_b(FullAdder_2781_io_b),
    .io_ci(FullAdder_2781_io_ci),
    .io_s(FullAdder_2781_io_s),
    .io_co(FullAdder_2781_io_co)
  );
  FullAdder FullAdder_2782 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2782_io_a),
    .io_b(FullAdder_2782_io_b),
    .io_ci(FullAdder_2782_io_ci),
    .io_s(FullAdder_2782_io_s),
    .io_co(FullAdder_2782_io_co)
  );
  FullAdder FullAdder_2783 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2783_io_a),
    .io_b(FullAdder_2783_io_b),
    .io_ci(FullAdder_2783_io_ci),
    .io_s(FullAdder_2783_io_s),
    .io_co(FullAdder_2783_io_co)
  );
  HalfAdder HalfAdder_90 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_90_io_a),
    .io_b(HalfAdder_90_io_b),
    .io_s(HalfAdder_90_io_s),
    .io_co(HalfAdder_90_io_co)
  );
  HalfAdder HalfAdder_91 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_91_io_a),
    .io_b(HalfAdder_91_io_b),
    .io_s(HalfAdder_91_io_s),
    .io_co(HalfAdder_91_io_co)
  );
  HalfAdder HalfAdder_92 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_92_io_a),
    .io_b(HalfAdder_92_io_b),
    .io_s(HalfAdder_92_io_s),
    .io_co(HalfAdder_92_io_co)
  );
  HalfAdder HalfAdder_93 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_93_io_a),
    .io_b(HalfAdder_93_io_b),
    .io_s(HalfAdder_93_io_s),
    .io_co(HalfAdder_93_io_co)
  );
  HalfAdder HalfAdder_94 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_94_io_a),
    .io_b(HalfAdder_94_io_b),
    .io_s(HalfAdder_94_io_s),
    .io_co(HalfAdder_94_io_co)
  );
  HalfAdder HalfAdder_95 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_95_io_a),
    .io_b(HalfAdder_95_io_b),
    .io_s(HalfAdder_95_io_s),
    .io_co(HalfAdder_95_io_co)
  );
  FullAdder FullAdder_2784 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2784_io_a),
    .io_b(FullAdder_2784_io_b),
    .io_ci(FullAdder_2784_io_ci),
    .io_s(FullAdder_2784_io_s),
    .io_co(FullAdder_2784_io_co)
  );
  HalfAdder HalfAdder_96 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_96_io_a),
    .io_b(HalfAdder_96_io_b),
    .io_s(HalfAdder_96_io_s),
    .io_co(HalfAdder_96_io_co)
  );
  FullAdder FullAdder_2785 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2785_io_a),
    .io_b(FullAdder_2785_io_b),
    .io_ci(FullAdder_2785_io_ci),
    .io_s(FullAdder_2785_io_s),
    .io_co(FullAdder_2785_io_co)
  );
  FullAdder FullAdder_2786 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2786_io_a),
    .io_b(FullAdder_2786_io_b),
    .io_ci(FullAdder_2786_io_ci),
    .io_s(FullAdder_2786_io_s),
    .io_co(FullAdder_2786_io_co)
  );
  FullAdder FullAdder_2787 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2787_io_a),
    .io_b(FullAdder_2787_io_b),
    .io_ci(FullAdder_2787_io_ci),
    .io_s(FullAdder_2787_io_s),
    .io_co(FullAdder_2787_io_co)
  );
  FullAdder FullAdder_2788 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2788_io_a),
    .io_b(FullAdder_2788_io_b),
    .io_ci(FullAdder_2788_io_ci),
    .io_s(FullAdder_2788_io_s),
    .io_co(FullAdder_2788_io_co)
  );
  FullAdder FullAdder_2789 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2789_io_a),
    .io_b(FullAdder_2789_io_b),
    .io_ci(FullAdder_2789_io_ci),
    .io_s(FullAdder_2789_io_s),
    .io_co(FullAdder_2789_io_co)
  );
  FullAdder FullAdder_2790 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2790_io_a),
    .io_b(FullAdder_2790_io_b),
    .io_ci(FullAdder_2790_io_ci),
    .io_s(FullAdder_2790_io_s),
    .io_co(FullAdder_2790_io_co)
  );
  FullAdder FullAdder_2791 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2791_io_a),
    .io_b(FullAdder_2791_io_b),
    .io_ci(FullAdder_2791_io_ci),
    .io_s(FullAdder_2791_io_s),
    .io_co(FullAdder_2791_io_co)
  );
  FullAdder FullAdder_2792 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2792_io_a),
    .io_b(FullAdder_2792_io_b),
    .io_ci(FullAdder_2792_io_ci),
    .io_s(FullAdder_2792_io_s),
    .io_co(FullAdder_2792_io_co)
  );
  FullAdder FullAdder_2793 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2793_io_a),
    .io_b(FullAdder_2793_io_b),
    .io_ci(FullAdder_2793_io_ci),
    .io_s(FullAdder_2793_io_s),
    .io_co(FullAdder_2793_io_co)
  );
  FullAdder FullAdder_2794 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2794_io_a),
    .io_b(FullAdder_2794_io_b),
    .io_ci(FullAdder_2794_io_ci),
    .io_s(FullAdder_2794_io_s),
    .io_co(FullAdder_2794_io_co)
  );
  FullAdder FullAdder_2795 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2795_io_a),
    .io_b(FullAdder_2795_io_b),
    .io_ci(FullAdder_2795_io_ci),
    .io_s(FullAdder_2795_io_s),
    .io_co(FullAdder_2795_io_co)
  );
  FullAdder FullAdder_2796 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2796_io_a),
    .io_b(FullAdder_2796_io_b),
    .io_ci(FullAdder_2796_io_ci),
    .io_s(FullAdder_2796_io_s),
    .io_co(FullAdder_2796_io_co)
  );
  FullAdder FullAdder_2797 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2797_io_a),
    .io_b(FullAdder_2797_io_b),
    .io_ci(FullAdder_2797_io_ci),
    .io_s(FullAdder_2797_io_s),
    .io_co(FullAdder_2797_io_co)
  );
  FullAdder FullAdder_2798 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2798_io_a),
    .io_b(FullAdder_2798_io_b),
    .io_ci(FullAdder_2798_io_ci),
    .io_s(FullAdder_2798_io_s),
    .io_co(FullAdder_2798_io_co)
  );
  FullAdder FullAdder_2799 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2799_io_a),
    .io_b(FullAdder_2799_io_b),
    .io_ci(FullAdder_2799_io_ci),
    .io_s(FullAdder_2799_io_s),
    .io_co(FullAdder_2799_io_co)
  );
  FullAdder FullAdder_2800 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2800_io_a),
    .io_b(FullAdder_2800_io_b),
    .io_ci(FullAdder_2800_io_ci),
    .io_s(FullAdder_2800_io_s),
    .io_co(FullAdder_2800_io_co)
  );
  FullAdder FullAdder_2801 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2801_io_a),
    .io_b(FullAdder_2801_io_b),
    .io_ci(FullAdder_2801_io_ci),
    .io_s(FullAdder_2801_io_s),
    .io_co(FullAdder_2801_io_co)
  );
  FullAdder FullAdder_2802 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2802_io_a),
    .io_b(FullAdder_2802_io_b),
    .io_ci(FullAdder_2802_io_ci),
    .io_s(FullAdder_2802_io_s),
    .io_co(FullAdder_2802_io_co)
  );
  FullAdder FullAdder_2803 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2803_io_a),
    .io_b(FullAdder_2803_io_b),
    .io_ci(FullAdder_2803_io_ci),
    .io_s(FullAdder_2803_io_s),
    .io_co(FullAdder_2803_io_co)
  );
  FullAdder FullAdder_2804 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2804_io_a),
    .io_b(FullAdder_2804_io_b),
    .io_ci(FullAdder_2804_io_ci),
    .io_s(FullAdder_2804_io_s),
    .io_co(FullAdder_2804_io_co)
  );
  FullAdder FullAdder_2805 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2805_io_a),
    .io_b(FullAdder_2805_io_b),
    .io_ci(FullAdder_2805_io_ci),
    .io_s(FullAdder_2805_io_s),
    .io_co(FullAdder_2805_io_co)
  );
  FullAdder FullAdder_2806 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2806_io_a),
    .io_b(FullAdder_2806_io_b),
    .io_ci(FullAdder_2806_io_ci),
    .io_s(FullAdder_2806_io_s),
    .io_co(FullAdder_2806_io_co)
  );
  FullAdder FullAdder_2807 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2807_io_a),
    .io_b(FullAdder_2807_io_b),
    .io_ci(FullAdder_2807_io_ci),
    .io_s(FullAdder_2807_io_s),
    .io_co(FullAdder_2807_io_co)
  );
  FullAdder FullAdder_2808 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2808_io_a),
    .io_b(FullAdder_2808_io_b),
    .io_ci(FullAdder_2808_io_ci),
    .io_s(FullAdder_2808_io_s),
    .io_co(FullAdder_2808_io_co)
  );
  FullAdder FullAdder_2809 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2809_io_a),
    .io_b(FullAdder_2809_io_b),
    .io_ci(FullAdder_2809_io_ci),
    .io_s(FullAdder_2809_io_s),
    .io_co(FullAdder_2809_io_co)
  );
  FullAdder FullAdder_2810 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2810_io_a),
    .io_b(FullAdder_2810_io_b),
    .io_ci(FullAdder_2810_io_ci),
    .io_s(FullAdder_2810_io_s),
    .io_co(FullAdder_2810_io_co)
  );
  FullAdder FullAdder_2811 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2811_io_a),
    .io_b(FullAdder_2811_io_b),
    .io_ci(FullAdder_2811_io_ci),
    .io_s(FullAdder_2811_io_s),
    .io_co(FullAdder_2811_io_co)
  );
  FullAdder FullAdder_2812 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2812_io_a),
    .io_b(FullAdder_2812_io_b),
    .io_ci(FullAdder_2812_io_ci),
    .io_s(FullAdder_2812_io_s),
    .io_co(FullAdder_2812_io_co)
  );
  FullAdder FullAdder_2813 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2813_io_a),
    .io_b(FullAdder_2813_io_b),
    .io_ci(FullAdder_2813_io_ci),
    .io_s(FullAdder_2813_io_s),
    .io_co(FullAdder_2813_io_co)
  );
  FullAdder FullAdder_2814 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2814_io_a),
    .io_b(FullAdder_2814_io_b),
    .io_ci(FullAdder_2814_io_ci),
    .io_s(FullAdder_2814_io_s),
    .io_co(FullAdder_2814_io_co)
  );
  FullAdder FullAdder_2815 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2815_io_a),
    .io_b(FullAdder_2815_io_b),
    .io_ci(FullAdder_2815_io_ci),
    .io_s(FullAdder_2815_io_s),
    .io_co(FullAdder_2815_io_co)
  );
  FullAdder FullAdder_2816 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2816_io_a),
    .io_b(FullAdder_2816_io_b),
    .io_ci(FullAdder_2816_io_ci),
    .io_s(FullAdder_2816_io_s),
    .io_co(FullAdder_2816_io_co)
  );
  FullAdder FullAdder_2817 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2817_io_a),
    .io_b(FullAdder_2817_io_b),
    .io_ci(FullAdder_2817_io_ci),
    .io_s(FullAdder_2817_io_s),
    .io_co(FullAdder_2817_io_co)
  );
  FullAdder FullAdder_2818 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2818_io_a),
    .io_b(FullAdder_2818_io_b),
    .io_ci(FullAdder_2818_io_ci),
    .io_s(FullAdder_2818_io_s),
    .io_co(FullAdder_2818_io_co)
  );
  FullAdder FullAdder_2819 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2819_io_a),
    .io_b(FullAdder_2819_io_b),
    .io_ci(FullAdder_2819_io_ci),
    .io_s(FullAdder_2819_io_s),
    .io_co(FullAdder_2819_io_co)
  );
  FullAdder FullAdder_2820 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2820_io_a),
    .io_b(FullAdder_2820_io_b),
    .io_ci(FullAdder_2820_io_ci),
    .io_s(FullAdder_2820_io_s),
    .io_co(FullAdder_2820_io_co)
  );
  FullAdder FullAdder_2821 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2821_io_a),
    .io_b(FullAdder_2821_io_b),
    .io_ci(FullAdder_2821_io_ci),
    .io_s(FullAdder_2821_io_s),
    .io_co(FullAdder_2821_io_co)
  );
  HalfAdder HalfAdder_97 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_97_io_a),
    .io_b(HalfAdder_97_io_b),
    .io_s(HalfAdder_97_io_s),
    .io_co(HalfAdder_97_io_co)
  );
  FullAdder FullAdder_2822 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2822_io_a),
    .io_b(FullAdder_2822_io_b),
    .io_ci(FullAdder_2822_io_ci),
    .io_s(FullAdder_2822_io_s),
    .io_co(FullAdder_2822_io_co)
  );
  FullAdder FullAdder_2823 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2823_io_a),
    .io_b(FullAdder_2823_io_b),
    .io_ci(FullAdder_2823_io_ci),
    .io_s(FullAdder_2823_io_s),
    .io_co(FullAdder_2823_io_co)
  );
  FullAdder FullAdder_2824 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2824_io_a),
    .io_b(FullAdder_2824_io_b),
    .io_ci(FullAdder_2824_io_ci),
    .io_s(FullAdder_2824_io_s),
    .io_co(FullAdder_2824_io_co)
  );
  FullAdder FullAdder_2825 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2825_io_a),
    .io_b(FullAdder_2825_io_b),
    .io_ci(FullAdder_2825_io_ci),
    .io_s(FullAdder_2825_io_s),
    .io_co(FullAdder_2825_io_co)
  );
  FullAdder FullAdder_2826 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2826_io_a),
    .io_b(FullAdder_2826_io_b),
    .io_ci(FullAdder_2826_io_ci),
    .io_s(FullAdder_2826_io_s),
    .io_co(FullAdder_2826_io_co)
  );
  FullAdder FullAdder_2827 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2827_io_a),
    .io_b(FullAdder_2827_io_b),
    .io_ci(FullAdder_2827_io_ci),
    .io_s(FullAdder_2827_io_s),
    .io_co(FullAdder_2827_io_co)
  );
  FullAdder FullAdder_2828 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2828_io_a),
    .io_b(FullAdder_2828_io_b),
    .io_ci(FullAdder_2828_io_ci),
    .io_s(FullAdder_2828_io_s),
    .io_co(FullAdder_2828_io_co)
  );
  FullAdder FullAdder_2829 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2829_io_a),
    .io_b(FullAdder_2829_io_b),
    .io_ci(FullAdder_2829_io_ci),
    .io_s(FullAdder_2829_io_s),
    .io_co(FullAdder_2829_io_co)
  );
  FullAdder FullAdder_2830 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2830_io_a),
    .io_b(FullAdder_2830_io_b),
    .io_ci(FullAdder_2830_io_ci),
    .io_s(FullAdder_2830_io_s),
    .io_co(FullAdder_2830_io_co)
  );
  FullAdder FullAdder_2831 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2831_io_a),
    .io_b(FullAdder_2831_io_b),
    .io_ci(FullAdder_2831_io_ci),
    .io_s(FullAdder_2831_io_s),
    .io_co(FullAdder_2831_io_co)
  );
  FullAdder FullAdder_2832 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2832_io_a),
    .io_b(FullAdder_2832_io_b),
    .io_ci(FullAdder_2832_io_ci),
    .io_s(FullAdder_2832_io_s),
    .io_co(FullAdder_2832_io_co)
  );
  FullAdder FullAdder_2833 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2833_io_a),
    .io_b(FullAdder_2833_io_b),
    .io_ci(FullAdder_2833_io_ci),
    .io_s(FullAdder_2833_io_s),
    .io_co(FullAdder_2833_io_co)
  );
  FullAdder FullAdder_2834 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2834_io_a),
    .io_b(FullAdder_2834_io_b),
    .io_ci(FullAdder_2834_io_ci),
    .io_s(FullAdder_2834_io_s),
    .io_co(FullAdder_2834_io_co)
  );
  FullAdder FullAdder_2835 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2835_io_a),
    .io_b(FullAdder_2835_io_b),
    .io_ci(FullAdder_2835_io_ci),
    .io_s(FullAdder_2835_io_s),
    .io_co(FullAdder_2835_io_co)
  );
  FullAdder FullAdder_2836 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2836_io_a),
    .io_b(FullAdder_2836_io_b),
    .io_ci(FullAdder_2836_io_ci),
    .io_s(FullAdder_2836_io_s),
    .io_co(FullAdder_2836_io_co)
  );
  FullAdder FullAdder_2837 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2837_io_a),
    .io_b(FullAdder_2837_io_b),
    .io_ci(FullAdder_2837_io_ci),
    .io_s(FullAdder_2837_io_s),
    .io_co(FullAdder_2837_io_co)
  );
  FullAdder FullAdder_2838 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2838_io_a),
    .io_b(FullAdder_2838_io_b),
    .io_ci(FullAdder_2838_io_ci),
    .io_s(FullAdder_2838_io_s),
    .io_co(FullAdder_2838_io_co)
  );
  FullAdder FullAdder_2839 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2839_io_a),
    .io_b(FullAdder_2839_io_b),
    .io_ci(FullAdder_2839_io_ci),
    .io_s(FullAdder_2839_io_s),
    .io_co(FullAdder_2839_io_co)
  );
  HalfAdder HalfAdder_98 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_98_io_a),
    .io_b(HalfAdder_98_io_b),
    .io_s(HalfAdder_98_io_s),
    .io_co(HalfAdder_98_io_co)
  );
  FullAdder FullAdder_2840 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2840_io_a),
    .io_b(FullAdder_2840_io_b),
    .io_ci(FullAdder_2840_io_ci),
    .io_s(FullAdder_2840_io_s),
    .io_co(FullAdder_2840_io_co)
  );
  FullAdder FullAdder_2841 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2841_io_a),
    .io_b(FullAdder_2841_io_b),
    .io_ci(FullAdder_2841_io_ci),
    .io_s(FullAdder_2841_io_s),
    .io_co(FullAdder_2841_io_co)
  );
  FullAdder FullAdder_2842 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2842_io_a),
    .io_b(FullAdder_2842_io_b),
    .io_ci(FullAdder_2842_io_ci),
    .io_s(FullAdder_2842_io_s),
    .io_co(FullAdder_2842_io_co)
  );
  HalfAdder HalfAdder_99 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_99_io_a),
    .io_b(HalfAdder_99_io_b),
    .io_s(HalfAdder_99_io_s),
    .io_co(HalfAdder_99_io_co)
  );
  FullAdder FullAdder_2843 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2843_io_a),
    .io_b(FullAdder_2843_io_b),
    .io_ci(FullAdder_2843_io_ci),
    .io_s(FullAdder_2843_io_s),
    .io_co(FullAdder_2843_io_co)
  );
  FullAdder FullAdder_2844 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2844_io_a),
    .io_b(FullAdder_2844_io_b),
    .io_ci(FullAdder_2844_io_ci),
    .io_s(FullAdder_2844_io_s),
    .io_co(FullAdder_2844_io_co)
  );
  FullAdder FullAdder_2845 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2845_io_a),
    .io_b(FullAdder_2845_io_b),
    .io_ci(FullAdder_2845_io_ci),
    .io_s(FullAdder_2845_io_s),
    .io_co(FullAdder_2845_io_co)
  );
  HalfAdder HalfAdder_100 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_100_io_a),
    .io_b(HalfAdder_100_io_b),
    .io_s(HalfAdder_100_io_s),
    .io_co(HalfAdder_100_io_co)
  );
  FullAdder FullAdder_2846 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2846_io_a),
    .io_b(FullAdder_2846_io_b),
    .io_ci(FullAdder_2846_io_ci),
    .io_s(FullAdder_2846_io_s),
    .io_co(FullAdder_2846_io_co)
  );
  FullAdder FullAdder_2847 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2847_io_a),
    .io_b(FullAdder_2847_io_b),
    .io_ci(FullAdder_2847_io_ci),
    .io_s(FullAdder_2847_io_s),
    .io_co(FullAdder_2847_io_co)
  );
  FullAdder FullAdder_2848 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2848_io_a),
    .io_b(FullAdder_2848_io_b),
    .io_ci(FullAdder_2848_io_ci),
    .io_s(FullAdder_2848_io_s),
    .io_co(FullAdder_2848_io_co)
  );
  FullAdder FullAdder_2849 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2849_io_a),
    .io_b(FullAdder_2849_io_b),
    .io_ci(FullAdder_2849_io_ci),
    .io_s(FullAdder_2849_io_s),
    .io_co(FullAdder_2849_io_co)
  );
  FullAdder FullAdder_2850 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2850_io_a),
    .io_b(FullAdder_2850_io_b),
    .io_ci(FullAdder_2850_io_ci),
    .io_s(FullAdder_2850_io_s),
    .io_co(FullAdder_2850_io_co)
  );
  FullAdder FullAdder_2851 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2851_io_a),
    .io_b(FullAdder_2851_io_b),
    .io_ci(FullAdder_2851_io_ci),
    .io_s(FullAdder_2851_io_s),
    .io_co(FullAdder_2851_io_co)
  );
  FullAdder FullAdder_2852 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2852_io_a),
    .io_b(FullAdder_2852_io_b),
    .io_ci(FullAdder_2852_io_ci),
    .io_s(FullAdder_2852_io_s),
    .io_co(FullAdder_2852_io_co)
  );
  FullAdder FullAdder_2853 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2853_io_a),
    .io_b(FullAdder_2853_io_b),
    .io_ci(FullAdder_2853_io_ci),
    .io_s(FullAdder_2853_io_s),
    .io_co(FullAdder_2853_io_co)
  );
  FullAdder FullAdder_2854 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2854_io_a),
    .io_b(FullAdder_2854_io_b),
    .io_ci(FullAdder_2854_io_ci),
    .io_s(FullAdder_2854_io_s),
    .io_co(FullAdder_2854_io_co)
  );
  FullAdder FullAdder_2855 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2855_io_a),
    .io_b(FullAdder_2855_io_b),
    .io_ci(FullAdder_2855_io_ci),
    .io_s(FullAdder_2855_io_s),
    .io_co(FullAdder_2855_io_co)
  );
  FullAdder FullAdder_2856 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2856_io_a),
    .io_b(FullAdder_2856_io_b),
    .io_ci(FullAdder_2856_io_ci),
    .io_s(FullAdder_2856_io_s),
    .io_co(FullAdder_2856_io_co)
  );
  FullAdder FullAdder_2857 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2857_io_a),
    .io_b(FullAdder_2857_io_b),
    .io_ci(FullAdder_2857_io_ci),
    .io_s(FullAdder_2857_io_s),
    .io_co(FullAdder_2857_io_co)
  );
  FullAdder FullAdder_2858 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2858_io_a),
    .io_b(FullAdder_2858_io_b),
    .io_ci(FullAdder_2858_io_ci),
    .io_s(FullAdder_2858_io_s),
    .io_co(FullAdder_2858_io_co)
  );
  FullAdder FullAdder_2859 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2859_io_a),
    .io_b(FullAdder_2859_io_b),
    .io_ci(FullAdder_2859_io_ci),
    .io_s(FullAdder_2859_io_s),
    .io_co(FullAdder_2859_io_co)
  );
  FullAdder FullAdder_2860 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2860_io_a),
    .io_b(FullAdder_2860_io_b),
    .io_ci(FullAdder_2860_io_ci),
    .io_s(FullAdder_2860_io_s),
    .io_co(FullAdder_2860_io_co)
  );
  FullAdder FullAdder_2861 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2861_io_a),
    .io_b(FullAdder_2861_io_b),
    .io_ci(FullAdder_2861_io_ci),
    .io_s(FullAdder_2861_io_s),
    .io_co(FullAdder_2861_io_co)
  );
  FullAdder FullAdder_2862 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2862_io_a),
    .io_b(FullAdder_2862_io_b),
    .io_ci(FullAdder_2862_io_ci),
    .io_s(FullAdder_2862_io_s),
    .io_co(FullAdder_2862_io_co)
  );
  FullAdder FullAdder_2863 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2863_io_a),
    .io_b(FullAdder_2863_io_b),
    .io_ci(FullAdder_2863_io_ci),
    .io_s(FullAdder_2863_io_s),
    .io_co(FullAdder_2863_io_co)
  );
  FullAdder FullAdder_2864 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2864_io_a),
    .io_b(FullAdder_2864_io_b),
    .io_ci(FullAdder_2864_io_ci),
    .io_s(FullAdder_2864_io_s),
    .io_co(FullAdder_2864_io_co)
  );
  FullAdder FullAdder_2865 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2865_io_a),
    .io_b(FullAdder_2865_io_b),
    .io_ci(FullAdder_2865_io_ci),
    .io_s(FullAdder_2865_io_s),
    .io_co(FullAdder_2865_io_co)
  );
  FullAdder FullAdder_2866 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2866_io_a),
    .io_b(FullAdder_2866_io_b),
    .io_ci(FullAdder_2866_io_ci),
    .io_s(FullAdder_2866_io_s),
    .io_co(FullAdder_2866_io_co)
  );
  FullAdder FullAdder_2867 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2867_io_a),
    .io_b(FullAdder_2867_io_b),
    .io_ci(FullAdder_2867_io_ci),
    .io_s(FullAdder_2867_io_s),
    .io_co(FullAdder_2867_io_co)
  );
  FullAdder FullAdder_2868 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2868_io_a),
    .io_b(FullAdder_2868_io_b),
    .io_ci(FullAdder_2868_io_ci),
    .io_s(FullAdder_2868_io_s),
    .io_co(FullAdder_2868_io_co)
  );
  FullAdder FullAdder_2869 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2869_io_a),
    .io_b(FullAdder_2869_io_b),
    .io_ci(FullAdder_2869_io_ci),
    .io_s(FullAdder_2869_io_s),
    .io_co(FullAdder_2869_io_co)
  );
  FullAdder FullAdder_2870 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2870_io_a),
    .io_b(FullAdder_2870_io_b),
    .io_ci(FullAdder_2870_io_ci),
    .io_s(FullAdder_2870_io_s),
    .io_co(FullAdder_2870_io_co)
  );
  FullAdder FullAdder_2871 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2871_io_a),
    .io_b(FullAdder_2871_io_b),
    .io_ci(FullAdder_2871_io_ci),
    .io_s(FullAdder_2871_io_s),
    .io_co(FullAdder_2871_io_co)
  );
  FullAdder FullAdder_2872 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2872_io_a),
    .io_b(FullAdder_2872_io_b),
    .io_ci(FullAdder_2872_io_ci),
    .io_s(FullAdder_2872_io_s),
    .io_co(FullAdder_2872_io_co)
  );
  FullAdder FullAdder_2873 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2873_io_a),
    .io_b(FullAdder_2873_io_b),
    .io_ci(FullAdder_2873_io_ci),
    .io_s(FullAdder_2873_io_s),
    .io_co(FullAdder_2873_io_co)
  );
  FullAdder FullAdder_2874 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2874_io_a),
    .io_b(FullAdder_2874_io_b),
    .io_ci(FullAdder_2874_io_ci),
    .io_s(FullAdder_2874_io_s),
    .io_co(FullAdder_2874_io_co)
  );
  FullAdder FullAdder_2875 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2875_io_a),
    .io_b(FullAdder_2875_io_b),
    .io_ci(FullAdder_2875_io_ci),
    .io_s(FullAdder_2875_io_s),
    .io_co(FullAdder_2875_io_co)
  );
  FullAdder FullAdder_2876 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2876_io_a),
    .io_b(FullAdder_2876_io_b),
    .io_ci(FullAdder_2876_io_ci),
    .io_s(FullAdder_2876_io_s),
    .io_co(FullAdder_2876_io_co)
  );
  FullAdder FullAdder_2877 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2877_io_a),
    .io_b(FullAdder_2877_io_b),
    .io_ci(FullAdder_2877_io_ci),
    .io_s(FullAdder_2877_io_s),
    .io_co(FullAdder_2877_io_co)
  );
  FullAdder FullAdder_2878 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2878_io_a),
    .io_b(FullAdder_2878_io_b),
    .io_ci(FullAdder_2878_io_ci),
    .io_s(FullAdder_2878_io_s),
    .io_co(FullAdder_2878_io_co)
  );
  HalfAdder HalfAdder_101 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_101_io_a),
    .io_b(HalfAdder_101_io_b),
    .io_s(HalfAdder_101_io_s),
    .io_co(HalfAdder_101_io_co)
  );
  FullAdder FullAdder_2879 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2879_io_a),
    .io_b(FullAdder_2879_io_b),
    .io_ci(FullAdder_2879_io_ci),
    .io_s(FullAdder_2879_io_s),
    .io_co(FullAdder_2879_io_co)
  );
  FullAdder FullAdder_2880 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2880_io_a),
    .io_b(FullAdder_2880_io_b),
    .io_ci(FullAdder_2880_io_ci),
    .io_s(FullAdder_2880_io_s),
    .io_co(FullAdder_2880_io_co)
  );
  FullAdder FullAdder_2881 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2881_io_a),
    .io_b(FullAdder_2881_io_b),
    .io_ci(FullAdder_2881_io_ci),
    .io_s(FullAdder_2881_io_s),
    .io_co(FullAdder_2881_io_co)
  );
  FullAdder FullAdder_2882 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2882_io_a),
    .io_b(FullAdder_2882_io_b),
    .io_ci(FullAdder_2882_io_ci),
    .io_s(FullAdder_2882_io_s),
    .io_co(FullAdder_2882_io_co)
  );
  FullAdder FullAdder_2883 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2883_io_a),
    .io_b(FullAdder_2883_io_b),
    .io_ci(FullAdder_2883_io_ci),
    .io_s(FullAdder_2883_io_s),
    .io_co(FullAdder_2883_io_co)
  );
  FullAdder FullAdder_2884 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2884_io_a),
    .io_b(FullAdder_2884_io_b),
    .io_ci(FullAdder_2884_io_ci),
    .io_s(FullAdder_2884_io_s),
    .io_co(FullAdder_2884_io_co)
  );
  FullAdder FullAdder_2885 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2885_io_a),
    .io_b(FullAdder_2885_io_b),
    .io_ci(FullAdder_2885_io_ci),
    .io_s(FullAdder_2885_io_s),
    .io_co(FullAdder_2885_io_co)
  );
  FullAdder FullAdder_2886 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2886_io_a),
    .io_b(FullAdder_2886_io_b),
    .io_ci(FullAdder_2886_io_ci),
    .io_s(FullAdder_2886_io_s),
    .io_co(FullAdder_2886_io_co)
  );
  FullAdder FullAdder_2887 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2887_io_a),
    .io_b(FullAdder_2887_io_b),
    .io_ci(FullAdder_2887_io_ci),
    .io_s(FullAdder_2887_io_s),
    .io_co(FullAdder_2887_io_co)
  );
  FullAdder FullAdder_2888 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2888_io_a),
    .io_b(FullAdder_2888_io_b),
    .io_ci(FullAdder_2888_io_ci),
    .io_s(FullAdder_2888_io_s),
    .io_co(FullAdder_2888_io_co)
  );
  FullAdder FullAdder_2889 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2889_io_a),
    .io_b(FullAdder_2889_io_b),
    .io_ci(FullAdder_2889_io_ci),
    .io_s(FullAdder_2889_io_s),
    .io_co(FullAdder_2889_io_co)
  );
  FullAdder FullAdder_2890 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2890_io_a),
    .io_b(FullAdder_2890_io_b),
    .io_ci(FullAdder_2890_io_ci),
    .io_s(FullAdder_2890_io_s),
    .io_co(FullAdder_2890_io_co)
  );
  FullAdder FullAdder_2891 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2891_io_a),
    .io_b(FullAdder_2891_io_b),
    .io_ci(FullAdder_2891_io_ci),
    .io_s(FullAdder_2891_io_s),
    .io_co(FullAdder_2891_io_co)
  );
  FullAdder FullAdder_2892 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2892_io_a),
    .io_b(FullAdder_2892_io_b),
    .io_ci(FullAdder_2892_io_ci),
    .io_s(FullAdder_2892_io_s),
    .io_co(FullAdder_2892_io_co)
  );
  FullAdder FullAdder_2893 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2893_io_a),
    .io_b(FullAdder_2893_io_b),
    .io_ci(FullAdder_2893_io_ci),
    .io_s(FullAdder_2893_io_s),
    .io_co(FullAdder_2893_io_co)
  );
  FullAdder FullAdder_2894 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2894_io_a),
    .io_b(FullAdder_2894_io_b),
    .io_ci(FullAdder_2894_io_ci),
    .io_s(FullAdder_2894_io_s),
    .io_co(FullAdder_2894_io_co)
  );
  FullAdder FullAdder_2895 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2895_io_a),
    .io_b(FullAdder_2895_io_b),
    .io_ci(FullAdder_2895_io_ci),
    .io_s(FullAdder_2895_io_s),
    .io_co(FullAdder_2895_io_co)
  );
  FullAdder FullAdder_2896 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2896_io_a),
    .io_b(FullAdder_2896_io_b),
    .io_ci(FullAdder_2896_io_ci),
    .io_s(FullAdder_2896_io_s),
    .io_co(FullAdder_2896_io_co)
  );
  FullAdder FullAdder_2897 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2897_io_a),
    .io_b(FullAdder_2897_io_b),
    .io_ci(FullAdder_2897_io_ci),
    .io_s(FullAdder_2897_io_s),
    .io_co(FullAdder_2897_io_co)
  );
  FullAdder FullAdder_2898 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2898_io_a),
    .io_b(FullAdder_2898_io_b),
    .io_ci(FullAdder_2898_io_ci),
    .io_s(FullAdder_2898_io_s),
    .io_co(FullAdder_2898_io_co)
  );
  FullAdder FullAdder_2899 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2899_io_a),
    .io_b(FullAdder_2899_io_b),
    .io_ci(FullAdder_2899_io_ci),
    .io_s(FullAdder_2899_io_s),
    .io_co(FullAdder_2899_io_co)
  );
  FullAdder FullAdder_2900 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2900_io_a),
    .io_b(FullAdder_2900_io_b),
    .io_ci(FullAdder_2900_io_ci),
    .io_s(FullAdder_2900_io_s),
    .io_co(FullAdder_2900_io_co)
  );
  FullAdder FullAdder_2901 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2901_io_a),
    .io_b(FullAdder_2901_io_b),
    .io_ci(FullAdder_2901_io_ci),
    .io_s(FullAdder_2901_io_s),
    .io_co(FullAdder_2901_io_co)
  );
  FullAdder FullAdder_2902 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2902_io_a),
    .io_b(FullAdder_2902_io_b),
    .io_ci(FullAdder_2902_io_ci),
    .io_s(FullAdder_2902_io_s),
    .io_co(FullAdder_2902_io_co)
  );
  FullAdder FullAdder_2903 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2903_io_a),
    .io_b(FullAdder_2903_io_b),
    .io_ci(FullAdder_2903_io_ci),
    .io_s(FullAdder_2903_io_s),
    .io_co(FullAdder_2903_io_co)
  );
  FullAdder FullAdder_2904 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2904_io_a),
    .io_b(FullAdder_2904_io_b),
    .io_ci(FullAdder_2904_io_ci),
    .io_s(FullAdder_2904_io_s),
    .io_co(FullAdder_2904_io_co)
  );
  FullAdder FullAdder_2905 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2905_io_a),
    .io_b(FullAdder_2905_io_b),
    .io_ci(FullAdder_2905_io_ci),
    .io_s(FullAdder_2905_io_s),
    .io_co(FullAdder_2905_io_co)
  );
  FullAdder FullAdder_2906 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2906_io_a),
    .io_b(FullAdder_2906_io_b),
    .io_ci(FullAdder_2906_io_ci),
    .io_s(FullAdder_2906_io_s),
    .io_co(FullAdder_2906_io_co)
  );
  FullAdder FullAdder_2907 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2907_io_a),
    .io_b(FullAdder_2907_io_b),
    .io_ci(FullAdder_2907_io_ci),
    .io_s(FullAdder_2907_io_s),
    .io_co(FullAdder_2907_io_co)
  );
  FullAdder FullAdder_2908 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2908_io_a),
    .io_b(FullAdder_2908_io_b),
    .io_ci(FullAdder_2908_io_ci),
    .io_s(FullAdder_2908_io_s),
    .io_co(FullAdder_2908_io_co)
  );
  FullAdder FullAdder_2909 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2909_io_a),
    .io_b(FullAdder_2909_io_b),
    .io_ci(FullAdder_2909_io_ci),
    .io_s(FullAdder_2909_io_s),
    .io_co(FullAdder_2909_io_co)
  );
  FullAdder FullAdder_2910 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2910_io_a),
    .io_b(FullAdder_2910_io_b),
    .io_ci(FullAdder_2910_io_ci),
    .io_s(FullAdder_2910_io_s),
    .io_co(FullAdder_2910_io_co)
  );
  FullAdder FullAdder_2911 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2911_io_a),
    .io_b(FullAdder_2911_io_b),
    .io_ci(FullAdder_2911_io_ci),
    .io_s(FullAdder_2911_io_s),
    .io_co(FullAdder_2911_io_co)
  );
  FullAdder FullAdder_2912 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2912_io_a),
    .io_b(FullAdder_2912_io_b),
    .io_ci(FullAdder_2912_io_ci),
    .io_s(FullAdder_2912_io_s),
    .io_co(FullAdder_2912_io_co)
  );
  FullAdder FullAdder_2913 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2913_io_a),
    .io_b(FullAdder_2913_io_b),
    .io_ci(FullAdder_2913_io_ci),
    .io_s(FullAdder_2913_io_s),
    .io_co(FullAdder_2913_io_co)
  );
  FullAdder FullAdder_2914 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2914_io_a),
    .io_b(FullAdder_2914_io_b),
    .io_ci(FullAdder_2914_io_ci),
    .io_s(FullAdder_2914_io_s),
    .io_co(FullAdder_2914_io_co)
  );
  FullAdder FullAdder_2915 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2915_io_a),
    .io_b(FullAdder_2915_io_b),
    .io_ci(FullAdder_2915_io_ci),
    .io_s(FullAdder_2915_io_s),
    .io_co(FullAdder_2915_io_co)
  );
  FullAdder FullAdder_2916 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2916_io_a),
    .io_b(FullAdder_2916_io_b),
    .io_ci(FullAdder_2916_io_ci),
    .io_s(FullAdder_2916_io_s),
    .io_co(FullAdder_2916_io_co)
  );
  FullAdder FullAdder_2917 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2917_io_a),
    .io_b(FullAdder_2917_io_b),
    .io_ci(FullAdder_2917_io_ci),
    .io_s(FullAdder_2917_io_s),
    .io_co(FullAdder_2917_io_co)
  );
  FullAdder FullAdder_2918 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2918_io_a),
    .io_b(FullAdder_2918_io_b),
    .io_ci(FullAdder_2918_io_ci),
    .io_s(FullAdder_2918_io_s),
    .io_co(FullAdder_2918_io_co)
  );
  FullAdder FullAdder_2919 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2919_io_a),
    .io_b(FullAdder_2919_io_b),
    .io_ci(FullAdder_2919_io_ci),
    .io_s(FullAdder_2919_io_s),
    .io_co(FullAdder_2919_io_co)
  );
  FullAdder FullAdder_2920 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2920_io_a),
    .io_b(FullAdder_2920_io_b),
    .io_ci(FullAdder_2920_io_ci),
    .io_s(FullAdder_2920_io_s),
    .io_co(FullAdder_2920_io_co)
  );
  FullAdder FullAdder_2921 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2921_io_a),
    .io_b(FullAdder_2921_io_b),
    .io_ci(FullAdder_2921_io_ci),
    .io_s(FullAdder_2921_io_s),
    .io_co(FullAdder_2921_io_co)
  );
  FullAdder FullAdder_2922 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2922_io_a),
    .io_b(FullAdder_2922_io_b),
    .io_ci(FullAdder_2922_io_ci),
    .io_s(FullAdder_2922_io_s),
    .io_co(FullAdder_2922_io_co)
  );
  FullAdder FullAdder_2923 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2923_io_a),
    .io_b(FullAdder_2923_io_b),
    .io_ci(FullAdder_2923_io_ci),
    .io_s(FullAdder_2923_io_s),
    .io_co(FullAdder_2923_io_co)
  );
  FullAdder FullAdder_2924 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2924_io_a),
    .io_b(FullAdder_2924_io_b),
    .io_ci(FullAdder_2924_io_ci),
    .io_s(FullAdder_2924_io_s),
    .io_co(FullAdder_2924_io_co)
  );
  FullAdder FullAdder_2925 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2925_io_a),
    .io_b(FullAdder_2925_io_b),
    .io_ci(FullAdder_2925_io_ci),
    .io_s(FullAdder_2925_io_s),
    .io_co(FullAdder_2925_io_co)
  );
  FullAdder FullAdder_2926 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2926_io_a),
    .io_b(FullAdder_2926_io_b),
    .io_ci(FullAdder_2926_io_ci),
    .io_s(FullAdder_2926_io_s),
    .io_co(FullAdder_2926_io_co)
  );
  FullAdder FullAdder_2927 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2927_io_a),
    .io_b(FullAdder_2927_io_b),
    .io_ci(FullAdder_2927_io_ci),
    .io_s(FullAdder_2927_io_s),
    .io_co(FullAdder_2927_io_co)
  );
  FullAdder FullAdder_2928 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2928_io_a),
    .io_b(FullAdder_2928_io_b),
    .io_ci(FullAdder_2928_io_ci),
    .io_s(FullAdder_2928_io_s),
    .io_co(FullAdder_2928_io_co)
  );
  FullAdder FullAdder_2929 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2929_io_a),
    .io_b(FullAdder_2929_io_b),
    .io_ci(FullAdder_2929_io_ci),
    .io_s(FullAdder_2929_io_s),
    .io_co(FullAdder_2929_io_co)
  );
  FullAdder FullAdder_2930 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2930_io_a),
    .io_b(FullAdder_2930_io_b),
    .io_ci(FullAdder_2930_io_ci),
    .io_s(FullAdder_2930_io_s),
    .io_co(FullAdder_2930_io_co)
  );
  FullAdder FullAdder_2931 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2931_io_a),
    .io_b(FullAdder_2931_io_b),
    .io_ci(FullAdder_2931_io_ci),
    .io_s(FullAdder_2931_io_s),
    .io_co(FullAdder_2931_io_co)
  );
  FullAdder FullAdder_2932 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2932_io_a),
    .io_b(FullAdder_2932_io_b),
    .io_ci(FullAdder_2932_io_ci),
    .io_s(FullAdder_2932_io_s),
    .io_co(FullAdder_2932_io_co)
  );
  HalfAdder HalfAdder_102 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_102_io_a),
    .io_b(HalfAdder_102_io_b),
    .io_s(HalfAdder_102_io_s),
    .io_co(HalfAdder_102_io_co)
  );
  FullAdder FullAdder_2933 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2933_io_a),
    .io_b(FullAdder_2933_io_b),
    .io_ci(FullAdder_2933_io_ci),
    .io_s(FullAdder_2933_io_s),
    .io_co(FullAdder_2933_io_co)
  );
  FullAdder FullAdder_2934 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2934_io_a),
    .io_b(FullAdder_2934_io_b),
    .io_ci(FullAdder_2934_io_ci),
    .io_s(FullAdder_2934_io_s),
    .io_co(FullAdder_2934_io_co)
  );
  FullAdder FullAdder_2935 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2935_io_a),
    .io_b(FullAdder_2935_io_b),
    .io_ci(FullAdder_2935_io_ci),
    .io_s(FullAdder_2935_io_s),
    .io_co(FullAdder_2935_io_co)
  );
  FullAdder FullAdder_2936 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2936_io_a),
    .io_b(FullAdder_2936_io_b),
    .io_ci(FullAdder_2936_io_ci),
    .io_s(FullAdder_2936_io_s),
    .io_co(FullAdder_2936_io_co)
  );
  FullAdder FullAdder_2937 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2937_io_a),
    .io_b(FullAdder_2937_io_b),
    .io_ci(FullAdder_2937_io_ci),
    .io_s(FullAdder_2937_io_s),
    .io_co(FullAdder_2937_io_co)
  );
  FullAdder FullAdder_2938 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2938_io_a),
    .io_b(FullAdder_2938_io_b),
    .io_ci(FullAdder_2938_io_ci),
    .io_s(FullAdder_2938_io_s),
    .io_co(FullAdder_2938_io_co)
  );
  FullAdder FullAdder_2939 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2939_io_a),
    .io_b(FullAdder_2939_io_b),
    .io_ci(FullAdder_2939_io_ci),
    .io_s(FullAdder_2939_io_s),
    .io_co(FullAdder_2939_io_co)
  );
  FullAdder FullAdder_2940 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2940_io_a),
    .io_b(FullAdder_2940_io_b),
    .io_ci(FullAdder_2940_io_ci),
    .io_s(FullAdder_2940_io_s),
    .io_co(FullAdder_2940_io_co)
  );
  FullAdder FullAdder_2941 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2941_io_a),
    .io_b(FullAdder_2941_io_b),
    .io_ci(FullAdder_2941_io_ci),
    .io_s(FullAdder_2941_io_s),
    .io_co(FullAdder_2941_io_co)
  );
  FullAdder FullAdder_2942 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2942_io_a),
    .io_b(FullAdder_2942_io_b),
    .io_ci(FullAdder_2942_io_ci),
    .io_s(FullAdder_2942_io_s),
    .io_co(FullAdder_2942_io_co)
  );
  FullAdder FullAdder_2943 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2943_io_a),
    .io_b(FullAdder_2943_io_b),
    .io_ci(FullAdder_2943_io_ci),
    .io_s(FullAdder_2943_io_s),
    .io_co(FullAdder_2943_io_co)
  );
  FullAdder FullAdder_2944 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2944_io_a),
    .io_b(FullAdder_2944_io_b),
    .io_ci(FullAdder_2944_io_ci),
    .io_s(FullAdder_2944_io_s),
    .io_co(FullAdder_2944_io_co)
  );
  FullAdder FullAdder_2945 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2945_io_a),
    .io_b(FullAdder_2945_io_b),
    .io_ci(FullAdder_2945_io_ci),
    .io_s(FullAdder_2945_io_s),
    .io_co(FullAdder_2945_io_co)
  );
  FullAdder FullAdder_2946 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2946_io_a),
    .io_b(FullAdder_2946_io_b),
    .io_ci(FullAdder_2946_io_ci),
    .io_s(FullAdder_2946_io_s),
    .io_co(FullAdder_2946_io_co)
  );
  FullAdder FullAdder_2947 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2947_io_a),
    .io_b(FullAdder_2947_io_b),
    .io_ci(FullAdder_2947_io_ci),
    .io_s(FullAdder_2947_io_s),
    .io_co(FullAdder_2947_io_co)
  );
  FullAdder FullAdder_2948 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2948_io_a),
    .io_b(FullAdder_2948_io_b),
    .io_ci(FullAdder_2948_io_ci),
    .io_s(FullAdder_2948_io_s),
    .io_co(FullAdder_2948_io_co)
  );
  FullAdder FullAdder_2949 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2949_io_a),
    .io_b(FullAdder_2949_io_b),
    .io_ci(FullAdder_2949_io_ci),
    .io_s(FullAdder_2949_io_s),
    .io_co(FullAdder_2949_io_co)
  );
  FullAdder FullAdder_2950 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2950_io_a),
    .io_b(FullAdder_2950_io_b),
    .io_ci(FullAdder_2950_io_ci),
    .io_s(FullAdder_2950_io_s),
    .io_co(FullAdder_2950_io_co)
  );
  FullAdder FullAdder_2951 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2951_io_a),
    .io_b(FullAdder_2951_io_b),
    .io_ci(FullAdder_2951_io_ci),
    .io_s(FullAdder_2951_io_s),
    .io_co(FullAdder_2951_io_co)
  );
  FullAdder FullAdder_2952 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2952_io_a),
    .io_b(FullAdder_2952_io_b),
    .io_ci(FullAdder_2952_io_ci),
    .io_s(FullAdder_2952_io_s),
    .io_co(FullAdder_2952_io_co)
  );
  FullAdder FullAdder_2953 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2953_io_a),
    .io_b(FullAdder_2953_io_b),
    .io_ci(FullAdder_2953_io_ci),
    .io_s(FullAdder_2953_io_s),
    .io_co(FullAdder_2953_io_co)
  );
  FullAdder FullAdder_2954 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2954_io_a),
    .io_b(FullAdder_2954_io_b),
    .io_ci(FullAdder_2954_io_ci),
    .io_s(FullAdder_2954_io_s),
    .io_co(FullAdder_2954_io_co)
  );
  FullAdder FullAdder_2955 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2955_io_a),
    .io_b(FullAdder_2955_io_b),
    .io_ci(FullAdder_2955_io_ci),
    .io_s(FullAdder_2955_io_s),
    .io_co(FullAdder_2955_io_co)
  );
  FullAdder FullAdder_2956 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2956_io_a),
    .io_b(FullAdder_2956_io_b),
    .io_ci(FullAdder_2956_io_ci),
    .io_s(FullAdder_2956_io_s),
    .io_co(FullAdder_2956_io_co)
  );
  FullAdder FullAdder_2957 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2957_io_a),
    .io_b(FullAdder_2957_io_b),
    .io_ci(FullAdder_2957_io_ci),
    .io_s(FullAdder_2957_io_s),
    .io_co(FullAdder_2957_io_co)
  );
  FullAdder FullAdder_2958 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2958_io_a),
    .io_b(FullAdder_2958_io_b),
    .io_ci(FullAdder_2958_io_ci),
    .io_s(FullAdder_2958_io_s),
    .io_co(FullAdder_2958_io_co)
  );
  FullAdder FullAdder_2959 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2959_io_a),
    .io_b(FullAdder_2959_io_b),
    .io_ci(FullAdder_2959_io_ci),
    .io_s(FullAdder_2959_io_s),
    .io_co(FullAdder_2959_io_co)
  );
  FullAdder FullAdder_2960 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2960_io_a),
    .io_b(FullAdder_2960_io_b),
    .io_ci(FullAdder_2960_io_ci),
    .io_s(FullAdder_2960_io_s),
    .io_co(FullAdder_2960_io_co)
  );
  FullAdder FullAdder_2961 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2961_io_a),
    .io_b(FullAdder_2961_io_b),
    .io_ci(FullAdder_2961_io_ci),
    .io_s(FullAdder_2961_io_s),
    .io_co(FullAdder_2961_io_co)
  );
  FullAdder FullAdder_2962 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2962_io_a),
    .io_b(FullAdder_2962_io_b),
    .io_ci(FullAdder_2962_io_ci),
    .io_s(FullAdder_2962_io_s),
    .io_co(FullAdder_2962_io_co)
  );
  FullAdder FullAdder_2963 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2963_io_a),
    .io_b(FullAdder_2963_io_b),
    .io_ci(FullAdder_2963_io_ci),
    .io_s(FullAdder_2963_io_s),
    .io_co(FullAdder_2963_io_co)
  );
  FullAdder FullAdder_2964 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2964_io_a),
    .io_b(FullAdder_2964_io_b),
    .io_ci(FullAdder_2964_io_ci),
    .io_s(FullAdder_2964_io_s),
    .io_co(FullAdder_2964_io_co)
  );
  FullAdder FullAdder_2965 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2965_io_a),
    .io_b(FullAdder_2965_io_b),
    .io_ci(FullAdder_2965_io_ci),
    .io_s(FullAdder_2965_io_s),
    .io_co(FullAdder_2965_io_co)
  );
  FullAdder FullAdder_2966 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2966_io_a),
    .io_b(FullAdder_2966_io_b),
    .io_ci(FullAdder_2966_io_ci),
    .io_s(FullAdder_2966_io_s),
    .io_co(FullAdder_2966_io_co)
  );
  FullAdder FullAdder_2967 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2967_io_a),
    .io_b(FullAdder_2967_io_b),
    .io_ci(FullAdder_2967_io_ci),
    .io_s(FullAdder_2967_io_s),
    .io_co(FullAdder_2967_io_co)
  );
  FullAdder FullAdder_2968 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2968_io_a),
    .io_b(FullAdder_2968_io_b),
    .io_ci(FullAdder_2968_io_ci),
    .io_s(FullAdder_2968_io_s),
    .io_co(FullAdder_2968_io_co)
  );
  FullAdder FullAdder_2969 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2969_io_a),
    .io_b(FullAdder_2969_io_b),
    .io_ci(FullAdder_2969_io_ci),
    .io_s(FullAdder_2969_io_s),
    .io_co(FullAdder_2969_io_co)
  );
  FullAdder FullAdder_2970 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2970_io_a),
    .io_b(FullAdder_2970_io_b),
    .io_ci(FullAdder_2970_io_ci),
    .io_s(FullAdder_2970_io_s),
    .io_co(FullAdder_2970_io_co)
  );
  FullAdder FullAdder_2971 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2971_io_a),
    .io_b(FullAdder_2971_io_b),
    .io_ci(FullAdder_2971_io_ci),
    .io_s(FullAdder_2971_io_s),
    .io_co(FullAdder_2971_io_co)
  );
  FullAdder FullAdder_2972 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2972_io_a),
    .io_b(FullAdder_2972_io_b),
    .io_ci(FullAdder_2972_io_ci),
    .io_s(FullAdder_2972_io_s),
    .io_co(FullAdder_2972_io_co)
  );
  FullAdder FullAdder_2973 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2973_io_a),
    .io_b(FullAdder_2973_io_b),
    .io_ci(FullAdder_2973_io_ci),
    .io_s(FullAdder_2973_io_s),
    .io_co(FullAdder_2973_io_co)
  );
  FullAdder FullAdder_2974 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2974_io_a),
    .io_b(FullAdder_2974_io_b),
    .io_ci(FullAdder_2974_io_ci),
    .io_s(FullAdder_2974_io_s),
    .io_co(FullAdder_2974_io_co)
  );
  FullAdder FullAdder_2975 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2975_io_a),
    .io_b(FullAdder_2975_io_b),
    .io_ci(FullAdder_2975_io_ci),
    .io_s(FullAdder_2975_io_s),
    .io_co(FullAdder_2975_io_co)
  );
  FullAdder FullAdder_2976 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2976_io_a),
    .io_b(FullAdder_2976_io_b),
    .io_ci(FullAdder_2976_io_ci),
    .io_s(FullAdder_2976_io_s),
    .io_co(FullAdder_2976_io_co)
  );
  FullAdder FullAdder_2977 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2977_io_a),
    .io_b(FullAdder_2977_io_b),
    .io_ci(FullAdder_2977_io_ci),
    .io_s(FullAdder_2977_io_s),
    .io_co(FullAdder_2977_io_co)
  );
  FullAdder FullAdder_2978 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2978_io_a),
    .io_b(FullAdder_2978_io_b),
    .io_ci(FullAdder_2978_io_ci),
    .io_s(FullAdder_2978_io_s),
    .io_co(FullAdder_2978_io_co)
  );
  FullAdder FullAdder_2979 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2979_io_a),
    .io_b(FullAdder_2979_io_b),
    .io_ci(FullAdder_2979_io_ci),
    .io_s(FullAdder_2979_io_s),
    .io_co(FullAdder_2979_io_co)
  );
  FullAdder FullAdder_2980 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2980_io_a),
    .io_b(FullAdder_2980_io_b),
    .io_ci(FullAdder_2980_io_ci),
    .io_s(FullAdder_2980_io_s),
    .io_co(FullAdder_2980_io_co)
  );
  FullAdder FullAdder_2981 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2981_io_a),
    .io_b(FullAdder_2981_io_b),
    .io_ci(FullAdder_2981_io_ci),
    .io_s(FullAdder_2981_io_s),
    .io_co(FullAdder_2981_io_co)
  );
  FullAdder FullAdder_2982 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2982_io_a),
    .io_b(FullAdder_2982_io_b),
    .io_ci(FullAdder_2982_io_ci),
    .io_s(FullAdder_2982_io_s),
    .io_co(FullAdder_2982_io_co)
  );
  FullAdder FullAdder_2983 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2983_io_a),
    .io_b(FullAdder_2983_io_b),
    .io_ci(FullAdder_2983_io_ci),
    .io_s(FullAdder_2983_io_s),
    .io_co(FullAdder_2983_io_co)
  );
  FullAdder FullAdder_2984 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2984_io_a),
    .io_b(FullAdder_2984_io_b),
    .io_ci(FullAdder_2984_io_ci),
    .io_s(FullAdder_2984_io_s),
    .io_co(FullAdder_2984_io_co)
  );
  FullAdder FullAdder_2985 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2985_io_a),
    .io_b(FullAdder_2985_io_b),
    .io_ci(FullAdder_2985_io_ci),
    .io_s(FullAdder_2985_io_s),
    .io_co(FullAdder_2985_io_co)
  );
  FullAdder FullAdder_2986 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2986_io_a),
    .io_b(FullAdder_2986_io_b),
    .io_ci(FullAdder_2986_io_ci),
    .io_s(FullAdder_2986_io_s),
    .io_co(FullAdder_2986_io_co)
  );
  HalfAdder HalfAdder_103 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_103_io_a),
    .io_b(HalfAdder_103_io_b),
    .io_s(HalfAdder_103_io_s),
    .io_co(HalfAdder_103_io_co)
  );
  FullAdder FullAdder_2987 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2987_io_a),
    .io_b(FullAdder_2987_io_b),
    .io_ci(FullAdder_2987_io_ci),
    .io_s(FullAdder_2987_io_s),
    .io_co(FullAdder_2987_io_co)
  );
  FullAdder FullAdder_2988 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2988_io_a),
    .io_b(FullAdder_2988_io_b),
    .io_ci(FullAdder_2988_io_ci),
    .io_s(FullAdder_2988_io_s),
    .io_co(FullAdder_2988_io_co)
  );
  FullAdder FullAdder_2989 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2989_io_a),
    .io_b(FullAdder_2989_io_b),
    .io_ci(FullAdder_2989_io_ci),
    .io_s(FullAdder_2989_io_s),
    .io_co(FullAdder_2989_io_co)
  );
  FullAdder FullAdder_2990 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2990_io_a),
    .io_b(FullAdder_2990_io_b),
    .io_ci(FullAdder_2990_io_ci),
    .io_s(FullAdder_2990_io_s),
    .io_co(FullAdder_2990_io_co)
  );
  FullAdder FullAdder_2991 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2991_io_a),
    .io_b(FullAdder_2991_io_b),
    .io_ci(FullAdder_2991_io_ci),
    .io_s(FullAdder_2991_io_s),
    .io_co(FullAdder_2991_io_co)
  );
  FullAdder FullAdder_2992 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2992_io_a),
    .io_b(FullAdder_2992_io_b),
    .io_ci(FullAdder_2992_io_ci),
    .io_s(FullAdder_2992_io_s),
    .io_co(FullAdder_2992_io_co)
  );
  FullAdder FullAdder_2993 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2993_io_a),
    .io_b(FullAdder_2993_io_b),
    .io_ci(FullAdder_2993_io_ci),
    .io_s(FullAdder_2993_io_s),
    .io_co(FullAdder_2993_io_co)
  );
  FullAdder FullAdder_2994 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2994_io_a),
    .io_b(FullAdder_2994_io_b),
    .io_ci(FullAdder_2994_io_ci),
    .io_s(FullAdder_2994_io_s),
    .io_co(FullAdder_2994_io_co)
  );
  FullAdder FullAdder_2995 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2995_io_a),
    .io_b(FullAdder_2995_io_b),
    .io_ci(FullAdder_2995_io_ci),
    .io_s(FullAdder_2995_io_s),
    .io_co(FullAdder_2995_io_co)
  );
  FullAdder FullAdder_2996 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2996_io_a),
    .io_b(FullAdder_2996_io_b),
    .io_ci(FullAdder_2996_io_ci),
    .io_s(FullAdder_2996_io_s),
    .io_co(FullAdder_2996_io_co)
  );
  FullAdder FullAdder_2997 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2997_io_a),
    .io_b(FullAdder_2997_io_b),
    .io_ci(FullAdder_2997_io_ci),
    .io_s(FullAdder_2997_io_s),
    .io_co(FullAdder_2997_io_co)
  );
  FullAdder FullAdder_2998 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2998_io_a),
    .io_b(FullAdder_2998_io_b),
    .io_ci(FullAdder_2998_io_ci),
    .io_s(FullAdder_2998_io_s),
    .io_co(FullAdder_2998_io_co)
  );
  FullAdder FullAdder_2999 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_2999_io_a),
    .io_b(FullAdder_2999_io_b),
    .io_ci(FullAdder_2999_io_ci),
    .io_s(FullAdder_2999_io_s),
    .io_co(FullAdder_2999_io_co)
  );
  FullAdder FullAdder_3000 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3000_io_a),
    .io_b(FullAdder_3000_io_b),
    .io_ci(FullAdder_3000_io_ci),
    .io_s(FullAdder_3000_io_s),
    .io_co(FullAdder_3000_io_co)
  );
  FullAdder FullAdder_3001 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3001_io_a),
    .io_b(FullAdder_3001_io_b),
    .io_ci(FullAdder_3001_io_ci),
    .io_s(FullAdder_3001_io_s),
    .io_co(FullAdder_3001_io_co)
  );
  FullAdder FullAdder_3002 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3002_io_a),
    .io_b(FullAdder_3002_io_b),
    .io_ci(FullAdder_3002_io_ci),
    .io_s(FullAdder_3002_io_s),
    .io_co(FullAdder_3002_io_co)
  );
  FullAdder FullAdder_3003 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3003_io_a),
    .io_b(FullAdder_3003_io_b),
    .io_ci(FullAdder_3003_io_ci),
    .io_s(FullAdder_3003_io_s),
    .io_co(FullAdder_3003_io_co)
  );
  FullAdder FullAdder_3004 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3004_io_a),
    .io_b(FullAdder_3004_io_b),
    .io_ci(FullAdder_3004_io_ci),
    .io_s(FullAdder_3004_io_s),
    .io_co(FullAdder_3004_io_co)
  );
  FullAdder FullAdder_3005 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3005_io_a),
    .io_b(FullAdder_3005_io_b),
    .io_ci(FullAdder_3005_io_ci),
    .io_s(FullAdder_3005_io_s),
    .io_co(FullAdder_3005_io_co)
  );
  FullAdder FullAdder_3006 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3006_io_a),
    .io_b(FullAdder_3006_io_b),
    .io_ci(FullAdder_3006_io_ci),
    .io_s(FullAdder_3006_io_s),
    .io_co(FullAdder_3006_io_co)
  );
  FullAdder FullAdder_3007 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3007_io_a),
    .io_b(FullAdder_3007_io_b),
    .io_ci(FullAdder_3007_io_ci),
    .io_s(FullAdder_3007_io_s),
    .io_co(FullAdder_3007_io_co)
  );
  FullAdder FullAdder_3008 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3008_io_a),
    .io_b(FullAdder_3008_io_b),
    .io_ci(FullAdder_3008_io_ci),
    .io_s(FullAdder_3008_io_s),
    .io_co(FullAdder_3008_io_co)
  );
  FullAdder FullAdder_3009 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3009_io_a),
    .io_b(FullAdder_3009_io_b),
    .io_ci(FullAdder_3009_io_ci),
    .io_s(FullAdder_3009_io_s),
    .io_co(FullAdder_3009_io_co)
  );
  FullAdder FullAdder_3010 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3010_io_a),
    .io_b(FullAdder_3010_io_b),
    .io_ci(FullAdder_3010_io_ci),
    .io_s(FullAdder_3010_io_s),
    .io_co(FullAdder_3010_io_co)
  );
  FullAdder FullAdder_3011 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3011_io_a),
    .io_b(FullAdder_3011_io_b),
    .io_ci(FullAdder_3011_io_ci),
    .io_s(FullAdder_3011_io_s),
    .io_co(FullAdder_3011_io_co)
  );
  FullAdder FullAdder_3012 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3012_io_a),
    .io_b(FullAdder_3012_io_b),
    .io_ci(FullAdder_3012_io_ci),
    .io_s(FullAdder_3012_io_s),
    .io_co(FullAdder_3012_io_co)
  );
  FullAdder FullAdder_3013 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3013_io_a),
    .io_b(FullAdder_3013_io_b),
    .io_ci(FullAdder_3013_io_ci),
    .io_s(FullAdder_3013_io_s),
    .io_co(FullAdder_3013_io_co)
  );
  FullAdder FullAdder_3014 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3014_io_a),
    .io_b(FullAdder_3014_io_b),
    .io_ci(FullAdder_3014_io_ci),
    .io_s(FullAdder_3014_io_s),
    .io_co(FullAdder_3014_io_co)
  );
  FullAdder FullAdder_3015 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3015_io_a),
    .io_b(FullAdder_3015_io_b),
    .io_ci(FullAdder_3015_io_ci),
    .io_s(FullAdder_3015_io_s),
    .io_co(FullAdder_3015_io_co)
  );
  FullAdder FullAdder_3016 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3016_io_a),
    .io_b(FullAdder_3016_io_b),
    .io_ci(FullAdder_3016_io_ci),
    .io_s(FullAdder_3016_io_s),
    .io_co(FullAdder_3016_io_co)
  );
  FullAdder FullAdder_3017 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3017_io_a),
    .io_b(FullAdder_3017_io_b),
    .io_ci(FullAdder_3017_io_ci),
    .io_s(FullAdder_3017_io_s),
    .io_co(FullAdder_3017_io_co)
  );
  FullAdder FullAdder_3018 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3018_io_a),
    .io_b(FullAdder_3018_io_b),
    .io_ci(FullAdder_3018_io_ci),
    .io_s(FullAdder_3018_io_s),
    .io_co(FullAdder_3018_io_co)
  );
  FullAdder FullAdder_3019 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3019_io_a),
    .io_b(FullAdder_3019_io_b),
    .io_ci(FullAdder_3019_io_ci),
    .io_s(FullAdder_3019_io_s),
    .io_co(FullAdder_3019_io_co)
  );
  FullAdder FullAdder_3020 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3020_io_a),
    .io_b(FullAdder_3020_io_b),
    .io_ci(FullAdder_3020_io_ci),
    .io_s(FullAdder_3020_io_s),
    .io_co(FullAdder_3020_io_co)
  );
  FullAdder FullAdder_3021 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3021_io_a),
    .io_b(FullAdder_3021_io_b),
    .io_ci(FullAdder_3021_io_ci),
    .io_s(FullAdder_3021_io_s),
    .io_co(FullAdder_3021_io_co)
  );
  FullAdder FullAdder_3022 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3022_io_a),
    .io_b(FullAdder_3022_io_b),
    .io_ci(FullAdder_3022_io_ci),
    .io_s(FullAdder_3022_io_s),
    .io_co(FullAdder_3022_io_co)
  );
  FullAdder FullAdder_3023 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3023_io_a),
    .io_b(FullAdder_3023_io_b),
    .io_ci(FullAdder_3023_io_ci),
    .io_s(FullAdder_3023_io_s),
    .io_co(FullAdder_3023_io_co)
  );
  FullAdder FullAdder_3024 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3024_io_a),
    .io_b(FullAdder_3024_io_b),
    .io_ci(FullAdder_3024_io_ci),
    .io_s(FullAdder_3024_io_s),
    .io_co(FullAdder_3024_io_co)
  );
  FullAdder FullAdder_3025 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3025_io_a),
    .io_b(FullAdder_3025_io_b),
    .io_ci(FullAdder_3025_io_ci),
    .io_s(FullAdder_3025_io_s),
    .io_co(FullAdder_3025_io_co)
  );
  FullAdder FullAdder_3026 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3026_io_a),
    .io_b(FullAdder_3026_io_b),
    .io_ci(FullAdder_3026_io_ci),
    .io_s(FullAdder_3026_io_s),
    .io_co(FullAdder_3026_io_co)
  );
  HalfAdder HalfAdder_104 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_104_io_a),
    .io_b(HalfAdder_104_io_b),
    .io_s(HalfAdder_104_io_s),
    .io_co(HalfAdder_104_io_co)
  );
  FullAdder FullAdder_3027 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3027_io_a),
    .io_b(FullAdder_3027_io_b),
    .io_ci(FullAdder_3027_io_ci),
    .io_s(FullAdder_3027_io_s),
    .io_co(FullAdder_3027_io_co)
  );
  FullAdder FullAdder_3028 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3028_io_a),
    .io_b(FullAdder_3028_io_b),
    .io_ci(FullAdder_3028_io_ci),
    .io_s(FullAdder_3028_io_s),
    .io_co(FullAdder_3028_io_co)
  );
  FullAdder FullAdder_3029 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3029_io_a),
    .io_b(FullAdder_3029_io_b),
    .io_ci(FullAdder_3029_io_ci),
    .io_s(FullAdder_3029_io_s),
    .io_co(FullAdder_3029_io_co)
  );
  FullAdder FullAdder_3030 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3030_io_a),
    .io_b(FullAdder_3030_io_b),
    .io_ci(FullAdder_3030_io_ci),
    .io_s(FullAdder_3030_io_s),
    .io_co(FullAdder_3030_io_co)
  );
  FullAdder FullAdder_3031 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3031_io_a),
    .io_b(FullAdder_3031_io_b),
    .io_ci(FullAdder_3031_io_ci),
    .io_s(FullAdder_3031_io_s),
    .io_co(FullAdder_3031_io_co)
  );
  HalfAdder HalfAdder_105 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_105_io_a),
    .io_b(HalfAdder_105_io_b),
    .io_s(HalfAdder_105_io_s),
    .io_co(HalfAdder_105_io_co)
  );
  FullAdder FullAdder_3032 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3032_io_a),
    .io_b(FullAdder_3032_io_b),
    .io_ci(FullAdder_3032_io_ci),
    .io_s(FullAdder_3032_io_s),
    .io_co(FullAdder_3032_io_co)
  );
  FullAdder FullAdder_3033 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3033_io_a),
    .io_b(FullAdder_3033_io_b),
    .io_ci(FullAdder_3033_io_ci),
    .io_s(FullAdder_3033_io_s),
    .io_co(FullAdder_3033_io_co)
  );
  FullAdder FullAdder_3034 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3034_io_a),
    .io_b(FullAdder_3034_io_b),
    .io_ci(FullAdder_3034_io_ci),
    .io_s(FullAdder_3034_io_s),
    .io_co(FullAdder_3034_io_co)
  );
  FullAdder FullAdder_3035 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3035_io_a),
    .io_b(FullAdder_3035_io_b),
    .io_ci(FullAdder_3035_io_ci),
    .io_s(FullAdder_3035_io_s),
    .io_co(FullAdder_3035_io_co)
  );
  FullAdder FullAdder_3036 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3036_io_a),
    .io_b(FullAdder_3036_io_b),
    .io_ci(FullAdder_3036_io_ci),
    .io_s(FullAdder_3036_io_s),
    .io_co(FullAdder_3036_io_co)
  );
  FullAdder FullAdder_3037 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3037_io_a),
    .io_b(FullAdder_3037_io_b),
    .io_ci(FullAdder_3037_io_ci),
    .io_s(FullAdder_3037_io_s),
    .io_co(FullAdder_3037_io_co)
  );
  FullAdder FullAdder_3038 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3038_io_a),
    .io_b(FullAdder_3038_io_b),
    .io_ci(FullAdder_3038_io_ci),
    .io_s(FullAdder_3038_io_s),
    .io_co(FullAdder_3038_io_co)
  );
  FullAdder FullAdder_3039 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3039_io_a),
    .io_b(FullAdder_3039_io_b),
    .io_ci(FullAdder_3039_io_ci),
    .io_s(FullAdder_3039_io_s),
    .io_co(FullAdder_3039_io_co)
  );
  FullAdder FullAdder_3040 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3040_io_a),
    .io_b(FullAdder_3040_io_b),
    .io_ci(FullAdder_3040_io_ci),
    .io_s(FullAdder_3040_io_s),
    .io_co(FullAdder_3040_io_co)
  );
  FullAdder FullAdder_3041 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3041_io_a),
    .io_b(FullAdder_3041_io_b),
    .io_ci(FullAdder_3041_io_ci),
    .io_s(FullAdder_3041_io_s),
    .io_co(FullAdder_3041_io_co)
  );
  FullAdder FullAdder_3042 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3042_io_a),
    .io_b(FullAdder_3042_io_b),
    .io_ci(FullAdder_3042_io_ci),
    .io_s(FullAdder_3042_io_s),
    .io_co(FullAdder_3042_io_co)
  );
  FullAdder FullAdder_3043 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3043_io_a),
    .io_b(FullAdder_3043_io_b),
    .io_ci(FullAdder_3043_io_ci),
    .io_s(FullAdder_3043_io_s),
    .io_co(FullAdder_3043_io_co)
  );
  FullAdder FullAdder_3044 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3044_io_a),
    .io_b(FullAdder_3044_io_b),
    .io_ci(FullAdder_3044_io_ci),
    .io_s(FullAdder_3044_io_s),
    .io_co(FullAdder_3044_io_co)
  );
  FullAdder FullAdder_3045 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3045_io_a),
    .io_b(FullAdder_3045_io_b),
    .io_ci(FullAdder_3045_io_ci),
    .io_s(FullAdder_3045_io_s),
    .io_co(FullAdder_3045_io_co)
  );
  FullAdder FullAdder_3046 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3046_io_a),
    .io_b(FullAdder_3046_io_b),
    .io_ci(FullAdder_3046_io_ci),
    .io_s(FullAdder_3046_io_s),
    .io_co(FullAdder_3046_io_co)
  );
  FullAdder FullAdder_3047 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3047_io_a),
    .io_b(FullAdder_3047_io_b),
    .io_ci(FullAdder_3047_io_ci),
    .io_s(FullAdder_3047_io_s),
    .io_co(FullAdder_3047_io_co)
  );
  FullAdder FullAdder_3048 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3048_io_a),
    .io_b(FullAdder_3048_io_b),
    .io_ci(FullAdder_3048_io_ci),
    .io_s(FullAdder_3048_io_s),
    .io_co(FullAdder_3048_io_co)
  );
  FullAdder FullAdder_3049 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3049_io_a),
    .io_b(FullAdder_3049_io_b),
    .io_ci(FullAdder_3049_io_ci),
    .io_s(FullAdder_3049_io_s),
    .io_co(FullAdder_3049_io_co)
  );
  FullAdder FullAdder_3050 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3050_io_a),
    .io_b(FullAdder_3050_io_b),
    .io_ci(FullAdder_3050_io_ci),
    .io_s(FullAdder_3050_io_s),
    .io_co(FullAdder_3050_io_co)
  );
  FullAdder FullAdder_3051 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3051_io_a),
    .io_b(FullAdder_3051_io_b),
    .io_ci(FullAdder_3051_io_ci),
    .io_s(FullAdder_3051_io_s),
    .io_co(FullAdder_3051_io_co)
  );
  FullAdder FullAdder_3052 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3052_io_a),
    .io_b(FullAdder_3052_io_b),
    .io_ci(FullAdder_3052_io_ci),
    .io_s(FullAdder_3052_io_s),
    .io_co(FullAdder_3052_io_co)
  );
  FullAdder FullAdder_3053 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3053_io_a),
    .io_b(FullAdder_3053_io_b),
    .io_ci(FullAdder_3053_io_ci),
    .io_s(FullAdder_3053_io_s),
    .io_co(FullAdder_3053_io_co)
  );
  FullAdder FullAdder_3054 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3054_io_a),
    .io_b(FullAdder_3054_io_b),
    .io_ci(FullAdder_3054_io_ci),
    .io_s(FullAdder_3054_io_s),
    .io_co(FullAdder_3054_io_co)
  );
  FullAdder FullAdder_3055 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3055_io_a),
    .io_b(FullAdder_3055_io_b),
    .io_ci(FullAdder_3055_io_ci),
    .io_s(FullAdder_3055_io_s),
    .io_co(FullAdder_3055_io_co)
  );
  FullAdder FullAdder_3056 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3056_io_a),
    .io_b(FullAdder_3056_io_b),
    .io_ci(FullAdder_3056_io_ci),
    .io_s(FullAdder_3056_io_s),
    .io_co(FullAdder_3056_io_co)
  );
  FullAdder FullAdder_3057 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3057_io_a),
    .io_b(FullAdder_3057_io_b),
    .io_ci(FullAdder_3057_io_ci),
    .io_s(FullAdder_3057_io_s),
    .io_co(FullAdder_3057_io_co)
  );
  FullAdder FullAdder_3058 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3058_io_a),
    .io_b(FullAdder_3058_io_b),
    .io_ci(FullAdder_3058_io_ci),
    .io_s(FullAdder_3058_io_s),
    .io_co(FullAdder_3058_io_co)
  );
  FullAdder FullAdder_3059 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3059_io_a),
    .io_b(FullAdder_3059_io_b),
    .io_ci(FullAdder_3059_io_ci),
    .io_s(FullAdder_3059_io_s),
    .io_co(FullAdder_3059_io_co)
  );
  FullAdder FullAdder_3060 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3060_io_a),
    .io_b(FullAdder_3060_io_b),
    .io_ci(FullAdder_3060_io_ci),
    .io_s(FullAdder_3060_io_s),
    .io_co(FullAdder_3060_io_co)
  );
  FullAdder FullAdder_3061 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3061_io_a),
    .io_b(FullAdder_3061_io_b),
    .io_ci(FullAdder_3061_io_ci),
    .io_s(FullAdder_3061_io_s),
    .io_co(FullAdder_3061_io_co)
  );
  FullAdder FullAdder_3062 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3062_io_a),
    .io_b(FullAdder_3062_io_b),
    .io_ci(FullAdder_3062_io_ci),
    .io_s(FullAdder_3062_io_s),
    .io_co(FullAdder_3062_io_co)
  );
  FullAdder FullAdder_3063 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3063_io_a),
    .io_b(FullAdder_3063_io_b),
    .io_ci(FullAdder_3063_io_ci),
    .io_s(FullAdder_3063_io_s),
    .io_co(FullAdder_3063_io_co)
  );
  FullAdder FullAdder_3064 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3064_io_a),
    .io_b(FullAdder_3064_io_b),
    .io_ci(FullAdder_3064_io_ci),
    .io_s(FullAdder_3064_io_s),
    .io_co(FullAdder_3064_io_co)
  );
  FullAdder FullAdder_3065 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3065_io_a),
    .io_b(FullAdder_3065_io_b),
    .io_ci(FullAdder_3065_io_ci),
    .io_s(FullAdder_3065_io_s),
    .io_co(FullAdder_3065_io_co)
  );
  FullAdder FullAdder_3066 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3066_io_a),
    .io_b(FullAdder_3066_io_b),
    .io_ci(FullAdder_3066_io_ci),
    .io_s(FullAdder_3066_io_s),
    .io_co(FullAdder_3066_io_co)
  );
  FullAdder FullAdder_3067 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3067_io_a),
    .io_b(FullAdder_3067_io_b),
    .io_ci(FullAdder_3067_io_ci),
    .io_s(FullAdder_3067_io_s),
    .io_co(FullAdder_3067_io_co)
  );
  FullAdder FullAdder_3068 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3068_io_a),
    .io_b(FullAdder_3068_io_b),
    .io_ci(FullAdder_3068_io_ci),
    .io_s(FullAdder_3068_io_s),
    .io_co(FullAdder_3068_io_co)
  );
  FullAdder FullAdder_3069 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3069_io_a),
    .io_b(FullAdder_3069_io_b),
    .io_ci(FullAdder_3069_io_ci),
    .io_s(FullAdder_3069_io_s),
    .io_co(FullAdder_3069_io_co)
  );
  FullAdder FullAdder_3070 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3070_io_a),
    .io_b(FullAdder_3070_io_b),
    .io_ci(FullAdder_3070_io_ci),
    .io_s(FullAdder_3070_io_s),
    .io_co(FullAdder_3070_io_co)
  );
  FullAdder FullAdder_3071 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3071_io_a),
    .io_b(FullAdder_3071_io_b),
    .io_ci(FullAdder_3071_io_ci),
    .io_s(FullAdder_3071_io_s),
    .io_co(FullAdder_3071_io_co)
  );
  FullAdder FullAdder_3072 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3072_io_a),
    .io_b(FullAdder_3072_io_b),
    .io_ci(FullAdder_3072_io_ci),
    .io_s(FullAdder_3072_io_s),
    .io_co(FullAdder_3072_io_co)
  );
  FullAdder FullAdder_3073 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3073_io_a),
    .io_b(FullAdder_3073_io_b),
    .io_ci(FullAdder_3073_io_ci),
    .io_s(FullAdder_3073_io_s),
    .io_co(FullAdder_3073_io_co)
  );
  FullAdder FullAdder_3074 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3074_io_a),
    .io_b(FullAdder_3074_io_b),
    .io_ci(FullAdder_3074_io_ci),
    .io_s(FullAdder_3074_io_s),
    .io_co(FullAdder_3074_io_co)
  );
  FullAdder FullAdder_3075 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3075_io_a),
    .io_b(FullAdder_3075_io_b),
    .io_ci(FullAdder_3075_io_ci),
    .io_s(FullAdder_3075_io_s),
    .io_co(FullAdder_3075_io_co)
  );
  FullAdder FullAdder_3076 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3076_io_a),
    .io_b(FullAdder_3076_io_b),
    .io_ci(FullAdder_3076_io_ci),
    .io_s(FullAdder_3076_io_s),
    .io_co(FullAdder_3076_io_co)
  );
  HalfAdder HalfAdder_106 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_106_io_a),
    .io_b(HalfAdder_106_io_b),
    .io_s(HalfAdder_106_io_s),
    .io_co(HalfAdder_106_io_co)
  );
  FullAdder FullAdder_3077 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3077_io_a),
    .io_b(FullAdder_3077_io_b),
    .io_ci(FullAdder_3077_io_ci),
    .io_s(FullAdder_3077_io_s),
    .io_co(FullAdder_3077_io_co)
  );
  FullAdder FullAdder_3078 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3078_io_a),
    .io_b(FullAdder_3078_io_b),
    .io_ci(FullAdder_3078_io_ci),
    .io_s(FullAdder_3078_io_s),
    .io_co(FullAdder_3078_io_co)
  );
  FullAdder FullAdder_3079 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3079_io_a),
    .io_b(FullAdder_3079_io_b),
    .io_ci(FullAdder_3079_io_ci),
    .io_s(FullAdder_3079_io_s),
    .io_co(FullAdder_3079_io_co)
  );
  FullAdder FullAdder_3080 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3080_io_a),
    .io_b(FullAdder_3080_io_b),
    .io_ci(FullAdder_3080_io_ci),
    .io_s(FullAdder_3080_io_s),
    .io_co(FullAdder_3080_io_co)
  );
  FullAdder FullAdder_3081 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3081_io_a),
    .io_b(FullAdder_3081_io_b),
    .io_ci(FullAdder_3081_io_ci),
    .io_s(FullAdder_3081_io_s),
    .io_co(FullAdder_3081_io_co)
  );
  FullAdder FullAdder_3082 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3082_io_a),
    .io_b(FullAdder_3082_io_b),
    .io_ci(FullAdder_3082_io_ci),
    .io_s(FullAdder_3082_io_s),
    .io_co(FullAdder_3082_io_co)
  );
  FullAdder FullAdder_3083 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3083_io_a),
    .io_b(FullAdder_3083_io_b),
    .io_ci(FullAdder_3083_io_ci),
    .io_s(FullAdder_3083_io_s),
    .io_co(FullAdder_3083_io_co)
  );
  FullAdder FullAdder_3084 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3084_io_a),
    .io_b(FullAdder_3084_io_b),
    .io_ci(FullAdder_3084_io_ci),
    .io_s(FullAdder_3084_io_s),
    .io_co(FullAdder_3084_io_co)
  );
  FullAdder FullAdder_3085 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3085_io_a),
    .io_b(FullAdder_3085_io_b),
    .io_ci(FullAdder_3085_io_ci),
    .io_s(FullAdder_3085_io_s),
    .io_co(FullAdder_3085_io_co)
  );
  FullAdder FullAdder_3086 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3086_io_a),
    .io_b(FullAdder_3086_io_b),
    .io_ci(FullAdder_3086_io_ci),
    .io_s(FullAdder_3086_io_s),
    .io_co(FullAdder_3086_io_co)
  );
  FullAdder FullAdder_3087 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3087_io_a),
    .io_b(FullAdder_3087_io_b),
    .io_ci(FullAdder_3087_io_ci),
    .io_s(FullAdder_3087_io_s),
    .io_co(FullAdder_3087_io_co)
  );
  FullAdder FullAdder_3088 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3088_io_a),
    .io_b(FullAdder_3088_io_b),
    .io_ci(FullAdder_3088_io_ci),
    .io_s(FullAdder_3088_io_s),
    .io_co(FullAdder_3088_io_co)
  );
  FullAdder FullAdder_3089 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3089_io_a),
    .io_b(FullAdder_3089_io_b),
    .io_ci(FullAdder_3089_io_ci),
    .io_s(FullAdder_3089_io_s),
    .io_co(FullAdder_3089_io_co)
  );
  FullAdder FullAdder_3090 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3090_io_a),
    .io_b(FullAdder_3090_io_b),
    .io_ci(FullAdder_3090_io_ci),
    .io_s(FullAdder_3090_io_s),
    .io_co(FullAdder_3090_io_co)
  );
  FullAdder FullAdder_3091 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3091_io_a),
    .io_b(FullAdder_3091_io_b),
    .io_ci(FullAdder_3091_io_ci),
    .io_s(FullAdder_3091_io_s),
    .io_co(FullAdder_3091_io_co)
  );
  FullAdder FullAdder_3092 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3092_io_a),
    .io_b(FullAdder_3092_io_b),
    .io_ci(FullAdder_3092_io_ci),
    .io_s(FullAdder_3092_io_s),
    .io_co(FullAdder_3092_io_co)
  );
  FullAdder FullAdder_3093 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3093_io_a),
    .io_b(FullAdder_3093_io_b),
    .io_ci(FullAdder_3093_io_ci),
    .io_s(FullAdder_3093_io_s),
    .io_co(FullAdder_3093_io_co)
  );
  FullAdder FullAdder_3094 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3094_io_a),
    .io_b(FullAdder_3094_io_b),
    .io_ci(FullAdder_3094_io_ci),
    .io_s(FullAdder_3094_io_s),
    .io_co(FullAdder_3094_io_co)
  );
  FullAdder FullAdder_3095 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3095_io_a),
    .io_b(FullAdder_3095_io_b),
    .io_ci(FullAdder_3095_io_ci),
    .io_s(FullAdder_3095_io_s),
    .io_co(FullAdder_3095_io_co)
  );
  FullAdder FullAdder_3096 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3096_io_a),
    .io_b(FullAdder_3096_io_b),
    .io_ci(FullAdder_3096_io_ci),
    .io_s(FullAdder_3096_io_s),
    .io_co(FullAdder_3096_io_co)
  );
  FullAdder FullAdder_3097 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3097_io_a),
    .io_b(FullAdder_3097_io_b),
    .io_ci(FullAdder_3097_io_ci),
    .io_s(FullAdder_3097_io_s),
    .io_co(FullAdder_3097_io_co)
  );
  FullAdder FullAdder_3098 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3098_io_a),
    .io_b(FullAdder_3098_io_b),
    .io_ci(FullAdder_3098_io_ci),
    .io_s(FullAdder_3098_io_s),
    .io_co(FullAdder_3098_io_co)
  );
  FullAdder FullAdder_3099 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3099_io_a),
    .io_b(FullAdder_3099_io_b),
    .io_ci(FullAdder_3099_io_ci),
    .io_s(FullAdder_3099_io_s),
    .io_co(FullAdder_3099_io_co)
  );
  FullAdder FullAdder_3100 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3100_io_a),
    .io_b(FullAdder_3100_io_b),
    .io_ci(FullAdder_3100_io_ci),
    .io_s(FullAdder_3100_io_s),
    .io_co(FullAdder_3100_io_co)
  );
  FullAdder FullAdder_3101 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3101_io_a),
    .io_b(FullAdder_3101_io_b),
    .io_ci(FullAdder_3101_io_ci),
    .io_s(FullAdder_3101_io_s),
    .io_co(FullAdder_3101_io_co)
  );
  FullAdder FullAdder_3102 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3102_io_a),
    .io_b(FullAdder_3102_io_b),
    .io_ci(FullAdder_3102_io_ci),
    .io_s(FullAdder_3102_io_s),
    .io_co(FullAdder_3102_io_co)
  );
  FullAdder FullAdder_3103 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3103_io_a),
    .io_b(FullAdder_3103_io_b),
    .io_ci(FullAdder_3103_io_ci),
    .io_s(FullAdder_3103_io_s),
    .io_co(FullAdder_3103_io_co)
  );
  FullAdder FullAdder_3104 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3104_io_a),
    .io_b(FullAdder_3104_io_b),
    .io_ci(FullAdder_3104_io_ci),
    .io_s(FullAdder_3104_io_s),
    .io_co(FullAdder_3104_io_co)
  );
  FullAdder FullAdder_3105 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3105_io_a),
    .io_b(FullAdder_3105_io_b),
    .io_ci(FullAdder_3105_io_ci),
    .io_s(FullAdder_3105_io_s),
    .io_co(FullAdder_3105_io_co)
  );
  FullAdder FullAdder_3106 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3106_io_a),
    .io_b(FullAdder_3106_io_b),
    .io_ci(FullAdder_3106_io_ci),
    .io_s(FullAdder_3106_io_s),
    .io_co(FullAdder_3106_io_co)
  );
  FullAdder FullAdder_3107 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3107_io_a),
    .io_b(FullAdder_3107_io_b),
    .io_ci(FullAdder_3107_io_ci),
    .io_s(FullAdder_3107_io_s),
    .io_co(FullAdder_3107_io_co)
  );
  FullAdder FullAdder_3108 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3108_io_a),
    .io_b(FullAdder_3108_io_b),
    .io_ci(FullAdder_3108_io_ci),
    .io_s(FullAdder_3108_io_s),
    .io_co(FullAdder_3108_io_co)
  );
  FullAdder FullAdder_3109 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3109_io_a),
    .io_b(FullAdder_3109_io_b),
    .io_ci(FullAdder_3109_io_ci),
    .io_s(FullAdder_3109_io_s),
    .io_co(FullAdder_3109_io_co)
  );
  FullAdder FullAdder_3110 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3110_io_a),
    .io_b(FullAdder_3110_io_b),
    .io_ci(FullAdder_3110_io_ci),
    .io_s(FullAdder_3110_io_s),
    .io_co(FullAdder_3110_io_co)
  );
  FullAdder FullAdder_3111 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3111_io_a),
    .io_b(FullAdder_3111_io_b),
    .io_ci(FullAdder_3111_io_ci),
    .io_s(FullAdder_3111_io_s),
    .io_co(FullAdder_3111_io_co)
  );
  FullAdder FullAdder_3112 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3112_io_a),
    .io_b(FullAdder_3112_io_b),
    .io_ci(FullAdder_3112_io_ci),
    .io_s(FullAdder_3112_io_s),
    .io_co(FullAdder_3112_io_co)
  );
  FullAdder FullAdder_3113 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3113_io_a),
    .io_b(FullAdder_3113_io_b),
    .io_ci(FullAdder_3113_io_ci),
    .io_s(FullAdder_3113_io_s),
    .io_co(FullAdder_3113_io_co)
  );
  FullAdder FullAdder_3114 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3114_io_a),
    .io_b(FullAdder_3114_io_b),
    .io_ci(FullAdder_3114_io_ci),
    .io_s(FullAdder_3114_io_s),
    .io_co(FullAdder_3114_io_co)
  );
  FullAdder FullAdder_3115 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3115_io_a),
    .io_b(FullAdder_3115_io_b),
    .io_ci(FullAdder_3115_io_ci),
    .io_s(FullAdder_3115_io_s),
    .io_co(FullAdder_3115_io_co)
  );
  FullAdder FullAdder_3116 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3116_io_a),
    .io_b(FullAdder_3116_io_b),
    .io_ci(FullAdder_3116_io_ci),
    .io_s(FullAdder_3116_io_s),
    .io_co(FullAdder_3116_io_co)
  );
  FullAdder FullAdder_3117 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3117_io_a),
    .io_b(FullAdder_3117_io_b),
    .io_ci(FullAdder_3117_io_ci),
    .io_s(FullAdder_3117_io_s),
    .io_co(FullAdder_3117_io_co)
  );
  FullAdder FullAdder_3118 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3118_io_a),
    .io_b(FullAdder_3118_io_b),
    .io_ci(FullAdder_3118_io_ci),
    .io_s(FullAdder_3118_io_s),
    .io_co(FullAdder_3118_io_co)
  );
  HalfAdder HalfAdder_107 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_107_io_a),
    .io_b(HalfAdder_107_io_b),
    .io_s(HalfAdder_107_io_s),
    .io_co(HalfAdder_107_io_co)
  );
  FullAdder FullAdder_3119 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3119_io_a),
    .io_b(FullAdder_3119_io_b),
    .io_ci(FullAdder_3119_io_ci),
    .io_s(FullAdder_3119_io_s),
    .io_co(FullAdder_3119_io_co)
  );
  FullAdder FullAdder_3120 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3120_io_a),
    .io_b(FullAdder_3120_io_b),
    .io_ci(FullAdder_3120_io_ci),
    .io_s(FullAdder_3120_io_s),
    .io_co(FullAdder_3120_io_co)
  );
  FullAdder FullAdder_3121 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3121_io_a),
    .io_b(FullAdder_3121_io_b),
    .io_ci(FullAdder_3121_io_ci),
    .io_s(FullAdder_3121_io_s),
    .io_co(FullAdder_3121_io_co)
  );
  FullAdder FullAdder_3122 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3122_io_a),
    .io_b(FullAdder_3122_io_b),
    .io_ci(FullAdder_3122_io_ci),
    .io_s(FullAdder_3122_io_s),
    .io_co(FullAdder_3122_io_co)
  );
  FullAdder FullAdder_3123 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3123_io_a),
    .io_b(FullAdder_3123_io_b),
    .io_ci(FullAdder_3123_io_ci),
    .io_s(FullAdder_3123_io_s),
    .io_co(FullAdder_3123_io_co)
  );
  FullAdder FullAdder_3124 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3124_io_a),
    .io_b(FullAdder_3124_io_b),
    .io_ci(FullAdder_3124_io_ci),
    .io_s(FullAdder_3124_io_s),
    .io_co(FullAdder_3124_io_co)
  );
  FullAdder FullAdder_3125 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3125_io_a),
    .io_b(FullAdder_3125_io_b),
    .io_ci(FullAdder_3125_io_ci),
    .io_s(FullAdder_3125_io_s),
    .io_co(FullAdder_3125_io_co)
  );
  FullAdder FullAdder_3126 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3126_io_a),
    .io_b(FullAdder_3126_io_b),
    .io_ci(FullAdder_3126_io_ci),
    .io_s(FullAdder_3126_io_s),
    .io_co(FullAdder_3126_io_co)
  );
  FullAdder FullAdder_3127 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3127_io_a),
    .io_b(FullAdder_3127_io_b),
    .io_ci(FullAdder_3127_io_ci),
    .io_s(FullAdder_3127_io_s),
    .io_co(FullAdder_3127_io_co)
  );
  FullAdder FullAdder_3128 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3128_io_a),
    .io_b(FullAdder_3128_io_b),
    .io_ci(FullAdder_3128_io_ci),
    .io_s(FullAdder_3128_io_s),
    .io_co(FullAdder_3128_io_co)
  );
  FullAdder FullAdder_3129 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3129_io_a),
    .io_b(FullAdder_3129_io_b),
    .io_ci(FullAdder_3129_io_ci),
    .io_s(FullAdder_3129_io_s),
    .io_co(FullAdder_3129_io_co)
  );
  FullAdder FullAdder_3130 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3130_io_a),
    .io_b(FullAdder_3130_io_b),
    .io_ci(FullAdder_3130_io_ci),
    .io_s(FullAdder_3130_io_s),
    .io_co(FullAdder_3130_io_co)
  );
  FullAdder FullAdder_3131 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3131_io_a),
    .io_b(FullAdder_3131_io_b),
    .io_ci(FullAdder_3131_io_ci),
    .io_s(FullAdder_3131_io_s),
    .io_co(FullAdder_3131_io_co)
  );
  FullAdder FullAdder_3132 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3132_io_a),
    .io_b(FullAdder_3132_io_b),
    .io_ci(FullAdder_3132_io_ci),
    .io_s(FullAdder_3132_io_s),
    .io_co(FullAdder_3132_io_co)
  );
  FullAdder FullAdder_3133 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3133_io_a),
    .io_b(FullAdder_3133_io_b),
    .io_ci(FullAdder_3133_io_ci),
    .io_s(FullAdder_3133_io_s),
    .io_co(FullAdder_3133_io_co)
  );
  FullAdder FullAdder_3134 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3134_io_a),
    .io_b(FullAdder_3134_io_b),
    .io_ci(FullAdder_3134_io_ci),
    .io_s(FullAdder_3134_io_s),
    .io_co(FullAdder_3134_io_co)
  );
  FullAdder FullAdder_3135 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3135_io_a),
    .io_b(FullAdder_3135_io_b),
    .io_ci(FullAdder_3135_io_ci),
    .io_s(FullAdder_3135_io_s),
    .io_co(FullAdder_3135_io_co)
  );
  FullAdder FullAdder_3136 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3136_io_a),
    .io_b(FullAdder_3136_io_b),
    .io_ci(FullAdder_3136_io_ci),
    .io_s(FullAdder_3136_io_s),
    .io_co(FullAdder_3136_io_co)
  );
  FullAdder FullAdder_3137 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3137_io_a),
    .io_b(FullAdder_3137_io_b),
    .io_ci(FullAdder_3137_io_ci),
    .io_s(FullAdder_3137_io_s),
    .io_co(FullAdder_3137_io_co)
  );
  FullAdder FullAdder_3138 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3138_io_a),
    .io_b(FullAdder_3138_io_b),
    .io_ci(FullAdder_3138_io_ci),
    .io_s(FullAdder_3138_io_s),
    .io_co(FullAdder_3138_io_co)
  );
  FullAdder FullAdder_3139 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3139_io_a),
    .io_b(FullAdder_3139_io_b),
    .io_ci(FullAdder_3139_io_ci),
    .io_s(FullAdder_3139_io_s),
    .io_co(FullAdder_3139_io_co)
  );
  FullAdder FullAdder_3140 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3140_io_a),
    .io_b(FullAdder_3140_io_b),
    .io_ci(FullAdder_3140_io_ci),
    .io_s(FullAdder_3140_io_s),
    .io_co(FullAdder_3140_io_co)
  );
  FullAdder FullAdder_3141 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3141_io_a),
    .io_b(FullAdder_3141_io_b),
    .io_ci(FullAdder_3141_io_ci),
    .io_s(FullAdder_3141_io_s),
    .io_co(FullAdder_3141_io_co)
  );
  FullAdder FullAdder_3142 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3142_io_a),
    .io_b(FullAdder_3142_io_b),
    .io_ci(FullAdder_3142_io_ci),
    .io_s(FullAdder_3142_io_s),
    .io_co(FullAdder_3142_io_co)
  );
  FullAdder FullAdder_3143 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3143_io_a),
    .io_b(FullAdder_3143_io_b),
    .io_ci(FullAdder_3143_io_ci),
    .io_s(FullAdder_3143_io_s),
    .io_co(FullAdder_3143_io_co)
  );
  FullAdder FullAdder_3144 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3144_io_a),
    .io_b(FullAdder_3144_io_b),
    .io_ci(FullAdder_3144_io_ci),
    .io_s(FullAdder_3144_io_s),
    .io_co(FullAdder_3144_io_co)
  );
  FullAdder FullAdder_3145 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3145_io_a),
    .io_b(FullAdder_3145_io_b),
    .io_ci(FullAdder_3145_io_ci),
    .io_s(FullAdder_3145_io_s),
    .io_co(FullAdder_3145_io_co)
  );
  FullAdder FullAdder_3146 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3146_io_a),
    .io_b(FullAdder_3146_io_b),
    .io_ci(FullAdder_3146_io_ci),
    .io_s(FullAdder_3146_io_s),
    .io_co(FullAdder_3146_io_co)
  );
  FullAdder FullAdder_3147 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3147_io_a),
    .io_b(FullAdder_3147_io_b),
    .io_ci(FullAdder_3147_io_ci),
    .io_s(FullAdder_3147_io_s),
    .io_co(FullAdder_3147_io_co)
  );
  FullAdder FullAdder_3148 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3148_io_a),
    .io_b(FullAdder_3148_io_b),
    .io_ci(FullAdder_3148_io_ci),
    .io_s(FullAdder_3148_io_s),
    .io_co(FullAdder_3148_io_co)
  );
  FullAdder FullAdder_3149 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3149_io_a),
    .io_b(FullAdder_3149_io_b),
    .io_ci(FullAdder_3149_io_ci),
    .io_s(FullAdder_3149_io_s),
    .io_co(FullAdder_3149_io_co)
  );
  FullAdder FullAdder_3150 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3150_io_a),
    .io_b(FullAdder_3150_io_b),
    .io_ci(FullAdder_3150_io_ci),
    .io_s(FullAdder_3150_io_s),
    .io_co(FullAdder_3150_io_co)
  );
  FullAdder FullAdder_3151 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3151_io_a),
    .io_b(FullAdder_3151_io_b),
    .io_ci(FullAdder_3151_io_ci),
    .io_s(FullAdder_3151_io_s),
    .io_co(FullAdder_3151_io_co)
  );
  FullAdder FullAdder_3152 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3152_io_a),
    .io_b(FullAdder_3152_io_b),
    .io_ci(FullAdder_3152_io_ci),
    .io_s(FullAdder_3152_io_s),
    .io_co(FullAdder_3152_io_co)
  );
  FullAdder FullAdder_3153 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3153_io_a),
    .io_b(FullAdder_3153_io_b),
    .io_ci(FullAdder_3153_io_ci),
    .io_s(FullAdder_3153_io_s),
    .io_co(FullAdder_3153_io_co)
  );
  FullAdder FullAdder_3154 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3154_io_a),
    .io_b(FullAdder_3154_io_b),
    .io_ci(FullAdder_3154_io_ci),
    .io_s(FullAdder_3154_io_s),
    .io_co(FullAdder_3154_io_co)
  );
  FullAdder FullAdder_3155 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3155_io_a),
    .io_b(FullAdder_3155_io_b),
    .io_ci(FullAdder_3155_io_ci),
    .io_s(FullAdder_3155_io_s),
    .io_co(FullAdder_3155_io_co)
  );
  FullAdder FullAdder_3156 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3156_io_a),
    .io_b(FullAdder_3156_io_b),
    .io_ci(FullAdder_3156_io_ci),
    .io_s(FullAdder_3156_io_s),
    .io_co(FullAdder_3156_io_co)
  );
  FullAdder FullAdder_3157 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3157_io_a),
    .io_b(FullAdder_3157_io_b),
    .io_ci(FullAdder_3157_io_ci),
    .io_s(FullAdder_3157_io_s),
    .io_co(FullAdder_3157_io_co)
  );
  FullAdder FullAdder_3158 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3158_io_a),
    .io_b(FullAdder_3158_io_b),
    .io_ci(FullAdder_3158_io_ci),
    .io_s(FullAdder_3158_io_s),
    .io_co(FullAdder_3158_io_co)
  );
  FullAdder FullAdder_3159 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3159_io_a),
    .io_b(FullAdder_3159_io_b),
    .io_ci(FullAdder_3159_io_ci),
    .io_s(FullAdder_3159_io_s),
    .io_co(FullAdder_3159_io_co)
  );
  FullAdder FullAdder_3160 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3160_io_a),
    .io_b(FullAdder_3160_io_b),
    .io_ci(FullAdder_3160_io_ci),
    .io_s(FullAdder_3160_io_s),
    .io_co(FullAdder_3160_io_co)
  );
  FullAdder FullAdder_3161 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3161_io_a),
    .io_b(FullAdder_3161_io_b),
    .io_ci(FullAdder_3161_io_ci),
    .io_s(FullAdder_3161_io_s),
    .io_co(FullAdder_3161_io_co)
  );
  FullAdder FullAdder_3162 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3162_io_a),
    .io_b(FullAdder_3162_io_b),
    .io_ci(FullAdder_3162_io_ci),
    .io_s(FullAdder_3162_io_s),
    .io_co(FullAdder_3162_io_co)
  );
  FullAdder FullAdder_3163 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3163_io_a),
    .io_b(FullAdder_3163_io_b),
    .io_ci(FullAdder_3163_io_ci),
    .io_s(FullAdder_3163_io_s),
    .io_co(FullAdder_3163_io_co)
  );
  FullAdder FullAdder_3164 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3164_io_a),
    .io_b(FullAdder_3164_io_b),
    .io_ci(FullAdder_3164_io_ci),
    .io_s(FullAdder_3164_io_s),
    .io_co(FullAdder_3164_io_co)
  );
  FullAdder FullAdder_3165 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3165_io_a),
    .io_b(FullAdder_3165_io_b),
    .io_ci(FullAdder_3165_io_ci),
    .io_s(FullAdder_3165_io_s),
    .io_co(FullAdder_3165_io_co)
  );
  FullAdder FullAdder_3166 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3166_io_a),
    .io_b(FullAdder_3166_io_b),
    .io_ci(FullAdder_3166_io_ci),
    .io_s(FullAdder_3166_io_s),
    .io_co(FullAdder_3166_io_co)
  );
  FullAdder FullAdder_3167 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3167_io_a),
    .io_b(FullAdder_3167_io_b),
    .io_ci(FullAdder_3167_io_ci),
    .io_s(FullAdder_3167_io_s),
    .io_co(FullAdder_3167_io_co)
  );
  HalfAdder HalfAdder_108 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_108_io_a),
    .io_b(HalfAdder_108_io_b),
    .io_s(HalfAdder_108_io_s),
    .io_co(HalfAdder_108_io_co)
  );
  FullAdder FullAdder_3168 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3168_io_a),
    .io_b(FullAdder_3168_io_b),
    .io_ci(FullAdder_3168_io_ci),
    .io_s(FullAdder_3168_io_s),
    .io_co(FullAdder_3168_io_co)
  );
  FullAdder FullAdder_3169 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3169_io_a),
    .io_b(FullAdder_3169_io_b),
    .io_ci(FullAdder_3169_io_ci),
    .io_s(FullAdder_3169_io_s),
    .io_co(FullAdder_3169_io_co)
  );
  HalfAdder HalfAdder_109 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_109_io_a),
    .io_b(HalfAdder_109_io_b),
    .io_s(HalfAdder_109_io_s),
    .io_co(HalfAdder_109_io_co)
  );
  FullAdder FullAdder_3170 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3170_io_a),
    .io_b(FullAdder_3170_io_b),
    .io_ci(FullAdder_3170_io_ci),
    .io_s(FullAdder_3170_io_s),
    .io_co(FullAdder_3170_io_co)
  );
  FullAdder FullAdder_3171 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3171_io_a),
    .io_b(FullAdder_3171_io_b),
    .io_ci(FullAdder_3171_io_ci),
    .io_s(FullAdder_3171_io_s),
    .io_co(FullAdder_3171_io_co)
  );
  FullAdder FullAdder_3172 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3172_io_a),
    .io_b(FullAdder_3172_io_b),
    .io_ci(FullAdder_3172_io_ci),
    .io_s(FullAdder_3172_io_s),
    .io_co(FullAdder_3172_io_co)
  );
  HalfAdder HalfAdder_110 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_110_io_a),
    .io_b(HalfAdder_110_io_b),
    .io_s(HalfAdder_110_io_s),
    .io_co(HalfAdder_110_io_co)
  );
  HalfAdder HalfAdder_111 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_111_io_a),
    .io_b(HalfAdder_111_io_b),
    .io_s(HalfAdder_111_io_s),
    .io_co(HalfAdder_111_io_co)
  );
  FullAdder FullAdder_3173 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3173_io_a),
    .io_b(FullAdder_3173_io_b),
    .io_ci(FullAdder_3173_io_ci),
    .io_s(FullAdder_3173_io_s),
    .io_co(FullAdder_3173_io_co)
  );
  FullAdder FullAdder_3174 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3174_io_a),
    .io_b(FullAdder_3174_io_b),
    .io_ci(FullAdder_3174_io_ci),
    .io_s(FullAdder_3174_io_s),
    .io_co(FullAdder_3174_io_co)
  );
  FullAdder FullAdder_3175 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3175_io_a),
    .io_b(FullAdder_3175_io_b),
    .io_ci(FullAdder_3175_io_ci),
    .io_s(FullAdder_3175_io_s),
    .io_co(FullAdder_3175_io_co)
  );
  HalfAdder HalfAdder_112 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_112_io_a),
    .io_b(HalfAdder_112_io_b),
    .io_s(HalfAdder_112_io_s),
    .io_co(HalfAdder_112_io_co)
  );
  HalfAdder HalfAdder_113 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_113_io_a),
    .io_b(HalfAdder_113_io_b),
    .io_s(HalfAdder_113_io_s),
    .io_co(HalfAdder_113_io_co)
  );
  HalfAdder HalfAdder_114 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_114_io_a),
    .io_b(HalfAdder_114_io_b),
    .io_s(HalfAdder_114_io_s),
    .io_co(HalfAdder_114_io_co)
  );
  HalfAdder HalfAdder_115 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_115_io_a),
    .io_b(HalfAdder_115_io_b),
    .io_s(HalfAdder_115_io_s),
    .io_co(HalfAdder_115_io_co)
  );
  FullAdder FullAdder_3176 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3176_io_a),
    .io_b(FullAdder_3176_io_b),
    .io_ci(FullAdder_3176_io_ci),
    .io_s(FullAdder_3176_io_s),
    .io_co(FullAdder_3176_io_co)
  );
  HalfAdder HalfAdder_116 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_116_io_a),
    .io_b(HalfAdder_116_io_b),
    .io_s(HalfAdder_116_io_s),
    .io_co(HalfAdder_116_io_co)
  );
  HalfAdder HalfAdder_117 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_117_io_a),
    .io_b(HalfAdder_117_io_b),
    .io_s(HalfAdder_117_io_s),
    .io_co(HalfAdder_117_io_co)
  );
  FullAdder FullAdder_3177 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3177_io_a),
    .io_b(FullAdder_3177_io_b),
    .io_ci(FullAdder_3177_io_ci),
    .io_s(FullAdder_3177_io_s),
    .io_co(FullAdder_3177_io_co)
  );
  HalfAdder HalfAdder_118 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_118_io_a),
    .io_b(HalfAdder_118_io_b),
    .io_s(HalfAdder_118_io_s),
    .io_co(HalfAdder_118_io_co)
  );
  HalfAdder HalfAdder_119 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_119_io_a),
    .io_b(HalfAdder_119_io_b),
    .io_s(HalfAdder_119_io_s),
    .io_co(HalfAdder_119_io_co)
  );
  FullAdder FullAdder_3178 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3178_io_a),
    .io_b(FullAdder_3178_io_b),
    .io_ci(FullAdder_3178_io_ci),
    .io_s(FullAdder_3178_io_s),
    .io_co(FullAdder_3178_io_co)
  );
  FullAdder FullAdder_3179 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3179_io_a),
    .io_b(FullAdder_3179_io_b),
    .io_ci(FullAdder_3179_io_ci),
    .io_s(FullAdder_3179_io_s),
    .io_co(FullAdder_3179_io_co)
  );
  FullAdder FullAdder_3180 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3180_io_a),
    .io_b(FullAdder_3180_io_b),
    .io_ci(FullAdder_3180_io_ci),
    .io_s(FullAdder_3180_io_s),
    .io_co(FullAdder_3180_io_co)
  );
  FullAdder FullAdder_3181 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3181_io_a),
    .io_b(FullAdder_3181_io_b),
    .io_ci(FullAdder_3181_io_ci),
    .io_s(FullAdder_3181_io_s),
    .io_co(FullAdder_3181_io_co)
  );
  FullAdder FullAdder_3182 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3182_io_a),
    .io_b(FullAdder_3182_io_b),
    .io_ci(FullAdder_3182_io_ci),
    .io_s(FullAdder_3182_io_s),
    .io_co(FullAdder_3182_io_co)
  );
  FullAdder FullAdder_3183 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3183_io_a),
    .io_b(FullAdder_3183_io_b),
    .io_ci(FullAdder_3183_io_ci),
    .io_s(FullAdder_3183_io_s),
    .io_co(FullAdder_3183_io_co)
  );
  FullAdder FullAdder_3184 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3184_io_a),
    .io_b(FullAdder_3184_io_b),
    .io_ci(FullAdder_3184_io_ci),
    .io_s(FullAdder_3184_io_s),
    .io_co(FullAdder_3184_io_co)
  );
  FullAdder FullAdder_3185 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3185_io_a),
    .io_b(FullAdder_3185_io_b),
    .io_ci(FullAdder_3185_io_ci),
    .io_s(FullAdder_3185_io_s),
    .io_co(FullAdder_3185_io_co)
  );
  FullAdder FullAdder_3186 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3186_io_a),
    .io_b(FullAdder_3186_io_b),
    .io_ci(FullAdder_3186_io_ci),
    .io_s(FullAdder_3186_io_s),
    .io_co(FullAdder_3186_io_co)
  );
  FullAdder FullAdder_3187 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3187_io_a),
    .io_b(FullAdder_3187_io_b),
    .io_ci(FullAdder_3187_io_ci),
    .io_s(FullAdder_3187_io_s),
    .io_co(FullAdder_3187_io_co)
  );
  FullAdder FullAdder_3188 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3188_io_a),
    .io_b(FullAdder_3188_io_b),
    .io_ci(FullAdder_3188_io_ci),
    .io_s(FullAdder_3188_io_s),
    .io_co(FullAdder_3188_io_co)
  );
  HalfAdder HalfAdder_120 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_120_io_a),
    .io_b(HalfAdder_120_io_b),
    .io_s(HalfAdder_120_io_s),
    .io_co(HalfAdder_120_io_co)
  );
  FullAdder FullAdder_3189 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3189_io_a),
    .io_b(FullAdder_3189_io_b),
    .io_ci(FullAdder_3189_io_ci),
    .io_s(FullAdder_3189_io_s),
    .io_co(FullAdder_3189_io_co)
  );
  HalfAdder HalfAdder_121 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_121_io_a),
    .io_b(HalfAdder_121_io_b),
    .io_s(HalfAdder_121_io_s),
    .io_co(HalfAdder_121_io_co)
  );
  FullAdder FullAdder_3190 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3190_io_a),
    .io_b(FullAdder_3190_io_b),
    .io_ci(FullAdder_3190_io_ci),
    .io_s(FullAdder_3190_io_s),
    .io_co(FullAdder_3190_io_co)
  );
  FullAdder FullAdder_3191 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3191_io_a),
    .io_b(FullAdder_3191_io_b),
    .io_ci(FullAdder_3191_io_ci),
    .io_s(FullAdder_3191_io_s),
    .io_co(FullAdder_3191_io_co)
  );
  FullAdder FullAdder_3192 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3192_io_a),
    .io_b(FullAdder_3192_io_b),
    .io_ci(FullAdder_3192_io_ci),
    .io_s(FullAdder_3192_io_s),
    .io_co(FullAdder_3192_io_co)
  );
  FullAdder FullAdder_3193 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3193_io_a),
    .io_b(FullAdder_3193_io_b),
    .io_ci(FullAdder_3193_io_ci),
    .io_s(FullAdder_3193_io_s),
    .io_co(FullAdder_3193_io_co)
  );
  FullAdder FullAdder_3194 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3194_io_a),
    .io_b(FullAdder_3194_io_b),
    .io_ci(FullAdder_3194_io_ci),
    .io_s(FullAdder_3194_io_s),
    .io_co(FullAdder_3194_io_co)
  );
  FullAdder FullAdder_3195 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3195_io_a),
    .io_b(FullAdder_3195_io_b),
    .io_ci(FullAdder_3195_io_ci),
    .io_s(FullAdder_3195_io_s),
    .io_co(FullAdder_3195_io_co)
  );
  FullAdder FullAdder_3196 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3196_io_a),
    .io_b(FullAdder_3196_io_b),
    .io_ci(FullAdder_3196_io_ci),
    .io_s(FullAdder_3196_io_s),
    .io_co(FullAdder_3196_io_co)
  );
  FullAdder FullAdder_3197 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3197_io_a),
    .io_b(FullAdder_3197_io_b),
    .io_ci(FullAdder_3197_io_ci),
    .io_s(FullAdder_3197_io_s),
    .io_co(FullAdder_3197_io_co)
  );
  FullAdder FullAdder_3198 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3198_io_a),
    .io_b(FullAdder_3198_io_b),
    .io_ci(FullAdder_3198_io_ci),
    .io_s(FullAdder_3198_io_s),
    .io_co(FullAdder_3198_io_co)
  );
  FullAdder FullAdder_3199 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3199_io_a),
    .io_b(FullAdder_3199_io_b),
    .io_ci(FullAdder_3199_io_ci),
    .io_s(FullAdder_3199_io_s),
    .io_co(FullAdder_3199_io_co)
  );
  FullAdder FullAdder_3200 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3200_io_a),
    .io_b(FullAdder_3200_io_b),
    .io_ci(FullAdder_3200_io_ci),
    .io_s(FullAdder_3200_io_s),
    .io_co(FullAdder_3200_io_co)
  );
  FullAdder FullAdder_3201 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3201_io_a),
    .io_b(FullAdder_3201_io_b),
    .io_ci(FullAdder_3201_io_ci),
    .io_s(FullAdder_3201_io_s),
    .io_co(FullAdder_3201_io_co)
  );
  FullAdder FullAdder_3202 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3202_io_a),
    .io_b(FullAdder_3202_io_b),
    .io_ci(FullAdder_3202_io_ci),
    .io_s(FullAdder_3202_io_s),
    .io_co(FullAdder_3202_io_co)
  );
  FullAdder FullAdder_3203 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3203_io_a),
    .io_b(FullAdder_3203_io_b),
    .io_ci(FullAdder_3203_io_ci),
    .io_s(FullAdder_3203_io_s),
    .io_co(FullAdder_3203_io_co)
  );
  FullAdder FullAdder_3204 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3204_io_a),
    .io_b(FullAdder_3204_io_b),
    .io_ci(FullAdder_3204_io_ci),
    .io_s(FullAdder_3204_io_s),
    .io_co(FullAdder_3204_io_co)
  );
  FullAdder FullAdder_3205 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3205_io_a),
    .io_b(FullAdder_3205_io_b),
    .io_ci(FullAdder_3205_io_ci),
    .io_s(FullAdder_3205_io_s),
    .io_co(FullAdder_3205_io_co)
  );
  FullAdder FullAdder_3206 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3206_io_a),
    .io_b(FullAdder_3206_io_b),
    .io_ci(FullAdder_3206_io_ci),
    .io_s(FullAdder_3206_io_s),
    .io_co(FullAdder_3206_io_co)
  );
  FullAdder FullAdder_3207 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3207_io_a),
    .io_b(FullAdder_3207_io_b),
    .io_ci(FullAdder_3207_io_ci),
    .io_s(FullAdder_3207_io_s),
    .io_co(FullAdder_3207_io_co)
  );
  FullAdder FullAdder_3208 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3208_io_a),
    .io_b(FullAdder_3208_io_b),
    .io_ci(FullAdder_3208_io_ci),
    .io_s(FullAdder_3208_io_s),
    .io_co(FullAdder_3208_io_co)
  );
  FullAdder FullAdder_3209 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3209_io_a),
    .io_b(FullAdder_3209_io_b),
    .io_ci(FullAdder_3209_io_ci),
    .io_s(FullAdder_3209_io_s),
    .io_co(FullAdder_3209_io_co)
  );
  FullAdder FullAdder_3210 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3210_io_a),
    .io_b(FullAdder_3210_io_b),
    .io_ci(FullAdder_3210_io_ci),
    .io_s(FullAdder_3210_io_s),
    .io_co(FullAdder_3210_io_co)
  );
  FullAdder FullAdder_3211 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3211_io_a),
    .io_b(FullAdder_3211_io_b),
    .io_ci(FullAdder_3211_io_ci),
    .io_s(FullAdder_3211_io_s),
    .io_co(FullAdder_3211_io_co)
  );
  FullAdder FullAdder_3212 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3212_io_a),
    .io_b(FullAdder_3212_io_b),
    .io_ci(FullAdder_3212_io_ci),
    .io_s(FullAdder_3212_io_s),
    .io_co(FullAdder_3212_io_co)
  );
  FullAdder FullAdder_3213 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3213_io_a),
    .io_b(FullAdder_3213_io_b),
    .io_ci(FullAdder_3213_io_ci),
    .io_s(FullAdder_3213_io_s),
    .io_co(FullAdder_3213_io_co)
  );
  FullAdder FullAdder_3214 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3214_io_a),
    .io_b(FullAdder_3214_io_b),
    .io_ci(FullAdder_3214_io_ci),
    .io_s(FullAdder_3214_io_s),
    .io_co(FullAdder_3214_io_co)
  );
  HalfAdder HalfAdder_122 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_122_io_a),
    .io_b(HalfAdder_122_io_b),
    .io_s(HalfAdder_122_io_s),
    .io_co(HalfAdder_122_io_co)
  );
  FullAdder FullAdder_3215 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3215_io_a),
    .io_b(FullAdder_3215_io_b),
    .io_ci(FullAdder_3215_io_ci),
    .io_s(FullAdder_3215_io_s),
    .io_co(FullAdder_3215_io_co)
  );
  FullAdder FullAdder_3216 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3216_io_a),
    .io_b(FullAdder_3216_io_b),
    .io_ci(FullAdder_3216_io_ci),
    .io_s(FullAdder_3216_io_s),
    .io_co(FullAdder_3216_io_co)
  );
  HalfAdder HalfAdder_123 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_123_io_a),
    .io_b(HalfAdder_123_io_b),
    .io_s(HalfAdder_123_io_s),
    .io_co(HalfAdder_123_io_co)
  );
  FullAdder FullAdder_3217 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3217_io_a),
    .io_b(FullAdder_3217_io_b),
    .io_ci(FullAdder_3217_io_ci),
    .io_s(FullAdder_3217_io_s),
    .io_co(FullAdder_3217_io_co)
  );
  FullAdder FullAdder_3218 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3218_io_a),
    .io_b(FullAdder_3218_io_b),
    .io_ci(FullAdder_3218_io_ci),
    .io_s(FullAdder_3218_io_s),
    .io_co(FullAdder_3218_io_co)
  );
  HalfAdder HalfAdder_124 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_124_io_a),
    .io_b(HalfAdder_124_io_b),
    .io_s(HalfAdder_124_io_s),
    .io_co(HalfAdder_124_io_co)
  );
  FullAdder FullAdder_3219 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3219_io_a),
    .io_b(FullAdder_3219_io_b),
    .io_ci(FullAdder_3219_io_ci),
    .io_s(FullAdder_3219_io_s),
    .io_co(FullAdder_3219_io_co)
  );
  FullAdder FullAdder_3220 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3220_io_a),
    .io_b(FullAdder_3220_io_b),
    .io_ci(FullAdder_3220_io_ci),
    .io_s(FullAdder_3220_io_s),
    .io_co(FullAdder_3220_io_co)
  );
  FullAdder FullAdder_3221 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3221_io_a),
    .io_b(FullAdder_3221_io_b),
    .io_ci(FullAdder_3221_io_ci),
    .io_s(FullAdder_3221_io_s),
    .io_co(FullAdder_3221_io_co)
  );
  FullAdder FullAdder_3222 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3222_io_a),
    .io_b(FullAdder_3222_io_b),
    .io_ci(FullAdder_3222_io_ci),
    .io_s(FullAdder_3222_io_s),
    .io_co(FullAdder_3222_io_co)
  );
  FullAdder FullAdder_3223 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3223_io_a),
    .io_b(FullAdder_3223_io_b),
    .io_ci(FullAdder_3223_io_ci),
    .io_s(FullAdder_3223_io_s),
    .io_co(FullAdder_3223_io_co)
  );
  FullAdder FullAdder_3224 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3224_io_a),
    .io_b(FullAdder_3224_io_b),
    .io_ci(FullAdder_3224_io_ci),
    .io_s(FullAdder_3224_io_s),
    .io_co(FullAdder_3224_io_co)
  );
  FullAdder FullAdder_3225 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3225_io_a),
    .io_b(FullAdder_3225_io_b),
    .io_ci(FullAdder_3225_io_ci),
    .io_s(FullAdder_3225_io_s),
    .io_co(FullAdder_3225_io_co)
  );
  HalfAdder HalfAdder_125 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_125_io_a),
    .io_b(HalfAdder_125_io_b),
    .io_s(HalfAdder_125_io_s),
    .io_co(HalfAdder_125_io_co)
  );
  FullAdder FullAdder_3226 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3226_io_a),
    .io_b(FullAdder_3226_io_b),
    .io_ci(FullAdder_3226_io_ci),
    .io_s(FullAdder_3226_io_s),
    .io_co(FullAdder_3226_io_co)
  );
  FullAdder FullAdder_3227 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3227_io_a),
    .io_b(FullAdder_3227_io_b),
    .io_ci(FullAdder_3227_io_ci),
    .io_s(FullAdder_3227_io_s),
    .io_co(FullAdder_3227_io_co)
  );
  HalfAdder HalfAdder_126 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_126_io_a),
    .io_b(HalfAdder_126_io_b),
    .io_s(HalfAdder_126_io_s),
    .io_co(HalfAdder_126_io_co)
  );
  FullAdder FullAdder_3228 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3228_io_a),
    .io_b(FullAdder_3228_io_b),
    .io_ci(FullAdder_3228_io_ci),
    .io_s(FullAdder_3228_io_s),
    .io_co(FullAdder_3228_io_co)
  );
  FullAdder FullAdder_3229 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3229_io_a),
    .io_b(FullAdder_3229_io_b),
    .io_ci(FullAdder_3229_io_ci),
    .io_s(FullAdder_3229_io_s),
    .io_co(FullAdder_3229_io_co)
  );
  FullAdder FullAdder_3230 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3230_io_a),
    .io_b(FullAdder_3230_io_b),
    .io_ci(FullAdder_3230_io_ci),
    .io_s(FullAdder_3230_io_s),
    .io_co(FullAdder_3230_io_co)
  );
  FullAdder FullAdder_3231 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3231_io_a),
    .io_b(FullAdder_3231_io_b),
    .io_ci(FullAdder_3231_io_ci),
    .io_s(FullAdder_3231_io_s),
    .io_co(FullAdder_3231_io_co)
  );
  FullAdder FullAdder_3232 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3232_io_a),
    .io_b(FullAdder_3232_io_b),
    .io_ci(FullAdder_3232_io_ci),
    .io_s(FullAdder_3232_io_s),
    .io_co(FullAdder_3232_io_co)
  );
  FullAdder FullAdder_3233 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3233_io_a),
    .io_b(FullAdder_3233_io_b),
    .io_ci(FullAdder_3233_io_ci),
    .io_s(FullAdder_3233_io_s),
    .io_co(FullAdder_3233_io_co)
  );
  FullAdder FullAdder_3234 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3234_io_a),
    .io_b(FullAdder_3234_io_b),
    .io_ci(FullAdder_3234_io_ci),
    .io_s(FullAdder_3234_io_s),
    .io_co(FullAdder_3234_io_co)
  );
  FullAdder FullAdder_3235 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3235_io_a),
    .io_b(FullAdder_3235_io_b),
    .io_ci(FullAdder_3235_io_ci),
    .io_s(FullAdder_3235_io_s),
    .io_co(FullAdder_3235_io_co)
  );
  FullAdder FullAdder_3236 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3236_io_a),
    .io_b(FullAdder_3236_io_b),
    .io_ci(FullAdder_3236_io_ci),
    .io_s(FullAdder_3236_io_s),
    .io_co(FullAdder_3236_io_co)
  );
  FullAdder FullAdder_3237 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3237_io_a),
    .io_b(FullAdder_3237_io_b),
    .io_ci(FullAdder_3237_io_ci),
    .io_s(FullAdder_3237_io_s),
    .io_co(FullAdder_3237_io_co)
  );
  FullAdder FullAdder_3238 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3238_io_a),
    .io_b(FullAdder_3238_io_b),
    .io_ci(FullAdder_3238_io_ci),
    .io_s(FullAdder_3238_io_s),
    .io_co(FullAdder_3238_io_co)
  );
  FullAdder FullAdder_3239 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3239_io_a),
    .io_b(FullAdder_3239_io_b),
    .io_ci(FullAdder_3239_io_ci),
    .io_s(FullAdder_3239_io_s),
    .io_co(FullAdder_3239_io_co)
  );
  FullAdder FullAdder_3240 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3240_io_a),
    .io_b(FullAdder_3240_io_b),
    .io_ci(FullAdder_3240_io_ci),
    .io_s(FullAdder_3240_io_s),
    .io_co(FullAdder_3240_io_co)
  );
  FullAdder FullAdder_3241 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3241_io_a),
    .io_b(FullAdder_3241_io_b),
    .io_ci(FullAdder_3241_io_ci),
    .io_s(FullAdder_3241_io_s),
    .io_co(FullAdder_3241_io_co)
  );
  FullAdder FullAdder_3242 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3242_io_a),
    .io_b(FullAdder_3242_io_b),
    .io_ci(FullAdder_3242_io_ci),
    .io_s(FullAdder_3242_io_s),
    .io_co(FullAdder_3242_io_co)
  );
  FullAdder FullAdder_3243 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3243_io_a),
    .io_b(FullAdder_3243_io_b),
    .io_ci(FullAdder_3243_io_ci),
    .io_s(FullAdder_3243_io_s),
    .io_co(FullAdder_3243_io_co)
  );
  FullAdder FullAdder_3244 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3244_io_a),
    .io_b(FullAdder_3244_io_b),
    .io_ci(FullAdder_3244_io_ci),
    .io_s(FullAdder_3244_io_s),
    .io_co(FullAdder_3244_io_co)
  );
  FullAdder FullAdder_3245 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3245_io_a),
    .io_b(FullAdder_3245_io_b),
    .io_ci(FullAdder_3245_io_ci),
    .io_s(FullAdder_3245_io_s),
    .io_co(FullAdder_3245_io_co)
  );
  FullAdder FullAdder_3246 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3246_io_a),
    .io_b(FullAdder_3246_io_b),
    .io_ci(FullAdder_3246_io_ci),
    .io_s(FullAdder_3246_io_s),
    .io_co(FullAdder_3246_io_co)
  );
  FullAdder FullAdder_3247 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3247_io_a),
    .io_b(FullAdder_3247_io_b),
    .io_ci(FullAdder_3247_io_ci),
    .io_s(FullAdder_3247_io_s),
    .io_co(FullAdder_3247_io_co)
  );
  FullAdder FullAdder_3248 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3248_io_a),
    .io_b(FullAdder_3248_io_b),
    .io_ci(FullAdder_3248_io_ci),
    .io_s(FullAdder_3248_io_s),
    .io_co(FullAdder_3248_io_co)
  );
  FullAdder FullAdder_3249 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3249_io_a),
    .io_b(FullAdder_3249_io_b),
    .io_ci(FullAdder_3249_io_ci),
    .io_s(FullAdder_3249_io_s),
    .io_co(FullAdder_3249_io_co)
  );
  FullAdder FullAdder_3250 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3250_io_a),
    .io_b(FullAdder_3250_io_b),
    .io_ci(FullAdder_3250_io_ci),
    .io_s(FullAdder_3250_io_s),
    .io_co(FullAdder_3250_io_co)
  );
  FullAdder FullAdder_3251 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3251_io_a),
    .io_b(FullAdder_3251_io_b),
    .io_ci(FullAdder_3251_io_ci),
    .io_s(FullAdder_3251_io_s),
    .io_co(FullAdder_3251_io_co)
  );
  FullAdder FullAdder_3252 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3252_io_a),
    .io_b(FullAdder_3252_io_b),
    .io_ci(FullAdder_3252_io_ci),
    .io_s(FullAdder_3252_io_s),
    .io_co(FullAdder_3252_io_co)
  );
  FullAdder FullAdder_3253 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3253_io_a),
    .io_b(FullAdder_3253_io_b),
    .io_ci(FullAdder_3253_io_ci),
    .io_s(FullAdder_3253_io_s),
    .io_co(FullAdder_3253_io_co)
  );
  FullAdder FullAdder_3254 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3254_io_a),
    .io_b(FullAdder_3254_io_b),
    .io_ci(FullAdder_3254_io_ci),
    .io_s(FullAdder_3254_io_s),
    .io_co(FullAdder_3254_io_co)
  );
  FullAdder FullAdder_3255 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3255_io_a),
    .io_b(FullAdder_3255_io_b),
    .io_ci(FullAdder_3255_io_ci),
    .io_s(FullAdder_3255_io_s),
    .io_co(FullAdder_3255_io_co)
  );
  FullAdder FullAdder_3256 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3256_io_a),
    .io_b(FullAdder_3256_io_b),
    .io_ci(FullAdder_3256_io_ci),
    .io_s(FullAdder_3256_io_s),
    .io_co(FullAdder_3256_io_co)
  );
  FullAdder FullAdder_3257 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3257_io_a),
    .io_b(FullAdder_3257_io_b),
    .io_ci(FullAdder_3257_io_ci),
    .io_s(FullAdder_3257_io_s),
    .io_co(FullAdder_3257_io_co)
  );
  FullAdder FullAdder_3258 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3258_io_a),
    .io_b(FullAdder_3258_io_b),
    .io_ci(FullAdder_3258_io_ci),
    .io_s(FullAdder_3258_io_s),
    .io_co(FullAdder_3258_io_co)
  );
  FullAdder FullAdder_3259 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3259_io_a),
    .io_b(FullAdder_3259_io_b),
    .io_ci(FullAdder_3259_io_ci),
    .io_s(FullAdder_3259_io_s),
    .io_co(FullAdder_3259_io_co)
  );
  FullAdder FullAdder_3260 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3260_io_a),
    .io_b(FullAdder_3260_io_b),
    .io_ci(FullAdder_3260_io_ci),
    .io_s(FullAdder_3260_io_s),
    .io_co(FullAdder_3260_io_co)
  );
  FullAdder FullAdder_3261 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3261_io_a),
    .io_b(FullAdder_3261_io_b),
    .io_ci(FullAdder_3261_io_ci),
    .io_s(FullAdder_3261_io_s),
    .io_co(FullAdder_3261_io_co)
  );
  HalfAdder HalfAdder_127 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_127_io_a),
    .io_b(HalfAdder_127_io_b),
    .io_s(HalfAdder_127_io_s),
    .io_co(HalfAdder_127_io_co)
  );
  FullAdder FullAdder_3262 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3262_io_a),
    .io_b(FullAdder_3262_io_b),
    .io_ci(FullAdder_3262_io_ci),
    .io_s(FullAdder_3262_io_s),
    .io_co(FullAdder_3262_io_co)
  );
  FullAdder FullAdder_3263 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3263_io_a),
    .io_b(FullAdder_3263_io_b),
    .io_ci(FullAdder_3263_io_ci),
    .io_s(FullAdder_3263_io_s),
    .io_co(FullAdder_3263_io_co)
  );
  FullAdder FullAdder_3264 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3264_io_a),
    .io_b(FullAdder_3264_io_b),
    .io_ci(FullAdder_3264_io_ci),
    .io_s(FullAdder_3264_io_s),
    .io_co(FullAdder_3264_io_co)
  );
  HalfAdder HalfAdder_128 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_128_io_a),
    .io_b(HalfAdder_128_io_b),
    .io_s(HalfAdder_128_io_s),
    .io_co(HalfAdder_128_io_co)
  );
  FullAdder FullAdder_3265 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3265_io_a),
    .io_b(FullAdder_3265_io_b),
    .io_ci(FullAdder_3265_io_ci),
    .io_s(FullAdder_3265_io_s),
    .io_co(FullAdder_3265_io_co)
  );
  FullAdder FullAdder_3266 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3266_io_a),
    .io_b(FullAdder_3266_io_b),
    .io_ci(FullAdder_3266_io_ci),
    .io_s(FullAdder_3266_io_s),
    .io_co(FullAdder_3266_io_co)
  );
  FullAdder FullAdder_3267 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3267_io_a),
    .io_b(FullAdder_3267_io_b),
    .io_ci(FullAdder_3267_io_ci),
    .io_s(FullAdder_3267_io_s),
    .io_co(FullAdder_3267_io_co)
  );
  HalfAdder HalfAdder_129 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_129_io_a),
    .io_b(HalfAdder_129_io_b),
    .io_s(HalfAdder_129_io_s),
    .io_co(HalfAdder_129_io_co)
  );
  FullAdder FullAdder_3268 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3268_io_a),
    .io_b(FullAdder_3268_io_b),
    .io_ci(FullAdder_3268_io_ci),
    .io_s(FullAdder_3268_io_s),
    .io_co(FullAdder_3268_io_co)
  );
  FullAdder FullAdder_3269 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3269_io_a),
    .io_b(FullAdder_3269_io_b),
    .io_ci(FullAdder_3269_io_ci),
    .io_s(FullAdder_3269_io_s),
    .io_co(FullAdder_3269_io_co)
  );
  FullAdder FullAdder_3270 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3270_io_a),
    .io_b(FullAdder_3270_io_b),
    .io_ci(FullAdder_3270_io_ci),
    .io_s(FullAdder_3270_io_s),
    .io_co(FullAdder_3270_io_co)
  );
  FullAdder FullAdder_3271 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3271_io_a),
    .io_b(FullAdder_3271_io_b),
    .io_ci(FullAdder_3271_io_ci),
    .io_s(FullAdder_3271_io_s),
    .io_co(FullAdder_3271_io_co)
  );
  FullAdder FullAdder_3272 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3272_io_a),
    .io_b(FullAdder_3272_io_b),
    .io_ci(FullAdder_3272_io_ci),
    .io_s(FullAdder_3272_io_s),
    .io_co(FullAdder_3272_io_co)
  );
  FullAdder FullAdder_3273 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3273_io_a),
    .io_b(FullAdder_3273_io_b),
    .io_ci(FullAdder_3273_io_ci),
    .io_s(FullAdder_3273_io_s),
    .io_co(FullAdder_3273_io_co)
  );
  FullAdder FullAdder_3274 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3274_io_a),
    .io_b(FullAdder_3274_io_b),
    .io_ci(FullAdder_3274_io_ci),
    .io_s(FullAdder_3274_io_s),
    .io_co(FullAdder_3274_io_co)
  );
  FullAdder FullAdder_3275 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3275_io_a),
    .io_b(FullAdder_3275_io_b),
    .io_ci(FullAdder_3275_io_ci),
    .io_s(FullAdder_3275_io_s),
    .io_co(FullAdder_3275_io_co)
  );
  FullAdder FullAdder_3276 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3276_io_a),
    .io_b(FullAdder_3276_io_b),
    .io_ci(FullAdder_3276_io_ci),
    .io_s(FullAdder_3276_io_s),
    .io_co(FullAdder_3276_io_co)
  );
  FullAdder FullAdder_3277 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3277_io_a),
    .io_b(FullAdder_3277_io_b),
    .io_ci(FullAdder_3277_io_ci),
    .io_s(FullAdder_3277_io_s),
    .io_co(FullAdder_3277_io_co)
  );
  FullAdder FullAdder_3278 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3278_io_a),
    .io_b(FullAdder_3278_io_b),
    .io_ci(FullAdder_3278_io_ci),
    .io_s(FullAdder_3278_io_s),
    .io_co(FullAdder_3278_io_co)
  );
  FullAdder FullAdder_3279 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3279_io_a),
    .io_b(FullAdder_3279_io_b),
    .io_ci(FullAdder_3279_io_ci),
    .io_s(FullAdder_3279_io_s),
    .io_co(FullAdder_3279_io_co)
  );
  FullAdder FullAdder_3280 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3280_io_a),
    .io_b(FullAdder_3280_io_b),
    .io_ci(FullAdder_3280_io_ci),
    .io_s(FullAdder_3280_io_s),
    .io_co(FullAdder_3280_io_co)
  );
  FullAdder FullAdder_3281 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3281_io_a),
    .io_b(FullAdder_3281_io_b),
    .io_ci(FullAdder_3281_io_ci),
    .io_s(FullAdder_3281_io_s),
    .io_co(FullAdder_3281_io_co)
  );
  FullAdder FullAdder_3282 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3282_io_a),
    .io_b(FullAdder_3282_io_b),
    .io_ci(FullAdder_3282_io_ci),
    .io_s(FullAdder_3282_io_s),
    .io_co(FullAdder_3282_io_co)
  );
  FullAdder FullAdder_3283 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3283_io_a),
    .io_b(FullAdder_3283_io_b),
    .io_ci(FullAdder_3283_io_ci),
    .io_s(FullAdder_3283_io_s),
    .io_co(FullAdder_3283_io_co)
  );
  FullAdder FullAdder_3284 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3284_io_a),
    .io_b(FullAdder_3284_io_b),
    .io_ci(FullAdder_3284_io_ci),
    .io_s(FullAdder_3284_io_s),
    .io_co(FullAdder_3284_io_co)
  );
  FullAdder FullAdder_3285 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3285_io_a),
    .io_b(FullAdder_3285_io_b),
    .io_ci(FullAdder_3285_io_ci),
    .io_s(FullAdder_3285_io_s),
    .io_co(FullAdder_3285_io_co)
  );
  FullAdder FullAdder_3286 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3286_io_a),
    .io_b(FullAdder_3286_io_b),
    .io_ci(FullAdder_3286_io_ci),
    .io_s(FullAdder_3286_io_s),
    .io_co(FullAdder_3286_io_co)
  );
  FullAdder FullAdder_3287 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3287_io_a),
    .io_b(FullAdder_3287_io_b),
    .io_ci(FullAdder_3287_io_ci),
    .io_s(FullAdder_3287_io_s),
    .io_co(FullAdder_3287_io_co)
  );
  FullAdder FullAdder_3288 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3288_io_a),
    .io_b(FullAdder_3288_io_b),
    .io_ci(FullAdder_3288_io_ci),
    .io_s(FullAdder_3288_io_s),
    .io_co(FullAdder_3288_io_co)
  );
  FullAdder FullAdder_3289 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3289_io_a),
    .io_b(FullAdder_3289_io_b),
    .io_ci(FullAdder_3289_io_ci),
    .io_s(FullAdder_3289_io_s),
    .io_co(FullAdder_3289_io_co)
  );
  FullAdder FullAdder_3290 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3290_io_a),
    .io_b(FullAdder_3290_io_b),
    .io_ci(FullAdder_3290_io_ci),
    .io_s(FullAdder_3290_io_s),
    .io_co(FullAdder_3290_io_co)
  );
  FullAdder FullAdder_3291 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3291_io_a),
    .io_b(FullAdder_3291_io_b),
    .io_ci(FullAdder_3291_io_ci),
    .io_s(FullAdder_3291_io_s),
    .io_co(FullAdder_3291_io_co)
  );
  FullAdder FullAdder_3292 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3292_io_a),
    .io_b(FullAdder_3292_io_b),
    .io_ci(FullAdder_3292_io_ci),
    .io_s(FullAdder_3292_io_s),
    .io_co(FullAdder_3292_io_co)
  );
  FullAdder FullAdder_3293 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3293_io_a),
    .io_b(FullAdder_3293_io_b),
    .io_ci(FullAdder_3293_io_ci),
    .io_s(FullAdder_3293_io_s),
    .io_co(FullAdder_3293_io_co)
  );
  FullAdder FullAdder_3294 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3294_io_a),
    .io_b(FullAdder_3294_io_b),
    .io_ci(FullAdder_3294_io_ci),
    .io_s(FullAdder_3294_io_s),
    .io_co(FullAdder_3294_io_co)
  );
  FullAdder FullAdder_3295 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3295_io_a),
    .io_b(FullAdder_3295_io_b),
    .io_ci(FullAdder_3295_io_ci),
    .io_s(FullAdder_3295_io_s),
    .io_co(FullAdder_3295_io_co)
  );
  FullAdder FullAdder_3296 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3296_io_a),
    .io_b(FullAdder_3296_io_b),
    .io_ci(FullAdder_3296_io_ci),
    .io_s(FullAdder_3296_io_s),
    .io_co(FullAdder_3296_io_co)
  );
  FullAdder FullAdder_3297 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3297_io_a),
    .io_b(FullAdder_3297_io_b),
    .io_ci(FullAdder_3297_io_ci),
    .io_s(FullAdder_3297_io_s),
    .io_co(FullAdder_3297_io_co)
  );
  FullAdder FullAdder_3298 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3298_io_a),
    .io_b(FullAdder_3298_io_b),
    .io_ci(FullAdder_3298_io_ci),
    .io_s(FullAdder_3298_io_s),
    .io_co(FullAdder_3298_io_co)
  );
  FullAdder FullAdder_3299 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3299_io_a),
    .io_b(FullAdder_3299_io_b),
    .io_ci(FullAdder_3299_io_ci),
    .io_s(FullAdder_3299_io_s),
    .io_co(FullAdder_3299_io_co)
  );
  FullAdder FullAdder_3300 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3300_io_a),
    .io_b(FullAdder_3300_io_b),
    .io_ci(FullAdder_3300_io_ci),
    .io_s(FullAdder_3300_io_s),
    .io_co(FullAdder_3300_io_co)
  );
  FullAdder FullAdder_3301 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3301_io_a),
    .io_b(FullAdder_3301_io_b),
    .io_ci(FullAdder_3301_io_ci),
    .io_s(FullAdder_3301_io_s),
    .io_co(FullAdder_3301_io_co)
  );
  FullAdder FullAdder_3302 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3302_io_a),
    .io_b(FullAdder_3302_io_b),
    .io_ci(FullAdder_3302_io_ci),
    .io_s(FullAdder_3302_io_s),
    .io_co(FullAdder_3302_io_co)
  );
  FullAdder FullAdder_3303 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3303_io_a),
    .io_b(FullAdder_3303_io_b),
    .io_ci(FullAdder_3303_io_ci),
    .io_s(FullAdder_3303_io_s),
    .io_co(FullAdder_3303_io_co)
  );
  FullAdder FullAdder_3304 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3304_io_a),
    .io_b(FullAdder_3304_io_b),
    .io_ci(FullAdder_3304_io_ci),
    .io_s(FullAdder_3304_io_s),
    .io_co(FullAdder_3304_io_co)
  );
  FullAdder FullAdder_3305 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3305_io_a),
    .io_b(FullAdder_3305_io_b),
    .io_ci(FullAdder_3305_io_ci),
    .io_s(FullAdder_3305_io_s),
    .io_co(FullAdder_3305_io_co)
  );
  FullAdder FullAdder_3306 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3306_io_a),
    .io_b(FullAdder_3306_io_b),
    .io_ci(FullAdder_3306_io_ci),
    .io_s(FullAdder_3306_io_s),
    .io_co(FullAdder_3306_io_co)
  );
  FullAdder FullAdder_3307 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3307_io_a),
    .io_b(FullAdder_3307_io_b),
    .io_ci(FullAdder_3307_io_ci),
    .io_s(FullAdder_3307_io_s),
    .io_co(FullAdder_3307_io_co)
  );
  HalfAdder HalfAdder_130 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_130_io_a),
    .io_b(HalfAdder_130_io_b),
    .io_s(HalfAdder_130_io_s),
    .io_co(HalfAdder_130_io_co)
  );
  FullAdder FullAdder_3308 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3308_io_a),
    .io_b(FullAdder_3308_io_b),
    .io_ci(FullAdder_3308_io_ci),
    .io_s(FullAdder_3308_io_s),
    .io_co(FullAdder_3308_io_co)
  );
  FullAdder FullAdder_3309 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3309_io_a),
    .io_b(FullAdder_3309_io_b),
    .io_ci(FullAdder_3309_io_ci),
    .io_s(FullAdder_3309_io_s),
    .io_co(FullAdder_3309_io_co)
  );
  FullAdder FullAdder_3310 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3310_io_a),
    .io_b(FullAdder_3310_io_b),
    .io_ci(FullAdder_3310_io_ci),
    .io_s(FullAdder_3310_io_s),
    .io_co(FullAdder_3310_io_co)
  );
  FullAdder FullAdder_3311 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3311_io_a),
    .io_b(FullAdder_3311_io_b),
    .io_ci(FullAdder_3311_io_ci),
    .io_s(FullAdder_3311_io_s),
    .io_co(FullAdder_3311_io_co)
  );
  FullAdder FullAdder_3312 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3312_io_a),
    .io_b(FullAdder_3312_io_b),
    .io_ci(FullAdder_3312_io_ci),
    .io_s(FullAdder_3312_io_s),
    .io_co(FullAdder_3312_io_co)
  );
  FullAdder FullAdder_3313 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3313_io_a),
    .io_b(FullAdder_3313_io_b),
    .io_ci(FullAdder_3313_io_ci),
    .io_s(FullAdder_3313_io_s),
    .io_co(FullAdder_3313_io_co)
  );
  FullAdder FullAdder_3314 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3314_io_a),
    .io_b(FullAdder_3314_io_b),
    .io_ci(FullAdder_3314_io_ci),
    .io_s(FullAdder_3314_io_s),
    .io_co(FullAdder_3314_io_co)
  );
  FullAdder FullAdder_3315 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3315_io_a),
    .io_b(FullAdder_3315_io_b),
    .io_ci(FullAdder_3315_io_ci),
    .io_s(FullAdder_3315_io_s),
    .io_co(FullAdder_3315_io_co)
  );
  FullAdder FullAdder_3316 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3316_io_a),
    .io_b(FullAdder_3316_io_b),
    .io_ci(FullAdder_3316_io_ci),
    .io_s(FullAdder_3316_io_s),
    .io_co(FullAdder_3316_io_co)
  );
  FullAdder FullAdder_3317 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3317_io_a),
    .io_b(FullAdder_3317_io_b),
    .io_ci(FullAdder_3317_io_ci),
    .io_s(FullAdder_3317_io_s),
    .io_co(FullAdder_3317_io_co)
  );
  FullAdder FullAdder_3318 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3318_io_a),
    .io_b(FullAdder_3318_io_b),
    .io_ci(FullAdder_3318_io_ci),
    .io_s(FullAdder_3318_io_s),
    .io_co(FullAdder_3318_io_co)
  );
  FullAdder FullAdder_3319 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3319_io_a),
    .io_b(FullAdder_3319_io_b),
    .io_ci(FullAdder_3319_io_ci),
    .io_s(FullAdder_3319_io_s),
    .io_co(FullAdder_3319_io_co)
  );
  FullAdder FullAdder_3320 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3320_io_a),
    .io_b(FullAdder_3320_io_b),
    .io_ci(FullAdder_3320_io_ci),
    .io_s(FullAdder_3320_io_s),
    .io_co(FullAdder_3320_io_co)
  );
  FullAdder FullAdder_3321 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3321_io_a),
    .io_b(FullAdder_3321_io_b),
    .io_ci(FullAdder_3321_io_ci),
    .io_s(FullAdder_3321_io_s),
    .io_co(FullAdder_3321_io_co)
  );
  FullAdder FullAdder_3322 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3322_io_a),
    .io_b(FullAdder_3322_io_b),
    .io_ci(FullAdder_3322_io_ci),
    .io_s(FullAdder_3322_io_s),
    .io_co(FullAdder_3322_io_co)
  );
  FullAdder FullAdder_3323 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3323_io_a),
    .io_b(FullAdder_3323_io_b),
    .io_ci(FullAdder_3323_io_ci),
    .io_s(FullAdder_3323_io_s),
    .io_co(FullAdder_3323_io_co)
  );
  FullAdder FullAdder_3324 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3324_io_a),
    .io_b(FullAdder_3324_io_b),
    .io_ci(FullAdder_3324_io_ci),
    .io_s(FullAdder_3324_io_s),
    .io_co(FullAdder_3324_io_co)
  );
  FullAdder FullAdder_3325 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3325_io_a),
    .io_b(FullAdder_3325_io_b),
    .io_ci(FullAdder_3325_io_ci),
    .io_s(FullAdder_3325_io_s),
    .io_co(FullAdder_3325_io_co)
  );
  FullAdder FullAdder_3326 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3326_io_a),
    .io_b(FullAdder_3326_io_b),
    .io_ci(FullAdder_3326_io_ci),
    .io_s(FullAdder_3326_io_s),
    .io_co(FullAdder_3326_io_co)
  );
  FullAdder FullAdder_3327 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3327_io_a),
    .io_b(FullAdder_3327_io_b),
    .io_ci(FullAdder_3327_io_ci),
    .io_s(FullAdder_3327_io_s),
    .io_co(FullAdder_3327_io_co)
  );
  FullAdder FullAdder_3328 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3328_io_a),
    .io_b(FullAdder_3328_io_b),
    .io_ci(FullAdder_3328_io_ci),
    .io_s(FullAdder_3328_io_s),
    .io_co(FullAdder_3328_io_co)
  );
  FullAdder FullAdder_3329 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3329_io_a),
    .io_b(FullAdder_3329_io_b),
    .io_ci(FullAdder_3329_io_ci),
    .io_s(FullAdder_3329_io_s),
    .io_co(FullAdder_3329_io_co)
  );
  FullAdder FullAdder_3330 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3330_io_a),
    .io_b(FullAdder_3330_io_b),
    .io_ci(FullAdder_3330_io_ci),
    .io_s(FullAdder_3330_io_s),
    .io_co(FullAdder_3330_io_co)
  );
  FullAdder FullAdder_3331 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3331_io_a),
    .io_b(FullAdder_3331_io_b),
    .io_ci(FullAdder_3331_io_ci),
    .io_s(FullAdder_3331_io_s),
    .io_co(FullAdder_3331_io_co)
  );
  FullAdder FullAdder_3332 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3332_io_a),
    .io_b(FullAdder_3332_io_b),
    .io_ci(FullAdder_3332_io_ci),
    .io_s(FullAdder_3332_io_s),
    .io_co(FullAdder_3332_io_co)
  );
  FullAdder FullAdder_3333 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3333_io_a),
    .io_b(FullAdder_3333_io_b),
    .io_ci(FullAdder_3333_io_ci),
    .io_s(FullAdder_3333_io_s),
    .io_co(FullAdder_3333_io_co)
  );
  FullAdder FullAdder_3334 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3334_io_a),
    .io_b(FullAdder_3334_io_b),
    .io_ci(FullAdder_3334_io_ci),
    .io_s(FullAdder_3334_io_s),
    .io_co(FullAdder_3334_io_co)
  );
  FullAdder FullAdder_3335 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3335_io_a),
    .io_b(FullAdder_3335_io_b),
    .io_ci(FullAdder_3335_io_ci),
    .io_s(FullAdder_3335_io_s),
    .io_co(FullAdder_3335_io_co)
  );
  FullAdder FullAdder_3336 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3336_io_a),
    .io_b(FullAdder_3336_io_b),
    .io_ci(FullAdder_3336_io_ci),
    .io_s(FullAdder_3336_io_s),
    .io_co(FullAdder_3336_io_co)
  );
  FullAdder FullAdder_3337 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3337_io_a),
    .io_b(FullAdder_3337_io_b),
    .io_ci(FullAdder_3337_io_ci),
    .io_s(FullAdder_3337_io_s),
    .io_co(FullAdder_3337_io_co)
  );
  FullAdder FullAdder_3338 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3338_io_a),
    .io_b(FullAdder_3338_io_b),
    .io_ci(FullAdder_3338_io_ci),
    .io_s(FullAdder_3338_io_s),
    .io_co(FullAdder_3338_io_co)
  );
  FullAdder FullAdder_3339 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3339_io_a),
    .io_b(FullAdder_3339_io_b),
    .io_ci(FullAdder_3339_io_ci),
    .io_s(FullAdder_3339_io_s),
    .io_co(FullAdder_3339_io_co)
  );
  FullAdder FullAdder_3340 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3340_io_a),
    .io_b(FullAdder_3340_io_b),
    .io_ci(FullAdder_3340_io_ci),
    .io_s(FullAdder_3340_io_s),
    .io_co(FullAdder_3340_io_co)
  );
  FullAdder FullAdder_3341 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3341_io_a),
    .io_b(FullAdder_3341_io_b),
    .io_ci(FullAdder_3341_io_ci),
    .io_s(FullAdder_3341_io_s),
    .io_co(FullAdder_3341_io_co)
  );
  FullAdder FullAdder_3342 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3342_io_a),
    .io_b(FullAdder_3342_io_b),
    .io_ci(FullAdder_3342_io_ci),
    .io_s(FullAdder_3342_io_s),
    .io_co(FullAdder_3342_io_co)
  );
  FullAdder FullAdder_3343 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3343_io_a),
    .io_b(FullAdder_3343_io_b),
    .io_ci(FullAdder_3343_io_ci),
    .io_s(FullAdder_3343_io_s),
    .io_co(FullAdder_3343_io_co)
  );
  FullAdder FullAdder_3344 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3344_io_a),
    .io_b(FullAdder_3344_io_b),
    .io_ci(FullAdder_3344_io_ci),
    .io_s(FullAdder_3344_io_s),
    .io_co(FullAdder_3344_io_co)
  );
  FullAdder FullAdder_3345 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3345_io_a),
    .io_b(FullAdder_3345_io_b),
    .io_ci(FullAdder_3345_io_ci),
    .io_s(FullAdder_3345_io_s),
    .io_co(FullAdder_3345_io_co)
  );
  FullAdder FullAdder_3346 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3346_io_a),
    .io_b(FullAdder_3346_io_b),
    .io_ci(FullAdder_3346_io_ci),
    .io_s(FullAdder_3346_io_s),
    .io_co(FullAdder_3346_io_co)
  );
  FullAdder FullAdder_3347 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3347_io_a),
    .io_b(FullAdder_3347_io_b),
    .io_ci(FullAdder_3347_io_ci),
    .io_s(FullAdder_3347_io_s),
    .io_co(FullAdder_3347_io_co)
  );
  FullAdder FullAdder_3348 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3348_io_a),
    .io_b(FullAdder_3348_io_b),
    .io_ci(FullAdder_3348_io_ci),
    .io_s(FullAdder_3348_io_s),
    .io_co(FullAdder_3348_io_co)
  );
  HalfAdder HalfAdder_131 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_131_io_a),
    .io_b(HalfAdder_131_io_b),
    .io_s(HalfAdder_131_io_s),
    .io_co(HalfAdder_131_io_co)
  );
  FullAdder FullAdder_3349 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3349_io_a),
    .io_b(FullAdder_3349_io_b),
    .io_ci(FullAdder_3349_io_ci),
    .io_s(FullAdder_3349_io_s),
    .io_co(FullAdder_3349_io_co)
  );
  FullAdder FullAdder_3350 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3350_io_a),
    .io_b(FullAdder_3350_io_b),
    .io_ci(FullAdder_3350_io_ci),
    .io_s(FullAdder_3350_io_s),
    .io_co(FullAdder_3350_io_co)
  );
  FullAdder FullAdder_3351 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3351_io_a),
    .io_b(FullAdder_3351_io_b),
    .io_ci(FullAdder_3351_io_ci),
    .io_s(FullAdder_3351_io_s),
    .io_co(FullAdder_3351_io_co)
  );
  FullAdder FullAdder_3352 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3352_io_a),
    .io_b(FullAdder_3352_io_b),
    .io_ci(FullAdder_3352_io_ci),
    .io_s(FullAdder_3352_io_s),
    .io_co(FullAdder_3352_io_co)
  );
  FullAdder FullAdder_3353 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3353_io_a),
    .io_b(FullAdder_3353_io_b),
    .io_ci(FullAdder_3353_io_ci),
    .io_s(FullAdder_3353_io_s),
    .io_co(FullAdder_3353_io_co)
  );
  FullAdder FullAdder_3354 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3354_io_a),
    .io_b(FullAdder_3354_io_b),
    .io_ci(FullAdder_3354_io_ci),
    .io_s(FullAdder_3354_io_s),
    .io_co(FullAdder_3354_io_co)
  );
  FullAdder FullAdder_3355 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3355_io_a),
    .io_b(FullAdder_3355_io_b),
    .io_ci(FullAdder_3355_io_ci),
    .io_s(FullAdder_3355_io_s),
    .io_co(FullAdder_3355_io_co)
  );
  FullAdder FullAdder_3356 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3356_io_a),
    .io_b(FullAdder_3356_io_b),
    .io_ci(FullAdder_3356_io_ci),
    .io_s(FullAdder_3356_io_s),
    .io_co(FullAdder_3356_io_co)
  );
  FullAdder FullAdder_3357 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3357_io_a),
    .io_b(FullAdder_3357_io_b),
    .io_ci(FullAdder_3357_io_ci),
    .io_s(FullAdder_3357_io_s),
    .io_co(FullAdder_3357_io_co)
  );
  FullAdder FullAdder_3358 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3358_io_a),
    .io_b(FullAdder_3358_io_b),
    .io_ci(FullAdder_3358_io_ci),
    .io_s(FullAdder_3358_io_s),
    .io_co(FullAdder_3358_io_co)
  );
  FullAdder FullAdder_3359 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3359_io_a),
    .io_b(FullAdder_3359_io_b),
    .io_ci(FullAdder_3359_io_ci),
    .io_s(FullAdder_3359_io_s),
    .io_co(FullAdder_3359_io_co)
  );
  FullAdder FullAdder_3360 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3360_io_a),
    .io_b(FullAdder_3360_io_b),
    .io_ci(FullAdder_3360_io_ci),
    .io_s(FullAdder_3360_io_s),
    .io_co(FullAdder_3360_io_co)
  );
  FullAdder FullAdder_3361 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3361_io_a),
    .io_b(FullAdder_3361_io_b),
    .io_ci(FullAdder_3361_io_ci),
    .io_s(FullAdder_3361_io_s),
    .io_co(FullAdder_3361_io_co)
  );
  FullAdder FullAdder_3362 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3362_io_a),
    .io_b(FullAdder_3362_io_b),
    .io_ci(FullAdder_3362_io_ci),
    .io_s(FullAdder_3362_io_s),
    .io_co(FullAdder_3362_io_co)
  );
  FullAdder FullAdder_3363 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3363_io_a),
    .io_b(FullAdder_3363_io_b),
    .io_ci(FullAdder_3363_io_ci),
    .io_s(FullAdder_3363_io_s),
    .io_co(FullAdder_3363_io_co)
  );
  FullAdder FullAdder_3364 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3364_io_a),
    .io_b(FullAdder_3364_io_b),
    .io_ci(FullAdder_3364_io_ci),
    .io_s(FullAdder_3364_io_s),
    .io_co(FullAdder_3364_io_co)
  );
  FullAdder FullAdder_3365 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3365_io_a),
    .io_b(FullAdder_3365_io_b),
    .io_ci(FullAdder_3365_io_ci),
    .io_s(FullAdder_3365_io_s),
    .io_co(FullAdder_3365_io_co)
  );
  FullAdder FullAdder_3366 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3366_io_a),
    .io_b(FullAdder_3366_io_b),
    .io_ci(FullAdder_3366_io_ci),
    .io_s(FullAdder_3366_io_s),
    .io_co(FullAdder_3366_io_co)
  );
  FullAdder FullAdder_3367 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3367_io_a),
    .io_b(FullAdder_3367_io_b),
    .io_ci(FullAdder_3367_io_ci),
    .io_s(FullAdder_3367_io_s),
    .io_co(FullAdder_3367_io_co)
  );
  FullAdder FullAdder_3368 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3368_io_a),
    .io_b(FullAdder_3368_io_b),
    .io_ci(FullAdder_3368_io_ci),
    .io_s(FullAdder_3368_io_s),
    .io_co(FullAdder_3368_io_co)
  );
  FullAdder FullAdder_3369 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3369_io_a),
    .io_b(FullAdder_3369_io_b),
    .io_ci(FullAdder_3369_io_ci),
    .io_s(FullAdder_3369_io_s),
    .io_co(FullAdder_3369_io_co)
  );
  FullAdder FullAdder_3370 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3370_io_a),
    .io_b(FullAdder_3370_io_b),
    .io_ci(FullAdder_3370_io_ci),
    .io_s(FullAdder_3370_io_s),
    .io_co(FullAdder_3370_io_co)
  );
  FullAdder FullAdder_3371 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3371_io_a),
    .io_b(FullAdder_3371_io_b),
    .io_ci(FullAdder_3371_io_ci),
    .io_s(FullAdder_3371_io_s),
    .io_co(FullAdder_3371_io_co)
  );
  FullAdder FullAdder_3372 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3372_io_a),
    .io_b(FullAdder_3372_io_b),
    .io_ci(FullAdder_3372_io_ci),
    .io_s(FullAdder_3372_io_s),
    .io_co(FullAdder_3372_io_co)
  );
  FullAdder FullAdder_3373 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3373_io_a),
    .io_b(FullAdder_3373_io_b),
    .io_ci(FullAdder_3373_io_ci),
    .io_s(FullAdder_3373_io_s),
    .io_co(FullAdder_3373_io_co)
  );
  FullAdder FullAdder_3374 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3374_io_a),
    .io_b(FullAdder_3374_io_b),
    .io_ci(FullAdder_3374_io_ci),
    .io_s(FullAdder_3374_io_s),
    .io_co(FullAdder_3374_io_co)
  );
  FullAdder FullAdder_3375 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3375_io_a),
    .io_b(FullAdder_3375_io_b),
    .io_ci(FullAdder_3375_io_ci),
    .io_s(FullAdder_3375_io_s),
    .io_co(FullAdder_3375_io_co)
  );
  FullAdder FullAdder_3376 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3376_io_a),
    .io_b(FullAdder_3376_io_b),
    .io_ci(FullAdder_3376_io_ci),
    .io_s(FullAdder_3376_io_s),
    .io_co(FullAdder_3376_io_co)
  );
  FullAdder FullAdder_3377 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3377_io_a),
    .io_b(FullAdder_3377_io_b),
    .io_ci(FullAdder_3377_io_ci),
    .io_s(FullAdder_3377_io_s),
    .io_co(FullAdder_3377_io_co)
  );
  FullAdder FullAdder_3378 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3378_io_a),
    .io_b(FullAdder_3378_io_b),
    .io_ci(FullAdder_3378_io_ci),
    .io_s(FullAdder_3378_io_s),
    .io_co(FullAdder_3378_io_co)
  );
  FullAdder FullAdder_3379 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3379_io_a),
    .io_b(FullAdder_3379_io_b),
    .io_ci(FullAdder_3379_io_ci),
    .io_s(FullAdder_3379_io_s),
    .io_co(FullAdder_3379_io_co)
  );
  FullAdder FullAdder_3380 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3380_io_a),
    .io_b(FullAdder_3380_io_b),
    .io_ci(FullAdder_3380_io_ci),
    .io_s(FullAdder_3380_io_s),
    .io_co(FullAdder_3380_io_co)
  );
  FullAdder FullAdder_3381 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3381_io_a),
    .io_b(FullAdder_3381_io_b),
    .io_ci(FullAdder_3381_io_ci),
    .io_s(FullAdder_3381_io_s),
    .io_co(FullAdder_3381_io_co)
  );
  FullAdder FullAdder_3382 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3382_io_a),
    .io_b(FullAdder_3382_io_b),
    .io_ci(FullAdder_3382_io_ci),
    .io_s(FullAdder_3382_io_s),
    .io_co(FullAdder_3382_io_co)
  );
  FullAdder FullAdder_3383 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3383_io_a),
    .io_b(FullAdder_3383_io_b),
    .io_ci(FullAdder_3383_io_ci),
    .io_s(FullAdder_3383_io_s),
    .io_co(FullAdder_3383_io_co)
  );
  FullAdder FullAdder_3384 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3384_io_a),
    .io_b(FullAdder_3384_io_b),
    .io_ci(FullAdder_3384_io_ci),
    .io_s(FullAdder_3384_io_s),
    .io_co(FullAdder_3384_io_co)
  );
  FullAdder FullAdder_3385 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3385_io_a),
    .io_b(FullAdder_3385_io_b),
    .io_ci(FullAdder_3385_io_ci),
    .io_s(FullAdder_3385_io_s),
    .io_co(FullAdder_3385_io_co)
  );
  FullAdder FullAdder_3386 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3386_io_a),
    .io_b(FullAdder_3386_io_b),
    .io_ci(FullAdder_3386_io_ci),
    .io_s(FullAdder_3386_io_s),
    .io_co(FullAdder_3386_io_co)
  );
  FullAdder FullAdder_3387 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3387_io_a),
    .io_b(FullAdder_3387_io_b),
    .io_ci(FullAdder_3387_io_ci),
    .io_s(FullAdder_3387_io_s),
    .io_co(FullAdder_3387_io_co)
  );
  FullAdder FullAdder_3388 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3388_io_a),
    .io_b(FullAdder_3388_io_b),
    .io_ci(FullAdder_3388_io_ci),
    .io_s(FullAdder_3388_io_s),
    .io_co(FullAdder_3388_io_co)
  );
  HalfAdder HalfAdder_132 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_132_io_a),
    .io_b(HalfAdder_132_io_b),
    .io_s(HalfAdder_132_io_s),
    .io_co(HalfAdder_132_io_co)
  );
  FullAdder FullAdder_3389 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3389_io_a),
    .io_b(FullAdder_3389_io_b),
    .io_ci(FullAdder_3389_io_ci),
    .io_s(FullAdder_3389_io_s),
    .io_co(FullAdder_3389_io_co)
  );
  FullAdder FullAdder_3390 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3390_io_a),
    .io_b(FullAdder_3390_io_b),
    .io_ci(FullAdder_3390_io_ci),
    .io_s(FullAdder_3390_io_s),
    .io_co(FullAdder_3390_io_co)
  );
  FullAdder FullAdder_3391 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3391_io_a),
    .io_b(FullAdder_3391_io_b),
    .io_ci(FullAdder_3391_io_ci),
    .io_s(FullAdder_3391_io_s),
    .io_co(FullAdder_3391_io_co)
  );
  FullAdder FullAdder_3392 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3392_io_a),
    .io_b(FullAdder_3392_io_b),
    .io_ci(FullAdder_3392_io_ci),
    .io_s(FullAdder_3392_io_s),
    .io_co(FullAdder_3392_io_co)
  );
  FullAdder FullAdder_3393 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3393_io_a),
    .io_b(FullAdder_3393_io_b),
    .io_ci(FullAdder_3393_io_ci),
    .io_s(FullAdder_3393_io_s),
    .io_co(FullAdder_3393_io_co)
  );
  FullAdder FullAdder_3394 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3394_io_a),
    .io_b(FullAdder_3394_io_b),
    .io_ci(FullAdder_3394_io_ci),
    .io_s(FullAdder_3394_io_s),
    .io_co(FullAdder_3394_io_co)
  );
  FullAdder FullAdder_3395 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3395_io_a),
    .io_b(FullAdder_3395_io_b),
    .io_ci(FullAdder_3395_io_ci),
    .io_s(FullAdder_3395_io_s),
    .io_co(FullAdder_3395_io_co)
  );
  FullAdder FullAdder_3396 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3396_io_a),
    .io_b(FullAdder_3396_io_b),
    .io_ci(FullAdder_3396_io_ci),
    .io_s(FullAdder_3396_io_s),
    .io_co(FullAdder_3396_io_co)
  );
  FullAdder FullAdder_3397 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3397_io_a),
    .io_b(FullAdder_3397_io_b),
    .io_ci(FullAdder_3397_io_ci),
    .io_s(FullAdder_3397_io_s),
    .io_co(FullAdder_3397_io_co)
  );
  FullAdder FullAdder_3398 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3398_io_a),
    .io_b(FullAdder_3398_io_b),
    .io_ci(FullAdder_3398_io_ci),
    .io_s(FullAdder_3398_io_s),
    .io_co(FullAdder_3398_io_co)
  );
  FullAdder FullAdder_3399 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3399_io_a),
    .io_b(FullAdder_3399_io_b),
    .io_ci(FullAdder_3399_io_ci),
    .io_s(FullAdder_3399_io_s),
    .io_co(FullAdder_3399_io_co)
  );
  FullAdder FullAdder_3400 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3400_io_a),
    .io_b(FullAdder_3400_io_b),
    .io_ci(FullAdder_3400_io_ci),
    .io_s(FullAdder_3400_io_s),
    .io_co(FullAdder_3400_io_co)
  );
  FullAdder FullAdder_3401 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3401_io_a),
    .io_b(FullAdder_3401_io_b),
    .io_ci(FullAdder_3401_io_ci),
    .io_s(FullAdder_3401_io_s),
    .io_co(FullAdder_3401_io_co)
  );
  FullAdder FullAdder_3402 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3402_io_a),
    .io_b(FullAdder_3402_io_b),
    .io_ci(FullAdder_3402_io_ci),
    .io_s(FullAdder_3402_io_s),
    .io_co(FullAdder_3402_io_co)
  );
  HalfAdder HalfAdder_133 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_133_io_a),
    .io_b(HalfAdder_133_io_b),
    .io_s(HalfAdder_133_io_s),
    .io_co(HalfAdder_133_io_co)
  );
  FullAdder FullAdder_3403 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3403_io_a),
    .io_b(FullAdder_3403_io_b),
    .io_ci(FullAdder_3403_io_ci),
    .io_s(FullAdder_3403_io_s),
    .io_co(FullAdder_3403_io_co)
  );
  FullAdder FullAdder_3404 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3404_io_a),
    .io_b(FullAdder_3404_io_b),
    .io_ci(FullAdder_3404_io_ci),
    .io_s(FullAdder_3404_io_s),
    .io_co(FullAdder_3404_io_co)
  );
  FullAdder FullAdder_3405 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3405_io_a),
    .io_b(FullAdder_3405_io_b),
    .io_ci(FullAdder_3405_io_ci),
    .io_s(FullAdder_3405_io_s),
    .io_co(FullAdder_3405_io_co)
  );
  FullAdder FullAdder_3406 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3406_io_a),
    .io_b(FullAdder_3406_io_b),
    .io_ci(FullAdder_3406_io_ci),
    .io_s(FullAdder_3406_io_s),
    .io_co(FullAdder_3406_io_co)
  );
  FullAdder FullAdder_3407 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3407_io_a),
    .io_b(FullAdder_3407_io_b),
    .io_ci(FullAdder_3407_io_ci),
    .io_s(FullAdder_3407_io_s),
    .io_co(FullAdder_3407_io_co)
  );
  FullAdder FullAdder_3408 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3408_io_a),
    .io_b(FullAdder_3408_io_b),
    .io_ci(FullAdder_3408_io_ci),
    .io_s(FullAdder_3408_io_s),
    .io_co(FullAdder_3408_io_co)
  );
  FullAdder FullAdder_3409 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3409_io_a),
    .io_b(FullAdder_3409_io_b),
    .io_ci(FullAdder_3409_io_ci),
    .io_s(FullAdder_3409_io_s),
    .io_co(FullAdder_3409_io_co)
  );
  FullAdder FullAdder_3410 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3410_io_a),
    .io_b(FullAdder_3410_io_b),
    .io_ci(FullAdder_3410_io_ci),
    .io_s(FullAdder_3410_io_s),
    .io_co(FullAdder_3410_io_co)
  );
  FullAdder FullAdder_3411 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3411_io_a),
    .io_b(FullAdder_3411_io_b),
    .io_ci(FullAdder_3411_io_ci),
    .io_s(FullAdder_3411_io_s),
    .io_co(FullAdder_3411_io_co)
  );
  FullAdder FullAdder_3412 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3412_io_a),
    .io_b(FullAdder_3412_io_b),
    .io_ci(FullAdder_3412_io_ci),
    .io_s(FullAdder_3412_io_s),
    .io_co(FullAdder_3412_io_co)
  );
  FullAdder FullAdder_3413 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3413_io_a),
    .io_b(FullAdder_3413_io_b),
    .io_ci(FullAdder_3413_io_ci),
    .io_s(FullAdder_3413_io_s),
    .io_co(FullAdder_3413_io_co)
  );
  FullAdder FullAdder_3414 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3414_io_a),
    .io_b(FullAdder_3414_io_b),
    .io_ci(FullAdder_3414_io_ci),
    .io_s(FullAdder_3414_io_s),
    .io_co(FullAdder_3414_io_co)
  );
  FullAdder FullAdder_3415 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3415_io_a),
    .io_b(FullAdder_3415_io_b),
    .io_ci(FullAdder_3415_io_ci),
    .io_s(FullAdder_3415_io_s),
    .io_co(FullAdder_3415_io_co)
  );
  FullAdder FullAdder_3416 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3416_io_a),
    .io_b(FullAdder_3416_io_b),
    .io_ci(FullAdder_3416_io_ci),
    .io_s(FullAdder_3416_io_s),
    .io_co(FullAdder_3416_io_co)
  );
  FullAdder FullAdder_3417 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3417_io_a),
    .io_b(FullAdder_3417_io_b),
    .io_ci(FullAdder_3417_io_ci),
    .io_s(FullAdder_3417_io_s),
    .io_co(FullAdder_3417_io_co)
  );
  FullAdder FullAdder_3418 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3418_io_a),
    .io_b(FullAdder_3418_io_b),
    .io_ci(FullAdder_3418_io_ci),
    .io_s(FullAdder_3418_io_s),
    .io_co(FullAdder_3418_io_co)
  );
  FullAdder FullAdder_3419 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3419_io_a),
    .io_b(FullAdder_3419_io_b),
    .io_ci(FullAdder_3419_io_ci),
    .io_s(FullAdder_3419_io_s),
    .io_co(FullAdder_3419_io_co)
  );
  FullAdder FullAdder_3420 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3420_io_a),
    .io_b(FullAdder_3420_io_b),
    .io_ci(FullAdder_3420_io_ci),
    .io_s(FullAdder_3420_io_s),
    .io_co(FullAdder_3420_io_co)
  );
  FullAdder FullAdder_3421 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3421_io_a),
    .io_b(FullAdder_3421_io_b),
    .io_ci(FullAdder_3421_io_ci),
    .io_s(FullAdder_3421_io_s),
    .io_co(FullAdder_3421_io_co)
  );
  FullAdder FullAdder_3422 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3422_io_a),
    .io_b(FullAdder_3422_io_b),
    .io_ci(FullAdder_3422_io_ci),
    .io_s(FullAdder_3422_io_s),
    .io_co(FullAdder_3422_io_co)
  );
  FullAdder FullAdder_3423 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3423_io_a),
    .io_b(FullAdder_3423_io_b),
    .io_ci(FullAdder_3423_io_ci),
    .io_s(FullAdder_3423_io_s),
    .io_co(FullAdder_3423_io_co)
  );
  HalfAdder HalfAdder_134 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_134_io_a),
    .io_b(HalfAdder_134_io_b),
    .io_s(HalfAdder_134_io_s),
    .io_co(HalfAdder_134_io_co)
  );
  FullAdder FullAdder_3424 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3424_io_a),
    .io_b(FullAdder_3424_io_b),
    .io_ci(FullAdder_3424_io_ci),
    .io_s(FullAdder_3424_io_s),
    .io_co(FullAdder_3424_io_co)
  );
  HalfAdder HalfAdder_135 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_135_io_a),
    .io_b(HalfAdder_135_io_b),
    .io_s(HalfAdder_135_io_s),
    .io_co(HalfAdder_135_io_co)
  );
  FullAdder FullAdder_3425 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3425_io_a),
    .io_b(FullAdder_3425_io_b),
    .io_ci(FullAdder_3425_io_ci),
    .io_s(FullAdder_3425_io_s),
    .io_co(FullAdder_3425_io_co)
  );
  HalfAdder HalfAdder_136 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_136_io_a),
    .io_b(HalfAdder_136_io_b),
    .io_s(HalfAdder_136_io_s),
    .io_co(HalfAdder_136_io_co)
  );
  FullAdder FullAdder_3426 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3426_io_a),
    .io_b(FullAdder_3426_io_b),
    .io_ci(FullAdder_3426_io_ci),
    .io_s(FullAdder_3426_io_s),
    .io_co(FullAdder_3426_io_co)
  );
  FullAdder FullAdder_3427 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3427_io_a),
    .io_b(FullAdder_3427_io_b),
    .io_ci(FullAdder_3427_io_ci),
    .io_s(FullAdder_3427_io_s),
    .io_co(FullAdder_3427_io_co)
  );
  FullAdder FullAdder_3428 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3428_io_a),
    .io_b(FullAdder_3428_io_b),
    .io_ci(FullAdder_3428_io_ci),
    .io_s(FullAdder_3428_io_s),
    .io_co(FullAdder_3428_io_co)
  );
  FullAdder FullAdder_3429 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3429_io_a),
    .io_b(FullAdder_3429_io_b),
    .io_ci(FullAdder_3429_io_ci),
    .io_s(FullAdder_3429_io_s),
    .io_co(FullAdder_3429_io_co)
  );
  FullAdder FullAdder_3430 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3430_io_a),
    .io_b(FullAdder_3430_io_b),
    .io_ci(FullAdder_3430_io_ci),
    .io_s(FullAdder_3430_io_s),
    .io_co(FullAdder_3430_io_co)
  );
  FullAdder FullAdder_3431 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3431_io_a),
    .io_b(FullAdder_3431_io_b),
    .io_ci(FullAdder_3431_io_ci),
    .io_s(FullAdder_3431_io_s),
    .io_co(FullAdder_3431_io_co)
  );
  FullAdder FullAdder_3432 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3432_io_a),
    .io_b(FullAdder_3432_io_b),
    .io_ci(FullAdder_3432_io_ci),
    .io_s(FullAdder_3432_io_s),
    .io_co(FullAdder_3432_io_co)
  );
  FullAdder FullAdder_3433 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3433_io_a),
    .io_b(FullAdder_3433_io_b),
    .io_ci(FullAdder_3433_io_ci),
    .io_s(FullAdder_3433_io_s),
    .io_co(FullAdder_3433_io_co)
  );
  FullAdder FullAdder_3434 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3434_io_a),
    .io_b(FullAdder_3434_io_b),
    .io_ci(FullAdder_3434_io_ci),
    .io_s(FullAdder_3434_io_s),
    .io_co(FullAdder_3434_io_co)
  );
  HalfAdder HalfAdder_137 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_137_io_a),
    .io_b(HalfAdder_137_io_b),
    .io_s(HalfAdder_137_io_s),
    .io_co(HalfAdder_137_io_co)
  );
  HalfAdder HalfAdder_138 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_138_io_a),
    .io_b(HalfAdder_138_io_b),
    .io_s(HalfAdder_138_io_s),
    .io_co(HalfAdder_138_io_co)
  );
  HalfAdder HalfAdder_139 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_139_io_a),
    .io_b(HalfAdder_139_io_b),
    .io_s(HalfAdder_139_io_s),
    .io_co(HalfAdder_139_io_co)
  );
  HalfAdder HalfAdder_140 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_140_io_a),
    .io_b(HalfAdder_140_io_b),
    .io_s(HalfAdder_140_io_s),
    .io_co(HalfAdder_140_io_co)
  );
  HalfAdder HalfAdder_141 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_141_io_a),
    .io_b(HalfAdder_141_io_b),
    .io_s(HalfAdder_141_io_s),
    .io_co(HalfAdder_141_io_co)
  );
  HalfAdder HalfAdder_142 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_142_io_a),
    .io_b(HalfAdder_142_io_b),
    .io_s(HalfAdder_142_io_s),
    .io_co(HalfAdder_142_io_co)
  );
  HalfAdder HalfAdder_143 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_143_io_a),
    .io_b(HalfAdder_143_io_b),
    .io_s(HalfAdder_143_io_s),
    .io_co(HalfAdder_143_io_co)
  );
  HalfAdder HalfAdder_144 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_144_io_a),
    .io_b(HalfAdder_144_io_b),
    .io_s(HalfAdder_144_io_s),
    .io_co(HalfAdder_144_io_co)
  );
  HalfAdder HalfAdder_145 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_145_io_a),
    .io_b(HalfAdder_145_io_b),
    .io_s(HalfAdder_145_io_s),
    .io_co(HalfAdder_145_io_co)
  );
  HalfAdder HalfAdder_146 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_146_io_a),
    .io_b(HalfAdder_146_io_b),
    .io_s(HalfAdder_146_io_s),
    .io_co(HalfAdder_146_io_co)
  );
  HalfAdder HalfAdder_147 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_147_io_a),
    .io_b(HalfAdder_147_io_b),
    .io_s(HalfAdder_147_io_s),
    .io_co(HalfAdder_147_io_co)
  );
  HalfAdder HalfAdder_148 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_148_io_a),
    .io_b(HalfAdder_148_io_b),
    .io_s(HalfAdder_148_io_s),
    .io_co(HalfAdder_148_io_co)
  );
  HalfAdder HalfAdder_149 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_149_io_a),
    .io_b(HalfAdder_149_io_b),
    .io_s(HalfAdder_149_io_s),
    .io_co(HalfAdder_149_io_co)
  );
  FullAdder FullAdder_3435 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3435_io_a),
    .io_b(FullAdder_3435_io_b),
    .io_ci(FullAdder_3435_io_ci),
    .io_s(FullAdder_3435_io_s),
    .io_co(FullAdder_3435_io_co)
  );
  HalfAdder HalfAdder_150 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_150_io_a),
    .io_b(HalfAdder_150_io_b),
    .io_s(HalfAdder_150_io_s),
    .io_co(HalfAdder_150_io_co)
  );
  FullAdder FullAdder_3436 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3436_io_a),
    .io_b(FullAdder_3436_io_b),
    .io_ci(FullAdder_3436_io_ci),
    .io_s(FullAdder_3436_io_s),
    .io_co(FullAdder_3436_io_co)
  );
  FullAdder FullAdder_3437 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3437_io_a),
    .io_b(FullAdder_3437_io_b),
    .io_ci(FullAdder_3437_io_ci),
    .io_s(FullAdder_3437_io_s),
    .io_co(FullAdder_3437_io_co)
  );
  FullAdder FullAdder_3438 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3438_io_a),
    .io_b(FullAdder_3438_io_b),
    .io_ci(FullAdder_3438_io_ci),
    .io_s(FullAdder_3438_io_s),
    .io_co(FullAdder_3438_io_co)
  );
  FullAdder FullAdder_3439 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3439_io_a),
    .io_b(FullAdder_3439_io_b),
    .io_ci(FullAdder_3439_io_ci),
    .io_s(FullAdder_3439_io_s),
    .io_co(FullAdder_3439_io_co)
  );
  FullAdder FullAdder_3440 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3440_io_a),
    .io_b(FullAdder_3440_io_b),
    .io_ci(FullAdder_3440_io_ci),
    .io_s(FullAdder_3440_io_s),
    .io_co(FullAdder_3440_io_co)
  );
  FullAdder FullAdder_3441 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3441_io_a),
    .io_b(FullAdder_3441_io_b),
    .io_ci(FullAdder_3441_io_ci),
    .io_s(FullAdder_3441_io_s),
    .io_co(FullAdder_3441_io_co)
  );
  FullAdder FullAdder_3442 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3442_io_a),
    .io_b(FullAdder_3442_io_b),
    .io_ci(FullAdder_3442_io_ci),
    .io_s(FullAdder_3442_io_s),
    .io_co(FullAdder_3442_io_co)
  );
  FullAdder FullAdder_3443 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3443_io_a),
    .io_b(FullAdder_3443_io_b),
    .io_ci(FullAdder_3443_io_ci),
    .io_s(FullAdder_3443_io_s),
    .io_co(FullAdder_3443_io_co)
  );
  FullAdder FullAdder_3444 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3444_io_a),
    .io_b(FullAdder_3444_io_b),
    .io_ci(FullAdder_3444_io_ci),
    .io_s(FullAdder_3444_io_s),
    .io_co(FullAdder_3444_io_co)
  );
  FullAdder FullAdder_3445 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3445_io_a),
    .io_b(FullAdder_3445_io_b),
    .io_ci(FullAdder_3445_io_ci),
    .io_s(FullAdder_3445_io_s),
    .io_co(FullAdder_3445_io_co)
  );
  FullAdder FullAdder_3446 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3446_io_a),
    .io_b(FullAdder_3446_io_b),
    .io_ci(FullAdder_3446_io_ci),
    .io_s(FullAdder_3446_io_s),
    .io_co(FullAdder_3446_io_co)
  );
  FullAdder FullAdder_3447 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3447_io_a),
    .io_b(FullAdder_3447_io_b),
    .io_ci(FullAdder_3447_io_ci),
    .io_s(FullAdder_3447_io_s),
    .io_co(FullAdder_3447_io_co)
  );
  FullAdder FullAdder_3448 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3448_io_a),
    .io_b(FullAdder_3448_io_b),
    .io_ci(FullAdder_3448_io_ci),
    .io_s(FullAdder_3448_io_s),
    .io_co(FullAdder_3448_io_co)
  );
  FullAdder FullAdder_3449 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3449_io_a),
    .io_b(FullAdder_3449_io_b),
    .io_ci(FullAdder_3449_io_ci),
    .io_s(FullAdder_3449_io_s),
    .io_co(FullAdder_3449_io_co)
  );
  HalfAdder HalfAdder_151 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_151_io_a),
    .io_b(HalfAdder_151_io_b),
    .io_s(HalfAdder_151_io_s),
    .io_co(HalfAdder_151_io_co)
  );
  HalfAdder HalfAdder_152 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_152_io_a),
    .io_b(HalfAdder_152_io_b),
    .io_s(HalfAdder_152_io_s),
    .io_co(HalfAdder_152_io_co)
  );
  FullAdder FullAdder_3450 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3450_io_a),
    .io_b(FullAdder_3450_io_b),
    .io_ci(FullAdder_3450_io_ci),
    .io_s(FullAdder_3450_io_s),
    .io_co(FullAdder_3450_io_co)
  );
  FullAdder FullAdder_3451 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3451_io_a),
    .io_b(FullAdder_3451_io_b),
    .io_ci(FullAdder_3451_io_ci),
    .io_s(FullAdder_3451_io_s),
    .io_co(FullAdder_3451_io_co)
  );
  FullAdder FullAdder_3452 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3452_io_a),
    .io_b(FullAdder_3452_io_b),
    .io_ci(FullAdder_3452_io_ci),
    .io_s(FullAdder_3452_io_s),
    .io_co(FullAdder_3452_io_co)
  );
  FullAdder FullAdder_3453 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3453_io_a),
    .io_b(FullAdder_3453_io_b),
    .io_ci(FullAdder_3453_io_ci),
    .io_s(FullAdder_3453_io_s),
    .io_co(FullAdder_3453_io_co)
  );
  FullAdder FullAdder_3454 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3454_io_a),
    .io_b(FullAdder_3454_io_b),
    .io_ci(FullAdder_3454_io_ci),
    .io_s(FullAdder_3454_io_s),
    .io_co(FullAdder_3454_io_co)
  );
  HalfAdder HalfAdder_153 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_153_io_a),
    .io_b(HalfAdder_153_io_b),
    .io_s(HalfAdder_153_io_s),
    .io_co(HalfAdder_153_io_co)
  );
  FullAdder FullAdder_3455 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3455_io_a),
    .io_b(FullAdder_3455_io_b),
    .io_ci(FullAdder_3455_io_ci),
    .io_s(FullAdder_3455_io_s),
    .io_co(FullAdder_3455_io_co)
  );
  FullAdder FullAdder_3456 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3456_io_a),
    .io_b(FullAdder_3456_io_b),
    .io_ci(FullAdder_3456_io_ci),
    .io_s(FullAdder_3456_io_s),
    .io_co(FullAdder_3456_io_co)
  );
  FullAdder FullAdder_3457 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3457_io_a),
    .io_b(FullAdder_3457_io_b),
    .io_ci(FullAdder_3457_io_ci),
    .io_s(FullAdder_3457_io_s),
    .io_co(FullAdder_3457_io_co)
  );
  FullAdder FullAdder_3458 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3458_io_a),
    .io_b(FullAdder_3458_io_b),
    .io_ci(FullAdder_3458_io_ci),
    .io_s(FullAdder_3458_io_s),
    .io_co(FullAdder_3458_io_co)
  );
  FullAdder FullAdder_3459 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3459_io_a),
    .io_b(FullAdder_3459_io_b),
    .io_ci(FullAdder_3459_io_ci),
    .io_s(FullAdder_3459_io_s),
    .io_co(FullAdder_3459_io_co)
  );
  HalfAdder HalfAdder_154 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_154_io_a),
    .io_b(HalfAdder_154_io_b),
    .io_s(HalfAdder_154_io_s),
    .io_co(HalfAdder_154_io_co)
  );
  FullAdder FullAdder_3460 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3460_io_a),
    .io_b(FullAdder_3460_io_b),
    .io_ci(FullAdder_3460_io_ci),
    .io_s(FullAdder_3460_io_s),
    .io_co(FullAdder_3460_io_co)
  );
  FullAdder FullAdder_3461 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3461_io_a),
    .io_b(FullAdder_3461_io_b),
    .io_ci(FullAdder_3461_io_ci),
    .io_s(FullAdder_3461_io_s),
    .io_co(FullAdder_3461_io_co)
  );
  FullAdder FullAdder_3462 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3462_io_a),
    .io_b(FullAdder_3462_io_b),
    .io_ci(FullAdder_3462_io_ci),
    .io_s(FullAdder_3462_io_s),
    .io_co(FullAdder_3462_io_co)
  );
  FullAdder FullAdder_3463 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3463_io_a),
    .io_b(FullAdder_3463_io_b),
    .io_ci(FullAdder_3463_io_ci),
    .io_s(FullAdder_3463_io_s),
    .io_co(FullAdder_3463_io_co)
  );
  FullAdder FullAdder_3464 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3464_io_a),
    .io_b(FullAdder_3464_io_b),
    .io_ci(FullAdder_3464_io_ci),
    .io_s(FullAdder_3464_io_s),
    .io_co(FullAdder_3464_io_co)
  );
  FullAdder FullAdder_3465 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3465_io_a),
    .io_b(FullAdder_3465_io_b),
    .io_ci(FullAdder_3465_io_ci),
    .io_s(FullAdder_3465_io_s),
    .io_co(FullAdder_3465_io_co)
  );
  FullAdder FullAdder_3466 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3466_io_a),
    .io_b(FullAdder_3466_io_b),
    .io_ci(FullAdder_3466_io_ci),
    .io_s(FullAdder_3466_io_s),
    .io_co(FullAdder_3466_io_co)
  );
  HalfAdder HalfAdder_155 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_155_io_a),
    .io_b(HalfAdder_155_io_b),
    .io_s(HalfAdder_155_io_s),
    .io_co(HalfAdder_155_io_co)
  );
  HalfAdder HalfAdder_156 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_156_io_a),
    .io_b(HalfAdder_156_io_b),
    .io_s(HalfAdder_156_io_s),
    .io_co(HalfAdder_156_io_co)
  );
  HalfAdder HalfAdder_157 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_157_io_a),
    .io_b(HalfAdder_157_io_b),
    .io_s(HalfAdder_157_io_s),
    .io_co(HalfAdder_157_io_co)
  );
  FullAdder FullAdder_3467 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3467_io_a),
    .io_b(FullAdder_3467_io_b),
    .io_ci(FullAdder_3467_io_ci),
    .io_s(FullAdder_3467_io_s),
    .io_co(FullAdder_3467_io_co)
  );
  FullAdder FullAdder_3468 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3468_io_a),
    .io_b(FullAdder_3468_io_b),
    .io_ci(FullAdder_3468_io_ci),
    .io_s(FullAdder_3468_io_s),
    .io_co(FullAdder_3468_io_co)
  );
  FullAdder FullAdder_3469 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3469_io_a),
    .io_b(FullAdder_3469_io_b),
    .io_ci(FullAdder_3469_io_ci),
    .io_s(FullAdder_3469_io_s),
    .io_co(FullAdder_3469_io_co)
  );
  FullAdder FullAdder_3470 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3470_io_a),
    .io_b(FullAdder_3470_io_b),
    .io_ci(FullAdder_3470_io_ci),
    .io_s(FullAdder_3470_io_s),
    .io_co(FullAdder_3470_io_co)
  );
  FullAdder FullAdder_3471 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3471_io_a),
    .io_b(FullAdder_3471_io_b),
    .io_ci(FullAdder_3471_io_ci),
    .io_s(FullAdder_3471_io_s),
    .io_co(FullAdder_3471_io_co)
  );
  FullAdder FullAdder_3472 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3472_io_a),
    .io_b(FullAdder_3472_io_b),
    .io_ci(FullAdder_3472_io_ci),
    .io_s(FullAdder_3472_io_s),
    .io_co(FullAdder_3472_io_co)
  );
  FullAdder FullAdder_3473 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3473_io_a),
    .io_b(FullAdder_3473_io_b),
    .io_ci(FullAdder_3473_io_ci),
    .io_s(FullAdder_3473_io_s),
    .io_co(FullAdder_3473_io_co)
  );
  FullAdder FullAdder_3474 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3474_io_a),
    .io_b(FullAdder_3474_io_b),
    .io_ci(FullAdder_3474_io_ci),
    .io_s(FullAdder_3474_io_s),
    .io_co(FullAdder_3474_io_co)
  );
  FullAdder FullAdder_3475 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3475_io_a),
    .io_b(FullAdder_3475_io_b),
    .io_ci(FullAdder_3475_io_ci),
    .io_s(FullAdder_3475_io_s),
    .io_co(FullAdder_3475_io_co)
  );
  FullAdder FullAdder_3476 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3476_io_a),
    .io_b(FullAdder_3476_io_b),
    .io_ci(FullAdder_3476_io_ci),
    .io_s(FullAdder_3476_io_s),
    .io_co(FullAdder_3476_io_co)
  );
  FullAdder FullAdder_3477 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3477_io_a),
    .io_b(FullAdder_3477_io_b),
    .io_ci(FullAdder_3477_io_ci),
    .io_s(FullAdder_3477_io_s),
    .io_co(FullAdder_3477_io_co)
  );
  FullAdder FullAdder_3478 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3478_io_a),
    .io_b(FullAdder_3478_io_b),
    .io_ci(FullAdder_3478_io_ci),
    .io_s(FullAdder_3478_io_s),
    .io_co(FullAdder_3478_io_co)
  );
  FullAdder FullAdder_3479 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3479_io_a),
    .io_b(FullAdder_3479_io_b),
    .io_ci(FullAdder_3479_io_ci),
    .io_s(FullAdder_3479_io_s),
    .io_co(FullAdder_3479_io_co)
  );
  FullAdder FullAdder_3480 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3480_io_a),
    .io_b(FullAdder_3480_io_b),
    .io_ci(FullAdder_3480_io_ci),
    .io_s(FullAdder_3480_io_s),
    .io_co(FullAdder_3480_io_co)
  );
  FullAdder FullAdder_3481 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3481_io_a),
    .io_b(FullAdder_3481_io_b),
    .io_ci(FullAdder_3481_io_ci),
    .io_s(FullAdder_3481_io_s),
    .io_co(FullAdder_3481_io_co)
  );
  FullAdder FullAdder_3482 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3482_io_a),
    .io_b(FullAdder_3482_io_b),
    .io_ci(FullAdder_3482_io_ci),
    .io_s(FullAdder_3482_io_s),
    .io_co(FullAdder_3482_io_co)
  );
  FullAdder FullAdder_3483 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3483_io_a),
    .io_b(FullAdder_3483_io_b),
    .io_ci(FullAdder_3483_io_ci),
    .io_s(FullAdder_3483_io_s),
    .io_co(FullAdder_3483_io_co)
  );
  FullAdder FullAdder_3484 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3484_io_a),
    .io_b(FullAdder_3484_io_b),
    .io_ci(FullAdder_3484_io_ci),
    .io_s(FullAdder_3484_io_s),
    .io_co(FullAdder_3484_io_co)
  );
  HalfAdder HalfAdder_158 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_158_io_a),
    .io_b(HalfAdder_158_io_b),
    .io_s(HalfAdder_158_io_s),
    .io_co(HalfAdder_158_io_co)
  );
  FullAdder FullAdder_3485 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3485_io_a),
    .io_b(FullAdder_3485_io_b),
    .io_ci(FullAdder_3485_io_ci),
    .io_s(FullAdder_3485_io_s),
    .io_co(FullAdder_3485_io_co)
  );
  FullAdder FullAdder_3486 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3486_io_a),
    .io_b(FullAdder_3486_io_b),
    .io_ci(FullAdder_3486_io_ci),
    .io_s(FullAdder_3486_io_s),
    .io_co(FullAdder_3486_io_co)
  );
  FullAdder FullAdder_3487 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3487_io_a),
    .io_b(FullAdder_3487_io_b),
    .io_ci(FullAdder_3487_io_ci),
    .io_s(FullAdder_3487_io_s),
    .io_co(FullAdder_3487_io_co)
  );
  FullAdder FullAdder_3488 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3488_io_a),
    .io_b(FullAdder_3488_io_b),
    .io_ci(FullAdder_3488_io_ci),
    .io_s(FullAdder_3488_io_s),
    .io_co(FullAdder_3488_io_co)
  );
  FullAdder FullAdder_3489 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3489_io_a),
    .io_b(FullAdder_3489_io_b),
    .io_ci(FullAdder_3489_io_ci),
    .io_s(FullAdder_3489_io_s),
    .io_co(FullAdder_3489_io_co)
  );
  FullAdder FullAdder_3490 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3490_io_a),
    .io_b(FullAdder_3490_io_b),
    .io_ci(FullAdder_3490_io_ci),
    .io_s(FullAdder_3490_io_s),
    .io_co(FullAdder_3490_io_co)
  );
  HalfAdder HalfAdder_159 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_159_io_a),
    .io_b(HalfAdder_159_io_b),
    .io_s(HalfAdder_159_io_s),
    .io_co(HalfAdder_159_io_co)
  );
  FullAdder FullAdder_3491 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3491_io_a),
    .io_b(FullAdder_3491_io_b),
    .io_ci(FullAdder_3491_io_ci),
    .io_s(FullAdder_3491_io_s),
    .io_co(FullAdder_3491_io_co)
  );
  FullAdder FullAdder_3492 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3492_io_a),
    .io_b(FullAdder_3492_io_b),
    .io_ci(FullAdder_3492_io_ci),
    .io_s(FullAdder_3492_io_s),
    .io_co(FullAdder_3492_io_co)
  );
  FullAdder FullAdder_3493 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3493_io_a),
    .io_b(FullAdder_3493_io_b),
    .io_ci(FullAdder_3493_io_ci),
    .io_s(FullAdder_3493_io_s),
    .io_co(FullAdder_3493_io_co)
  );
  FullAdder FullAdder_3494 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3494_io_a),
    .io_b(FullAdder_3494_io_b),
    .io_ci(FullAdder_3494_io_ci),
    .io_s(FullAdder_3494_io_s),
    .io_co(FullAdder_3494_io_co)
  );
  HalfAdder HalfAdder_160 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_160_io_a),
    .io_b(HalfAdder_160_io_b),
    .io_s(HalfAdder_160_io_s),
    .io_co(HalfAdder_160_io_co)
  );
  FullAdder FullAdder_3495 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3495_io_a),
    .io_b(FullAdder_3495_io_b),
    .io_ci(FullAdder_3495_io_ci),
    .io_s(FullAdder_3495_io_s),
    .io_co(FullAdder_3495_io_co)
  );
  FullAdder FullAdder_3496 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3496_io_a),
    .io_b(FullAdder_3496_io_b),
    .io_ci(FullAdder_3496_io_ci),
    .io_s(FullAdder_3496_io_s),
    .io_co(FullAdder_3496_io_co)
  );
  HalfAdder HalfAdder_161 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_161_io_a),
    .io_b(HalfAdder_161_io_b),
    .io_s(HalfAdder_161_io_s),
    .io_co(HalfAdder_161_io_co)
  );
  FullAdder FullAdder_3497 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3497_io_a),
    .io_b(FullAdder_3497_io_b),
    .io_ci(FullAdder_3497_io_ci),
    .io_s(FullAdder_3497_io_s),
    .io_co(FullAdder_3497_io_co)
  );
  FullAdder FullAdder_3498 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3498_io_a),
    .io_b(FullAdder_3498_io_b),
    .io_ci(FullAdder_3498_io_ci),
    .io_s(FullAdder_3498_io_s),
    .io_co(FullAdder_3498_io_co)
  );
  FullAdder FullAdder_3499 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3499_io_a),
    .io_b(FullAdder_3499_io_b),
    .io_ci(FullAdder_3499_io_ci),
    .io_s(FullAdder_3499_io_s),
    .io_co(FullAdder_3499_io_co)
  );
  FullAdder FullAdder_3500 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3500_io_a),
    .io_b(FullAdder_3500_io_b),
    .io_ci(FullAdder_3500_io_ci),
    .io_s(FullAdder_3500_io_s),
    .io_co(FullAdder_3500_io_co)
  );
  FullAdder FullAdder_3501 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3501_io_a),
    .io_b(FullAdder_3501_io_b),
    .io_ci(FullAdder_3501_io_ci),
    .io_s(FullAdder_3501_io_s),
    .io_co(FullAdder_3501_io_co)
  );
  FullAdder FullAdder_3502 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3502_io_a),
    .io_b(FullAdder_3502_io_b),
    .io_ci(FullAdder_3502_io_ci),
    .io_s(FullAdder_3502_io_s),
    .io_co(FullAdder_3502_io_co)
  );
  FullAdder FullAdder_3503 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3503_io_a),
    .io_b(FullAdder_3503_io_b),
    .io_ci(FullAdder_3503_io_ci),
    .io_s(FullAdder_3503_io_s),
    .io_co(FullAdder_3503_io_co)
  );
  FullAdder FullAdder_3504 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3504_io_a),
    .io_b(FullAdder_3504_io_b),
    .io_ci(FullAdder_3504_io_ci),
    .io_s(FullAdder_3504_io_s),
    .io_co(FullAdder_3504_io_co)
  );
  HalfAdder HalfAdder_162 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_162_io_a),
    .io_b(HalfAdder_162_io_b),
    .io_s(HalfAdder_162_io_s),
    .io_co(HalfAdder_162_io_co)
  );
  FullAdder FullAdder_3505 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3505_io_a),
    .io_b(FullAdder_3505_io_b),
    .io_ci(FullAdder_3505_io_ci),
    .io_s(FullAdder_3505_io_s),
    .io_co(FullAdder_3505_io_co)
  );
  FullAdder FullAdder_3506 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3506_io_a),
    .io_b(FullAdder_3506_io_b),
    .io_ci(FullAdder_3506_io_ci),
    .io_s(FullAdder_3506_io_s),
    .io_co(FullAdder_3506_io_co)
  );
  HalfAdder HalfAdder_163 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_163_io_a),
    .io_b(HalfAdder_163_io_b),
    .io_s(HalfAdder_163_io_s),
    .io_co(HalfAdder_163_io_co)
  );
  FullAdder FullAdder_3507 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3507_io_a),
    .io_b(FullAdder_3507_io_b),
    .io_ci(FullAdder_3507_io_ci),
    .io_s(FullAdder_3507_io_s),
    .io_co(FullAdder_3507_io_co)
  );
  HalfAdder HalfAdder_164 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_164_io_a),
    .io_b(HalfAdder_164_io_b),
    .io_s(HalfAdder_164_io_s),
    .io_co(HalfAdder_164_io_co)
  );
  HalfAdder HalfAdder_165 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_165_io_a),
    .io_b(HalfAdder_165_io_b),
    .io_s(HalfAdder_165_io_s),
    .io_co(HalfAdder_165_io_co)
  );
  HalfAdder HalfAdder_166 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_166_io_a),
    .io_b(HalfAdder_166_io_b),
    .io_s(HalfAdder_166_io_s),
    .io_co(HalfAdder_166_io_co)
  );
  FullAdder FullAdder_3508 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3508_io_a),
    .io_b(FullAdder_3508_io_b),
    .io_ci(FullAdder_3508_io_ci),
    .io_s(FullAdder_3508_io_s),
    .io_co(FullAdder_3508_io_co)
  );
  FullAdder FullAdder_3509 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3509_io_a),
    .io_b(FullAdder_3509_io_b),
    .io_ci(FullAdder_3509_io_ci),
    .io_s(FullAdder_3509_io_s),
    .io_co(FullAdder_3509_io_co)
  );
  FullAdder FullAdder_3510 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3510_io_a),
    .io_b(FullAdder_3510_io_b),
    .io_ci(FullAdder_3510_io_ci),
    .io_s(FullAdder_3510_io_s),
    .io_co(FullAdder_3510_io_co)
  );
  FullAdder FullAdder_3511 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3511_io_a),
    .io_b(FullAdder_3511_io_b),
    .io_ci(FullAdder_3511_io_ci),
    .io_s(FullAdder_3511_io_s),
    .io_co(FullAdder_3511_io_co)
  );
  FullAdder FullAdder_3512 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3512_io_a),
    .io_b(FullAdder_3512_io_b),
    .io_ci(FullAdder_3512_io_ci),
    .io_s(FullAdder_3512_io_s),
    .io_co(FullAdder_3512_io_co)
  );
  FullAdder FullAdder_3513 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3513_io_a),
    .io_b(FullAdder_3513_io_b),
    .io_ci(FullAdder_3513_io_ci),
    .io_s(FullAdder_3513_io_s),
    .io_co(FullAdder_3513_io_co)
  );
  FullAdder FullAdder_3514 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3514_io_a),
    .io_b(FullAdder_3514_io_b),
    .io_ci(FullAdder_3514_io_ci),
    .io_s(FullAdder_3514_io_s),
    .io_co(FullAdder_3514_io_co)
  );
  FullAdder FullAdder_3515 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3515_io_a),
    .io_b(FullAdder_3515_io_b),
    .io_ci(FullAdder_3515_io_ci),
    .io_s(FullAdder_3515_io_s),
    .io_co(FullAdder_3515_io_co)
  );
  FullAdder FullAdder_3516 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3516_io_a),
    .io_b(FullAdder_3516_io_b),
    .io_ci(FullAdder_3516_io_ci),
    .io_s(FullAdder_3516_io_s),
    .io_co(FullAdder_3516_io_co)
  );
  FullAdder FullAdder_3517 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3517_io_a),
    .io_b(FullAdder_3517_io_b),
    .io_ci(FullAdder_3517_io_ci),
    .io_s(FullAdder_3517_io_s),
    .io_co(FullAdder_3517_io_co)
  );
  FullAdder FullAdder_3518 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3518_io_a),
    .io_b(FullAdder_3518_io_b),
    .io_ci(FullAdder_3518_io_ci),
    .io_s(FullAdder_3518_io_s),
    .io_co(FullAdder_3518_io_co)
  );
  FullAdder FullAdder_3519 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3519_io_a),
    .io_b(FullAdder_3519_io_b),
    .io_ci(FullAdder_3519_io_ci),
    .io_s(FullAdder_3519_io_s),
    .io_co(FullAdder_3519_io_co)
  );
  FullAdder FullAdder_3520 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3520_io_a),
    .io_b(FullAdder_3520_io_b),
    .io_ci(FullAdder_3520_io_ci),
    .io_s(FullAdder_3520_io_s),
    .io_co(FullAdder_3520_io_co)
  );
  FullAdder FullAdder_3521 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3521_io_a),
    .io_b(FullAdder_3521_io_b),
    .io_ci(FullAdder_3521_io_ci),
    .io_s(FullAdder_3521_io_s),
    .io_co(FullAdder_3521_io_co)
  );
  FullAdder FullAdder_3522 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3522_io_a),
    .io_b(FullAdder_3522_io_b),
    .io_ci(FullAdder_3522_io_ci),
    .io_s(FullAdder_3522_io_s),
    .io_co(FullAdder_3522_io_co)
  );
  FullAdder FullAdder_3523 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3523_io_a),
    .io_b(FullAdder_3523_io_b),
    .io_ci(FullAdder_3523_io_ci),
    .io_s(FullAdder_3523_io_s),
    .io_co(FullAdder_3523_io_co)
  );
  FullAdder FullAdder_3524 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3524_io_a),
    .io_b(FullAdder_3524_io_b),
    .io_ci(FullAdder_3524_io_ci),
    .io_s(FullAdder_3524_io_s),
    .io_co(FullAdder_3524_io_co)
  );
  FullAdder FullAdder_3525 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3525_io_a),
    .io_b(FullAdder_3525_io_b),
    .io_ci(FullAdder_3525_io_ci),
    .io_s(FullAdder_3525_io_s),
    .io_co(FullAdder_3525_io_co)
  );
  FullAdder FullAdder_3526 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3526_io_a),
    .io_b(FullAdder_3526_io_b),
    .io_ci(FullAdder_3526_io_ci),
    .io_s(FullAdder_3526_io_s),
    .io_co(FullAdder_3526_io_co)
  );
  FullAdder FullAdder_3527 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3527_io_a),
    .io_b(FullAdder_3527_io_b),
    .io_ci(FullAdder_3527_io_ci),
    .io_s(FullAdder_3527_io_s),
    .io_co(FullAdder_3527_io_co)
  );
  FullAdder FullAdder_3528 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3528_io_a),
    .io_b(FullAdder_3528_io_b),
    .io_ci(FullAdder_3528_io_ci),
    .io_s(FullAdder_3528_io_s),
    .io_co(FullAdder_3528_io_co)
  );
  FullAdder FullAdder_3529 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3529_io_a),
    .io_b(FullAdder_3529_io_b),
    .io_ci(FullAdder_3529_io_ci),
    .io_s(FullAdder_3529_io_s),
    .io_co(FullAdder_3529_io_co)
  );
  FullAdder FullAdder_3530 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3530_io_a),
    .io_b(FullAdder_3530_io_b),
    .io_ci(FullAdder_3530_io_ci),
    .io_s(FullAdder_3530_io_s),
    .io_co(FullAdder_3530_io_co)
  );
  FullAdder FullAdder_3531 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3531_io_a),
    .io_b(FullAdder_3531_io_b),
    .io_ci(FullAdder_3531_io_ci),
    .io_s(FullAdder_3531_io_s),
    .io_co(FullAdder_3531_io_co)
  );
  FullAdder FullAdder_3532 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3532_io_a),
    .io_b(FullAdder_3532_io_b),
    .io_ci(FullAdder_3532_io_ci),
    .io_s(FullAdder_3532_io_s),
    .io_co(FullAdder_3532_io_co)
  );
  FullAdder FullAdder_3533 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3533_io_a),
    .io_b(FullAdder_3533_io_b),
    .io_ci(FullAdder_3533_io_ci),
    .io_s(FullAdder_3533_io_s),
    .io_co(FullAdder_3533_io_co)
  );
  FullAdder FullAdder_3534 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3534_io_a),
    .io_b(FullAdder_3534_io_b),
    .io_ci(FullAdder_3534_io_ci),
    .io_s(FullAdder_3534_io_s),
    .io_co(FullAdder_3534_io_co)
  );
  HalfAdder HalfAdder_167 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_167_io_a),
    .io_b(HalfAdder_167_io_b),
    .io_s(HalfAdder_167_io_s),
    .io_co(HalfAdder_167_io_co)
  );
  FullAdder FullAdder_3535 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3535_io_a),
    .io_b(FullAdder_3535_io_b),
    .io_ci(FullAdder_3535_io_ci),
    .io_s(FullAdder_3535_io_s),
    .io_co(FullAdder_3535_io_co)
  );
  FullAdder FullAdder_3536 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3536_io_a),
    .io_b(FullAdder_3536_io_b),
    .io_ci(FullAdder_3536_io_ci),
    .io_s(FullAdder_3536_io_s),
    .io_co(FullAdder_3536_io_co)
  );
  FullAdder FullAdder_3537 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3537_io_a),
    .io_b(FullAdder_3537_io_b),
    .io_ci(FullAdder_3537_io_ci),
    .io_s(FullAdder_3537_io_s),
    .io_co(FullAdder_3537_io_co)
  );
  FullAdder FullAdder_3538 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3538_io_a),
    .io_b(FullAdder_3538_io_b),
    .io_ci(FullAdder_3538_io_ci),
    .io_s(FullAdder_3538_io_s),
    .io_co(FullAdder_3538_io_co)
  );
  FullAdder FullAdder_3539 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3539_io_a),
    .io_b(FullAdder_3539_io_b),
    .io_ci(FullAdder_3539_io_ci),
    .io_s(FullAdder_3539_io_s),
    .io_co(FullAdder_3539_io_co)
  );
  FullAdder FullAdder_3540 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3540_io_a),
    .io_b(FullAdder_3540_io_b),
    .io_ci(FullAdder_3540_io_ci),
    .io_s(FullAdder_3540_io_s),
    .io_co(FullAdder_3540_io_co)
  );
  FullAdder FullAdder_3541 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3541_io_a),
    .io_b(FullAdder_3541_io_b),
    .io_ci(FullAdder_3541_io_ci),
    .io_s(FullAdder_3541_io_s),
    .io_co(FullAdder_3541_io_co)
  );
  FullAdder FullAdder_3542 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3542_io_a),
    .io_b(FullAdder_3542_io_b),
    .io_ci(FullAdder_3542_io_ci),
    .io_s(FullAdder_3542_io_s),
    .io_co(FullAdder_3542_io_co)
  );
  FullAdder FullAdder_3543 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3543_io_a),
    .io_b(FullAdder_3543_io_b),
    .io_ci(FullAdder_3543_io_ci),
    .io_s(FullAdder_3543_io_s),
    .io_co(FullAdder_3543_io_co)
  );
  FullAdder FullAdder_3544 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3544_io_a),
    .io_b(FullAdder_3544_io_b),
    .io_ci(FullAdder_3544_io_ci),
    .io_s(FullAdder_3544_io_s),
    .io_co(FullAdder_3544_io_co)
  );
  FullAdder FullAdder_3545 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3545_io_a),
    .io_b(FullAdder_3545_io_b),
    .io_ci(FullAdder_3545_io_ci),
    .io_s(FullAdder_3545_io_s),
    .io_co(FullAdder_3545_io_co)
  );
  FullAdder FullAdder_3546 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3546_io_a),
    .io_b(FullAdder_3546_io_b),
    .io_ci(FullAdder_3546_io_ci),
    .io_s(FullAdder_3546_io_s),
    .io_co(FullAdder_3546_io_co)
  );
  FullAdder FullAdder_3547 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3547_io_a),
    .io_b(FullAdder_3547_io_b),
    .io_ci(FullAdder_3547_io_ci),
    .io_s(FullAdder_3547_io_s),
    .io_co(FullAdder_3547_io_co)
  );
  FullAdder FullAdder_3548 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3548_io_a),
    .io_b(FullAdder_3548_io_b),
    .io_ci(FullAdder_3548_io_ci),
    .io_s(FullAdder_3548_io_s),
    .io_co(FullAdder_3548_io_co)
  );
  FullAdder FullAdder_3549 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3549_io_a),
    .io_b(FullAdder_3549_io_b),
    .io_ci(FullAdder_3549_io_ci),
    .io_s(FullAdder_3549_io_s),
    .io_co(FullAdder_3549_io_co)
  );
  FullAdder FullAdder_3550 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3550_io_a),
    .io_b(FullAdder_3550_io_b),
    .io_ci(FullAdder_3550_io_ci),
    .io_s(FullAdder_3550_io_s),
    .io_co(FullAdder_3550_io_co)
  );
  FullAdder FullAdder_3551 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3551_io_a),
    .io_b(FullAdder_3551_io_b),
    .io_ci(FullAdder_3551_io_ci),
    .io_s(FullAdder_3551_io_s),
    .io_co(FullAdder_3551_io_co)
  );
  FullAdder FullAdder_3552 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3552_io_a),
    .io_b(FullAdder_3552_io_b),
    .io_ci(FullAdder_3552_io_ci),
    .io_s(FullAdder_3552_io_s),
    .io_co(FullAdder_3552_io_co)
  );
  FullAdder FullAdder_3553 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3553_io_a),
    .io_b(FullAdder_3553_io_b),
    .io_ci(FullAdder_3553_io_ci),
    .io_s(FullAdder_3553_io_s),
    .io_co(FullAdder_3553_io_co)
  );
  FullAdder FullAdder_3554 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3554_io_a),
    .io_b(FullAdder_3554_io_b),
    .io_ci(FullAdder_3554_io_ci),
    .io_s(FullAdder_3554_io_s),
    .io_co(FullAdder_3554_io_co)
  );
  FullAdder FullAdder_3555 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3555_io_a),
    .io_b(FullAdder_3555_io_b),
    .io_ci(FullAdder_3555_io_ci),
    .io_s(FullAdder_3555_io_s),
    .io_co(FullAdder_3555_io_co)
  );
  FullAdder FullAdder_3556 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3556_io_a),
    .io_b(FullAdder_3556_io_b),
    .io_ci(FullAdder_3556_io_ci),
    .io_s(FullAdder_3556_io_s),
    .io_co(FullAdder_3556_io_co)
  );
  FullAdder FullAdder_3557 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3557_io_a),
    .io_b(FullAdder_3557_io_b),
    .io_ci(FullAdder_3557_io_ci),
    .io_s(FullAdder_3557_io_s),
    .io_co(FullAdder_3557_io_co)
  );
  FullAdder FullAdder_3558 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3558_io_a),
    .io_b(FullAdder_3558_io_b),
    .io_ci(FullAdder_3558_io_ci),
    .io_s(FullAdder_3558_io_s),
    .io_co(FullAdder_3558_io_co)
  );
  FullAdder FullAdder_3559 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3559_io_a),
    .io_b(FullAdder_3559_io_b),
    .io_ci(FullAdder_3559_io_ci),
    .io_s(FullAdder_3559_io_s),
    .io_co(FullAdder_3559_io_co)
  );
  FullAdder FullAdder_3560 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3560_io_a),
    .io_b(FullAdder_3560_io_b),
    .io_ci(FullAdder_3560_io_ci),
    .io_s(FullAdder_3560_io_s),
    .io_co(FullAdder_3560_io_co)
  );
  FullAdder FullAdder_3561 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3561_io_a),
    .io_b(FullAdder_3561_io_b),
    .io_ci(FullAdder_3561_io_ci),
    .io_s(FullAdder_3561_io_s),
    .io_co(FullAdder_3561_io_co)
  );
  FullAdder FullAdder_3562 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3562_io_a),
    .io_b(FullAdder_3562_io_b),
    .io_ci(FullAdder_3562_io_ci),
    .io_s(FullAdder_3562_io_s),
    .io_co(FullAdder_3562_io_co)
  );
  FullAdder FullAdder_3563 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3563_io_a),
    .io_b(FullAdder_3563_io_b),
    .io_ci(FullAdder_3563_io_ci),
    .io_s(FullAdder_3563_io_s),
    .io_co(FullAdder_3563_io_co)
  );
  FullAdder FullAdder_3564 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3564_io_a),
    .io_b(FullAdder_3564_io_b),
    .io_ci(FullAdder_3564_io_ci),
    .io_s(FullAdder_3564_io_s),
    .io_co(FullAdder_3564_io_co)
  );
  FullAdder FullAdder_3565 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3565_io_a),
    .io_b(FullAdder_3565_io_b),
    .io_ci(FullAdder_3565_io_ci),
    .io_s(FullAdder_3565_io_s),
    .io_co(FullAdder_3565_io_co)
  );
  FullAdder FullAdder_3566 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3566_io_a),
    .io_b(FullAdder_3566_io_b),
    .io_ci(FullAdder_3566_io_ci),
    .io_s(FullAdder_3566_io_s),
    .io_co(FullAdder_3566_io_co)
  );
  HalfAdder HalfAdder_168 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_168_io_a),
    .io_b(HalfAdder_168_io_b),
    .io_s(HalfAdder_168_io_s),
    .io_co(HalfAdder_168_io_co)
  );
  FullAdder FullAdder_3567 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3567_io_a),
    .io_b(FullAdder_3567_io_b),
    .io_ci(FullAdder_3567_io_ci),
    .io_s(FullAdder_3567_io_s),
    .io_co(FullAdder_3567_io_co)
  );
  FullAdder FullAdder_3568 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3568_io_a),
    .io_b(FullAdder_3568_io_b),
    .io_ci(FullAdder_3568_io_ci),
    .io_s(FullAdder_3568_io_s),
    .io_co(FullAdder_3568_io_co)
  );
  FullAdder FullAdder_3569 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3569_io_a),
    .io_b(FullAdder_3569_io_b),
    .io_ci(FullAdder_3569_io_ci),
    .io_s(FullAdder_3569_io_s),
    .io_co(FullAdder_3569_io_co)
  );
  FullAdder FullAdder_3570 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3570_io_a),
    .io_b(FullAdder_3570_io_b),
    .io_ci(FullAdder_3570_io_ci),
    .io_s(FullAdder_3570_io_s),
    .io_co(FullAdder_3570_io_co)
  );
  FullAdder FullAdder_3571 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3571_io_a),
    .io_b(FullAdder_3571_io_b),
    .io_ci(FullAdder_3571_io_ci),
    .io_s(FullAdder_3571_io_s),
    .io_co(FullAdder_3571_io_co)
  );
  FullAdder FullAdder_3572 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3572_io_a),
    .io_b(FullAdder_3572_io_b),
    .io_ci(FullAdder_3572_io_ci),
    .io_s(FullAdder_3572_io_s),
    .io_co(FullAdder_3572_io_co)
  );
  FullAdder FullAdder_3573 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3573_io_a),
    .io_b(FullAdder_3573_io_b),
    .io_ci(FullAdder_3573_io_ci),
    .io_s(FullAdder_3573_io_s),
    .io_co(FullAdder_3573_io_co)
  );
  FullAdder FullAdder_3574 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3574_io_a),
    .io_b(FullAdder_3574_io_b),
    .io_ci(FullAdder_3574_io_ci),
    .io_s(FullAdder_3574_io_s),
    .io_co(FullAdder_3574_io_co)
  );
  FullAdder FullAdder_3575 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3575_io_a),
    .io_b(FullAdder_3575_io_b),
    .io_ci(FullAdder_3575_io_ci),
    .io_s(FullAdder_3575_io_s),
    .io_co(FullAdder_3575_io_co)
  );
  FullAdder FullAdder_3576 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3576_io_a),
    .io_b(FullAdder_3576_io_b),
    .io_ci(FullAdder_3576_io_ci),
    .io_s(FullAdder_3576_io_s),
    .io_co(FullAdder_3576_io_co)
  );
  HalfAdder HalfAdder_169 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_169_io_a),
    .io_b(HalfAdder_169_io_b),
    .io_s(HalfAdder_169_io_s),
    .io_co(HalfAdder_169_io_co)
  );
  FullAdder FullAdder_3577 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3577_io_a),
    .io_b(FullAdder_3577_io_b),
    .io_ci(FullAdder_3577_io_ci),
    .io_s(FullAdder_3577_io_s),
    .io_co(FullAdder_3577_io_co)
  );
  FullAdder FullAdder_3578 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3578_io_a),
    .io_b(FullAdder_3578_io_b),
    .io_ci(FullAdder_3578_io_ci),
    .io_s(FullAdder_3578_io_s),
    .io_co(FullAdder_3578_io_co)
  );
  HalfAdder HalfAdder_170 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_170_io_a),
    .io_b(HalfAdder_170_io_b),
    .io_s(HalfAdder_170_io_s),
    .io_co(HalfAdder_170_io_co)
  );
  FullAdder FullAdder_3579 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3579_io_a),
    .io_b(FullAdder_3579_io_b),
    .io_ci(FullAdder_3579_io_ci),
    .io_s(FullAdder_3579_io_s),
    .io_co(FullAdder_3579_io_co)
  );
  FullAdder FullAdder_3580 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3580_io_a),
    .io_b(FullAdder_3580_io_b),
    .io_ci(FullAdder_3580_io_ci),
    .io_s(FullAdder_3580_io_s),
    .io_co(FullAdder_3580_io_co)
  );
  FullAdder FullAdder_3581 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3581_io_a),
    .io_b(FullAdder_3581_io_b),
    .io_ci(FullAdder_3581_io_ci),
    .io_s(FullAdder_3581_io_s),
    .io_co(FullAdder_3581_io_co)
  );
  FullAdder FullAdder_3582 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3582_io_a),
    .io_b(FullAdder_3582_io_b),
    .io_ci(FullAdder_3582_io_ci),
    .io_s(FullAdder_3582_io_s),
    .io_co(FullAdder_3582_io_co)
  );
  FullAdder FullAdder_3583 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3583_io_a),
    .io_b(FullAdder_3583_io_b),
    .io_ci(FullAdder_3583_io_ci),
    .io_s(FullAdder_3583_io_s),
    .io_co(FullAdder_3583_io_co)
  );
  FullAdder FullAdder_3584 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3584_io_a),
    .io_b(FullAdder_3584_io_b),
    .io_ci(FullAdder_3584_io_ci),
    .io_s(FullAdder_3584_io_s),
    .io_co(FullAdder_3584_io_co)
  );
  FullAdder FullAdder_3585 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3585_io_a),
    .io_b(FullAdder_3585_io_b),
    .io_ci(FullAdder_3585_io_ci),
    .io_s(FullAdder_3585_io_s),
    .io_co(FullAdder_3585_io_co)
  );
  FullAdder FullAdder_3586 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3586_io_a),
    .io_b(FullAdder_3586_io_b),
    .io_ci(FullAdder_3586_io_ci),
    .io_s(FullAdder_3586_io_s),
    .io_co(FullAdder_3586_io_co)
  );
  FullAdder FullAdder_3587 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3587_io_a),
    .io_b(FullAdder_3587_io_b),
    .io_ci(FullAdder_3587_io_ci),
    .io_s(FullAdder_3587_io_s),
    .io_co(FullAdder_3587_io_co)
  );
  FullAdder FullAdder_3588 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3588_io_a),
    .io_b(FullAdder_3588_io_b),
    .io_ci(FullAdder_3588_io_ci),
    .io_s(FullAdder_3588_io_s),
    .io_co(FullAdder_3588_io_co)
  );
  FullAdder FullAdder_3589 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3589_io_a),
    .io_b(FullAdder_3589_io_b),
    .io_ci(FullAdder_3589_io_ci),
    .io_s(FullAdder_3589_io_s),
    .io_co(FullAdder_3589_io_co)
  );
  FullAdder FullAdder_3590 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3590_io_a),
    .io_b(FullAdder_3590_io_b),
    .io_ci(FullAdder_3590_io_ci),
    .io_s(FullAdder_3590_io_s),
    .io_co(FullAdder_3590_io_co)
  );
  FullAdder FullAdder_3591 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3591_io_a),
    .io_b(FullAdder_3591_io_b),
    .io_ci(FullAdder_3591_io_ci),
    .io_s(FullAdder_3591_io_s),
    .io_co(FullAdder_3591_io_co)
  );
  FullAdder FullAdder_3592 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3592_io_a),
    .io_b(FullAdder_3592_io_b),
    .io_ci(FullAdder_3592_io_ci),
    .io_s(FullAdder_3592_io_s),
    .io_co(FullAdder_3592_io_co)
  );
  HalfAdder HalfAdder_171 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_171_io_a),
    .io_b(HalfAdder_171_io_b),
    .io_s(HalfAdder_171_io_s),
    .io_co(HalfAdder_171_io_co)
  );
  FullAdder FullAdder_3593 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3593_io_a),
    .io_b(FullAdder_3593_io_b),
    .io_ci(FullAdder_3593_io_ci),
    .io_s(FullAdder_3593_io_s),
    .io_co(FullAdder_3593_io_co)
  );
  FullAdder FullAdder_3594 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3594_io_a),
    .io_b(FullAdder_3594_io_b),
    .io_ci(FullAdder_3594_io_ci),
    .io_s(FullAdder_3594_io_s),
    .io_co(FullAdder_3594_io_co)
  );
  HalfAdder HalfAdder_172 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_172_io_a),
    .io_b(HalfAdder_172_io_b),
    .io_s(HalfAdder_172_io_s),
    .io_co(HalfAdder_172_io_co)
  );
  FullAdder FullAdder_3595 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3595_io_a),
    .io_b(FullAdder_3595_io_b),
    .io_ci(FullAdder_3595_io_ci),
    .io_s(FullAdder_3595_io_s),
    .io_co(FullAdder_3595_io_co)
  );
  FullAdder FullAdder_3596 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3596_io_a),
    .io_b(FullAdder_3596_io_b),
    .io_ci(FullAdder_3596_io_ci),
    .io_s(FullAdder_3596_io_s),
    .io_co(FullAdder_3596_io_co)
  );
  FullAdder FullAdder_3597 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3597_io_a),
    .io_b(FullAdder_3597_io_b),
    .io_ci(FullAdder_3597_io_ci),
    .io_s(FullAdder_3597_io_s),
    .io_co(FullAdder_3597_io_co)
  );
  FullAdder FullAdder_3598 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3598_io_a),
    .io_b(FullAdder_3598_io_b),
    .io_ci(FullAdder_3598_io_ci),
    .io_s(FullAdder_3598_io_s),
    .io_co(FullAdder_3598_io_co)
  );
  HalfAdder HalfAdder_173 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_173_io_a),
    .io_b(HalfAdder_173_io_b),
    .io_s(HalfAdder_173_io_s),
    .io_co(HalfAdder_173_io_co)
  );
  FullAdder FullAdder_3599 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3599_io_a),
    .io_b(FullAdder_3599_io_b),
    .io_ci(FullAdder_3599_io_ci),
    .io_s(FullAdder_3599_io_s),
    .io_co(FullAdder_3599_io_co)
  );
  HalfAdder HalfAdder_174 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_174_io_a),
    .io_b(HalfAdder_174_io_b),
    .io_s(HalfAdder_174_io_s),
    .io_co(HalfAdder_174_io_co)
  );
  HalfAdder HalfAdder_175 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_175_io_a),
    .io_b(HalfAdder_175_io_b),
    .io_s(HalfAdder_175_io_s),
    .io_co(HalfAdder_175_io_co)
  );
  FullAdder FullAdder_3600 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3600_io_a),
    .io_b(FullAdder_3600_io_b),
    .io_ci(FullAdder_3600_io_ci),
    .io_s(FullAdder_3600_io_s),
    .io_co(FullAdder_3600_io_co)
  );
  HalfAdder HalfAdder_176 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_176_io_a),
    .io_b(HalfAdder_176_io_b),
    .io_s(HalfAdder_176_io_s),
    .io_co(HalfAdder_176_io_co)
  );
  HalfAdder HalfAdder_177 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_177_io_a),
    .io_b(HalfAdder_177_io_b),
    .io_s(HalfAdder_177_io_s),
    .io_co(HalfAdder_177_io_co)
  );
  HalfAdder HalfAdder_178 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_178_io_a),
    .io_b(HalfAdder_178_io_b),
    .io_s(HalfAdder_178_io_s),
    .io_co(HalfAdder_178_io_co)
  );
  FullAdder FullAdder_3601 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3601_io_a),
    .io_b(FullAdder_3601_io_b),
    .io_ci(FullAdder_3601_io_ci),
    .io_s(FullAdder_3601_io_s),
    .io_co(FullAdder_3601_io_co)
  );
  FullAdder FullAdder_3602 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3602_io_a),
    .io_b(FullAdder_3602_io_b),
    .io_ci(FullAdder_3602_io_ci),
    .io_s(FullAdder_3602_io_s),
    .io_co(FullAdder_3602_io_co)
  );
  FullAdder FullAdder_3603 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3603_io_a),
    .io_b(FullAdder_3603_io_b),
    .io_ci(FullAdder_3603_io_ci),
    .io_s(FullAdder_3603_io_s),
    .io_co(FullAdder_3603_io_co)
  );
  FullAdder FullAdder_3604 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3604_io_a),
    .io_b(FullAdder_3604_io_b),
    .io_ci(FullAdder_3604_io_ci),
    .io_s(FullAdder_3604_io_s),
    .io_co(FullAdder_3604_io_co)
  );
  HalfAdder HalfAdder_179 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_179_io_a),
    .io_b(HalfAdder_179_io_b),
    .io_s(HalfAdder_179_io_s),
    .io_co(HalfAdder_179_io_co)
  );
  FullAdder FullAdder_3605 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3605_io_a),
    .io_b(FullAdder_3605_io_b),
    .io_ci(FullAdder_3605_io_ci),
    .io_s(FullAdder_3605_io_s),
    .io_co(FullAdder_3605_io_co)
  );
  FullAdder FullAdder_3606 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3606_io_a),
    .io_b(FullAdder_3606_io_b),
    .io_ci(FullAdder_3606_io_ci),
    .io_s(FullAdder_3606_io_s),
    .io_co(FullAdder_3606_io_co)
  );
  FullAdder FullAdder_3607 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3607_io_a),
    .io_b(FullAdder_3607_io_b),
    .io_ci(FullAdder_3607_io_ci),
    .io_s(FullAdder_3607_io_s),
    .io_co(FullAdder_3607_io_co)
  );
  HalfAdder HalfAdder_180 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_180_io_a),
    .io_b(HalfAdder_180_io_b),
    .io_s(HalfAdder_180_io_s),
    .io_co(HalfAdder_180_io_co)
  );
  FullAdder FullAdder_3608 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3608_io_a),
    .io_b(FullAdder_3608_io_b),
    .io_ci(FullAdder_3608_io_ci),
    .io_s(FullAdder_3608_io_s),
    .io_co(FullAdder_3608_io_co)
  );
  FullAdder FullAdder_3609 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3609_io_a),
    .io_b(FullAdder_3609_io_b),
    .io_ci(FullAdder_3609_io_ci),
    .io_s(FullAdder_3609_io_s),
    .io_co(FullAdder_3609_io_co)
  );
  FullAdder FullAdder_3610 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3610_io_a),
    .io_b(FullAdder_3610_io_b),
    .io_ci(FullAdder_3610_io_ci),
    .io_s(FullAdder_3610_io_s),
    .io_co(FullAdder_3610_io_co)
  );
  FullAdder FullAdder_3611 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3611_io_a),
    .io_b(FullAdder_3611_io_b),
    .io_ci(FullAdder_3611_io_ci),
    .io_s(FullAdder_3611_io_s),
    .io_co(FullAdder_3611_io_co)
  );
  FullAdder FullAdder_3612 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3612_io_a),
    .io_b(FullAdder_3612_io_b),
    .io_ci(FullAdder_3612_io_ci),
    .io_s(FullAdder_3612_io_s),
    .io_co(FullAdder_3612_io_co)
  );
  HalfAdder HalfAdder_181 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_181_io_a),
    .io_b(HalfAdder_181_io_b),
    .io_s(HalfAdder_181_io_s),
    .io_co(HalfAdder_181_io_co)
  );
  FullAdder FullAdder_3613 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3613_io_a),
    .io_b(FullAdder_3613_io_b),
    .io_ci(FullAdder_3613_io_ci),
    .io_s(FullAdder_3613_io_s),
    .io_co(FullAdder_3613_io_co)
  );
  FullAdder FullAdder_3614 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3614_io_a),
    .io_b(FullAdder_3614_io_b),
    .io_ci(FullAdder_3614_io_ci),
    .io_s(FullAdder_3614_io_s),
    .io_co(FullAdder_3614_io_co)
  );
  FullAdder FullAdder_3615 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3615_io_a),
    .io_b(FullAdder_3615_io_b),
    .io_ci(FullAdder_3615_io_ci),
    .io_s(FullAdder_3615_io_s),
    .io_co(FullAdder_3615_io_co)
  );
  FullAdder FullAdder_3616 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3616_io_a),
    .io_b(FullAdder_3616_io_b),
    .io_ci(FullAdder_3616_io_ci),
    .io_s(FullAdder_3616_io_s),
    .io_co(FullAdder_3616_io_co)
  );
  FullAdder FullAdder_3617 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3617_io_a),
    .io_b(FullAdder_3617_io_b),
    .io_ci(FullAdder_3617_io_ci),
    .io_s(FullAdder_3617_io_s),
    .io_co(FullAdder_3617_io_co)
  );
  FullAdder FullAdder_3618 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3618_io_a),
    .io_b(FullAdder_3618_io_b),
    .io_ci(FullAdder_3618_io_ci),
    .io_s(FullAdder_3618_io_s),
    .io_co(FullAdder_3618_io_co)
  );
  HalfAdder HalfAdder_182 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_182_io_a),
    .io_b(HalfAdder_182_io_b),
    .io_s(HalfAdder_182_io_s),
    .io_co(HalfAdder_182_io_co)
  );
  HalfAdder HalfAdder_183 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_183_io_a),
    .io_b(HalfAdder_183_io_b),
    .io_s(HalfAdder_183_io_s),
    .io_co(HalfAdder_183_io_co)
  );
  FullAdder FullAdder_3619 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3619_io_a),
    .io_b(FullAdder_3619_io_b),
    .io_ci(FullAdder_3619_io_ci),
    .io_s(FullAdder_3619_io_s),
    .io_co(FullAdder_3619_io_co)
  );
  FullAdder FullAdder_3620 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3620_io_a),
    .io_b(FullAdder_3620_io_b),
    .io_ci(FullAdder_3620_io_ci),
    .io_s(FullAdder_3620_io_s),
    .io_co(FullAdder_3620_io_co)
  );
  FullAdder FullAdder_3621 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3621_io_a),
    .io_b(FullAdder_3621_io_b),
    .io_ci(FullAdder_3621_io_ci),
    .io_s(FullAdder_3621_io_s),
    .io_co(FullAdder_3621_io_co)
  );
  FullAdder FullAdder_3622 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3622_io_a),
    .io_b(FullAdder_3622_io_b),
    .io_ci(FullAdder_3622_io_ci),
    .io_s(FullAdder_3622_io_s),
    .io_co(FullAdder_3622_io_co)
  );
  HalfAdder HalfAdder_184 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_184_io_a),
    .io_b(HalfAdder_184_io_b),
    .io_s(HalfAdder_184_io_s),
    .io_co(HalfAdder_184_io_co)
  );
  HalfAdder HalfAdder_185 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_185_io_a),
    .io_b(HalfAdder_185_io_b),
    .io_s(HalfAdder_185_io_s),
    .io_co(HalfAdder_185_io_co)
  );
  HalfAdder HalfAdder_186 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_186_io_a),
    .io_b(HalfAdder_186_io_b),
    .io_s(HalfAdder_186_io_s),
    .io_co(HalfAdder_186_io_co)
  );
  FullAdder FullAdder_3623 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3623_io_a),
    .io_b(FullAdder_3623_io_b),
    .io_ci(FullAdder_3623_io_ci),
    .io_s(FullAdder_3623_io_s),
    .io_co(FullAdder_3623_io_co)
  );
  FullAdder FullAdder_3624 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3624_io_a),
    .io_b(FullAdder_3624_io_b),
    .io_ci(FullAdder_3624_io_ci),
    .io_s(FullAdder_3624_io_s),
    .io_co(FullAdder_3624_io_co)
  );
  HalfAdder HalfAdder_187 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_187_io_a),
    .io_b(HalfAdder_187_io_b),
    .io_s(HalfAdder_187_io_s),
    .io_co(HalfAdder_187_io_co)
  );
  FullAdder FullAdder_3625 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3625_io_a),
    .io_b(FullAdder_3625_io_b),
    .io_ci(FullAdder_3625_io_ci),
    .io_s(FullAdder_3625_io_s),
    .io_co(FullAdder_3625_io_co)
  );
  FullAdder FullAdder_3626 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3626_io_a),
    .io_b(FullAdder_3626_io_b),
    .io_ci(FullAdder_3626_io_ci),
    .io_s(FullAdder_3626_io_s),
    .io_co(FullAdder_3626_io_co)
  );
  HalfAdder HalfAdder_188 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_188_io_a),
    .io_b(HalfAdder_188_io_b),
    .io_s(HalfAdder_188_io_s),
    .io_co(HalfAdder_188_io_co)
  );
  HalfAdder HalfAdder_189 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_189_io_a),
    .io_b(HalfAdder_189_io_b),
    .io_s(HalfAdder_189_io_s),
    .io_co(HalfAdder_189_io_co)
  );
  FullAdder FullAdder_3627 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3627_io_a),
    .io_b(FullAdder_3627_io_b),
    .io_ci(FullAdder_3627_io_ci),
    .io_s(FullAdder_3627_io_s),
    .io_co(FullAdder_3627_io_co)
  );
  FullAdder FullAdder_3628 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3628_io_a),
    .io_b(FullAdder_3628_io_b),
    .io_ci(FullAdder_3628_io_ci),
    .io_s(FullAdder_3628_io_s),
    .io_co(FullAdder_3628_io_co)
  );
  FullAdder FullAdder_3629 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3629_io_a),
    .io_b(FullAdder_3629_io_b),
    .io_ci(FullAdder_3629_io_ci),
    .io_s(FullAdder_3629_io_s),
    .io_co(FullAdder_3629_io_co)
  );
  FullAdder FullAdder_3630 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3630_io_a),
    .io_b(FullAdder_3630_io_b),
    .io_ci(FullAdder_3630_io_ci),
    .io_s(FullAdder_3630_io_s),
    .io_co(FullAdder_3630_io_co)
  );
  FullAdder FullAdder_3631 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3631_io_a),
    .io_b(FullAdder_3631_io_b),
    .io_ci(FullAdder_3631_io_ci),
    .io_s(FullAdder_3631_io_s),
    .io_co(FullAdder_3631_io_co)
  );
  HalfAdder HalfAdder_190 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_190_io_a),
    .io_b(HalfAdder_190_io_b),
    .io_s(HalfAdder_190_io_s),
    .io_co(HalfAdder_190_io_co)
  );
  FullAdder FullAdder_3632 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3632_io_a),
    .io_b(FullAdder_3632_io_b),
    .io_ci(FullAdder_3632_io_ci),
    .io_s(FullAdder_3632_io_s),
    .io_co(FullAdder_3632_io_co)
  );
  FullAdder FullAdder_3633 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3633_io_a),
    .io_b(FullAdder_3633_io_b),
    .io_ci(FullAdder_3633_io_ci),
    .io_s(FullAdder_3633_io_s),
    .io_co(FullAdder_3633_io_co)
  );
  FullAdder FullAdder_3634 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3634_io_a),
    .io_b(FullAdder_3634_io_b),
    .io_ci(FullAdder_3634_io_ci),
    .io_s(FullAdder_3634_io_s),
    .io_co(FullAdder_3634_io_co)
  );
  FullAdder FullAdder_3635 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3635_io_a),
    .io_b(FullAdder_3635_io_b),
    .io_ci(FullAdder_3635_io_ci),
    .io_s(FullAdder_3635_io_s),
    .io_co(FullAdder_3635_io_co)
  );
  FullAdder FullAdder_3636 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3636_io_a),
    .io_b(FullAdder_3636_io_b),
    .io_ci(FullAdder_3636_io_ci),
    .io_s(FullAdder_3636_io_s),
    .io_co(FullAdder_3636_io_co)
  );
  FullAdder FullAdder_3637 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3637_io_a),
    .io_b(FullAdder_3637_io_b),
    .io_ci(FullAdder_3637_io_ci),
    .io_s(FullAdder_3637_io_s),
    .io_co(FullAdder_3637_io_co)
  );
  FullAdder FullAdder_3638 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3638_io_a),
    .io_b(FullAdder_3638_io_b),
    .io_ci(FullAdder_3638_io_ci),
    .io_s(FullAdder_3638_io_s),
    .io_co(FullAdder_3638_io_co)
  );
  FullAdder FullAdder_3639 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3639_io_a),
    .io_b(FullAdder_3639_io_b),
    .io_ci(FullAdder_3639_io_ci),
    .io_s(FullAdder_3639_io_s),
    .io_co(FullAdder_3639_io_co)
  );
  FullAdder FullAdder_3640 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3640_io_a),
    .io_b(FullAdder_3640_io_b),
    .io_ci(FullAdder_3640_io_ci),
    .io_s(FullAdder_3640_io_s),
    .io_co(FullAdder_3640_io_co)
  );
  FullAdder FullAdder_3641 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3641_io_a),
    .io_b(FullAdder_3641_io_b),
    .io_ci(FullAdder_3641_io_ci),
    .io_s(FullAdder_3641_io_s),
    .io_co(FullAdder_3641_io_co)
  );
  HalfAdder HalfAdder_191 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_191_io_a),
    .io_b(HalfAdder_191_io_b),
    .io_s(HalfAdder_191_io_s),
    .io_co(HalfAdder_191_io_co)
  );
  FullAdder FullAdder_3642 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3642_io_a),
    .io_b(FullAdder_3642_io_b),
    .io_ci(FullAdder_3642_io_ci),
    .io_s(FullAdder_3642_io_s),
    .io_co(FullAdder_3642_io_co)
  );
  FullAdder FullAdder_3643 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3643_io_a),
    .io_b(FullAdder_3643_io_b),
    .io_ci(FullAdder_3643_io_ci),
    .io_s(FullAdder_3643_io_s),
    .io_co(FullAdder_3643_io_co)
  );
  FullAdder FullAdder_3644 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3644_io_a),
    .io_b(FullAdder_3644_io_b),
    .io_ci(FullAdder_3644_io_ci),
    .io_s(FullAdder_3644_io_s),
    .io_co(FullAdder_3644_io_co)
  );
  FullAdder FullAdder_3645 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3645_io_a),
    .io_b(FullAdder_3645_io_b),
    .io_ci(FullAdder_3645_io_ci),
    .io_s(FullAdder_3645_io_s),
    .io_co(FullAdder_3645_io_co)
  );
  FullAdder FullAdder_3646 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3646_io_a),
    .io_b(FullAdder_3646_io_b),
    .io_ci(FullAdder_3646_io_ci),
    .io_s(FullAdder_3646_io_s),
    .io_co(FullAdder_3646_io_co)
  );
  FullAdder FullAdder_3647 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3647_io_a),
    .io_b(FullAdder_3647_io_b),
    .io_ci(FullAdder_3647_io_ci),
    .io_s(FullAdder_3647_io_s),
    .io_co(FullAdder_3647_io_co)
  );
  FullAdder FullAdder_3648 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3648_io_a),
    .io_b(FullAdder_3648_io_b),
    .io_ci(FullAdder_3648_io_ci),
    .io_s(FullAdder_3648_io_s),
    .io_co(FullAdder_3648_io_co)
  );
  FullAdder FullAdder_3649 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3649_io_a),
    .io_b(FullAdder_3649_io_b),
    .io_ci(FullAdder_3649_io_ci),
    .io_s(FullAdder_3649_io_s),
    .io_co(FullAdder_3649_io_co)
  );
  FullAdder FullAdder_3650 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3650_io_a),
    .io_b(FullAdder_3650_io_b),
    .io_ci(FullAdder_3650_io_ci),
    .io_s(FullAdder_3650_io_s),
    .io_co(FullAdder_3650_io_co)
  );
  FullAdder FullAdder_3651 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3651_io_a),
    .io_b(FullAdder_3651_io_b),
    .io_ci(FullAdder_3651_io_ci),
    .io_s(FullAdder_3651_io_s),
    .io_co(FullAdder_3651_io_co)
  );
  HalfAdder HalfAdder_192 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_192_io_a),
    .io_b(HalfAdder_192_io_b),
    .io_s(HalfAdder_192_io_s),
    .io_co(HalfAdder_192_io_co)
  );
  HalfAdder HalfAdder_193 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_193_io_a),
    .io_b(HalfAdder_193_io_b),
    .io_s(HalfAdder_193_io_s),
    .io_co(HalfAdder_193_io_co)
  );
  HalfAdder HalfAdder_194 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_194_io_a),
    .io_b(HalfAdder_194_io_b),
    .io_s(HalfAdder_194_io_s),
    .io_co(HalfAdder_194_io_co)
  );
  FullAdder FullAdder_3652 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3652_io_a),
    .io_b(FullAdder_3652_io_b),
    .io_ci(FullAdder_3652_io_ci),
    .io_s(FullAdder_3652_io_s),
    .io_co(FullAdder_3652_io_co)
  );
  FullAdder FullAdder_3653 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3653_io_a),
    .io_b(FullAdder_3653_io_b),
    .io_ci(FullAdder_3653_io_ci),
    .io_s(FullAdder_3653_io_s),
    .io_co(FullAdder_3653_io_co)
  );
  FullAdder FullAdder_3654 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3654_io_a),
    .io_b(FullAdder_3654_io_b),
    .io_ci(FullAdder_3654_io_ci),
    .io_s(FullAdder_3654_io_s),
    .io_co(FullAdder_3654_io_co)
  );
  FullAdder FullAdder_3655 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3655_io_a),
    .io_b(FullAdder_3655_io_b),
    .io_ci(FullAdder_3655_io_ci),
    .io_s(FullAdder_3655_io_s),
    .io_co(FullAdder_3655_io_co)
  );
  FullAdder FullAdder_3656 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3656_io_a),
    .io_b(FullAdder_3656_io_b),
    .io_ci(FullAdder_3656_io_ci),
    .io_s(FullAdder_3656_io_s),
    .io_co(FullAdder_3656_io_co)
  );
  FullAdder FullAdder_3657 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3657_io_a),
    .io_b(FullAdder_3657_io_b),
    .io_ci(FullAdder_3657_io_ci),
    .io_s(FullAdder_3657_io_s),
    .io_co(FullAdder_3657_io_co)
  );
  FullAdder FullAdder_3658 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3658_io_a),
    .io_b(FullAdder_3658_io_b),
    .io_ci(FullAdder_3658_io_ci),
    .io_s(FullAdder_3658_io_s),
    .io_co(FullAdder_3658_io_co)
  );
  FullAdder FullAdder_3659 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3659_io_a),
    .io_b(FullAdder_3659_io_b),
    .io_ci(FullAdder_3659_io_ci),
    .io_s(FullAdder_3659_io_s),
    .io_co(FullAdder_3659_io_co)
  );
  FullAdder FullAdder_3660 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3660_io_a),
    .io_b(FullAdder_3660_io_b),
    .io_ci(FullAdder_3660_io_ci),
    .io_s(FullAdder_3660_io_s),
    .io_co(FullAdder_3660_io_co)
  );
  HalfAdder HalfAdder_195 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_195_io_a),
    .io_b(HalfAdder_195_io_b),
    .io_s(HalfAdder_195_io_s),
    .io_co(HalfAdder_195_io_co)
  );
  FullAdder FullAdder_3661 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3661_io_a),
    .io_b(FullAdder_3661_io_b),
    .io_ci(FullAdder_3661_io_ci),
    .io_s(FullAdder_3661_io_s),
    .io_co(FullAdder_3661_io_co)
  );
  FullAdder FullAdder_3662 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3662_io_a),
    .io_b(FullAdder_3662_io_b),
    .io_ci(FullAdder_3662_io_ci),
    .io_s(FullAdder_3662_io_s),
    .io_co(FullAdder_3662_io_co)
  );
  FullAdder FullAdder_3663 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3663_io_a),
    .io_b(FullAdder_3663_io_b),
    .io_ci(FullAdder_3663_io_ci),
    .io_s(FullAdder_3663_io_s),
    .io_co(FullAdder_3663_io_co)
  );
  FullAdder FullAdder_3664 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3664_io_a),
    .io_b(FullAdder_3664_io_b),
    .io_ci(FullAdder_3664_io_ci),
    .io_s(FullAdder_3664_io_s),
    .io_co(FullAdder_3664_io_co)
  );
  FullAdder FullAdder_3665 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3665_io_a),
    .io_b(FullAdder_3665_io_b),
    .io_ci(FullAdder_3665_io_ci),
    .io_s(FullAdder_3665_io_s),
    .io_co(FullAdder_3665_io_co)
  );
  FullAdder FullAdder_3666 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3666_io_a),
    .io_b(FullAdder_3666_io_b),
    .io_ci(FullAdder_3666_io_ci),
    .io_s(FullAdder_3666_io_s),
    .io_co(FullAdder_3666_io_co)
  );
  FullAdder FullAdder_3667 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3667_io_a),
    .io_b(FullAdder_3667_io_b),
    .io_ci(FullAdder_3667_io_ci),
    .io_s(FullAdder_3667_io_s),
    .io_co(FullAdder_3667_io_co)
  );
  FullAdder FullAdder_3668 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3668_io_a),
    .io_b(FullAdder_3668_io_b),
    .io_ci(FullAdder_3668_io_ci),
    .io_s(FullAdder_3668_io_s),
    .io_co(FullAdder_3668_io_co)
  );
  FullAdder FullAdder_3669 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3669_io_a),
    .io_b(FullAdder_3669_io_b),
    .io_ci(FullAdder_3669_io_ci),
    .io_s(FullAdder_3669_io_s),
    .io_co(FullAdder_3669_io_co)
  );
  FullAdder FullAdder_3670 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3670_io_a),
    .io_b(FullAdder_3670_io_b),
    .io_ci(FullAdder_3670_io_ci),
    .io_s(FullAdder_3670_io_s),
    .io_co(FullAdder_3670_io_co)
  );
  FullAdder FullAdder_3671 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3671_io_a),
    .io_b(FullAdder_3671_io_b),
    .io_ci(FullAdder_3671_io_ci),
    .io_s(FullAdder_3671_io_s),
    .io_co(FullAdder_3671_io_co)
  );
  FullAdder FullAdder_3672 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3672_io_a),
    .io_b(FullAdder_3672_io_b),
    .io_ci(FullAdder_3672_io_ci),
    .io_s(FullAdder_3672_io_s),
    .io_co(FullAdder_3672_io_co)
  );
  FullAdder FullAdder_3673 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3673_io_a),
    .io_b(FullAdder_3673_io_b),
    .io_ci(FullAdder_3673_io_ci),
    .io_s(FullAdder_3673_io_s),
    .io_co(FullAdder_3673_io_co)
  );
  FullAdder FullAdder_3674 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3674_io_a),
    .io_b(FullAdder_3674_io_b),
    .io_ci(FullAdder_3674_io_ci),
    .io_s(FullAdder_3674_io_s),
    .io_co(FullAdder_3674_io_co)
  );
  FullAdder FullAdder_3675 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3675_io_a),
    .io_b(FullAdder_3675_io_b),
    .io_ci(FullAdder_3675_io_ci),
    .io_s(FullAdder_3675_io_s),
    .io_co(FullAdder_3675_io_co)
  );
  FullAdder FullAdder_3676 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3676_io_a),
    .io_b(FullAdder_3676_io_b),
    .io_ci(FullAdder_3676_io_ci),
    .io_s(FullAdder_3676_io_s),
    .io_co(FullAdder_3676_io_co)
  );
  FullAdder FullAdder_3677 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3677_io_a),
    .io_b(FullAdder_3677_io_b),
    .io_ci(FullAdder_3677_io_ci),
    .io_s(FullAdder_3677_io_s),
    .io_co(FullAdder_3677_io_co)
  );
  FullAdder FullAdder_3678 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3678_io_a),
    .io_b(FullAdder_3678_io_b),
    .io_ci(FullAdder_3678_io_ci),
    .io_s(FullAdder_3678_io_s),
    .io_co(FullAdder_3678_io_co)
  );
  HalfAdder HalfAdder_196 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_196_io_a),
    .io_b(HalfAdder_196_io_b),
    .io_s(HalfAdder_196_io_s),
    .io_co(HalfAdder_196_io_co)
  );
  FullAdder FullAdder_3679 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3679_io_a),
    .io_b(FullAdder_3679_io_b),
    .io_ci(FullAdder_3679_io_ci),
    .io_s(FullAdder_3679_io_s),
    .io_co(FullAdder_3679_io_co)
  );
  FullAdder FullAdder_3680 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3680_io_a),
    .io_b(FullAdder_3680_io_b),
    .io_ci(FullAdder_3680_io_ci),
    .io_s(FullAdder_3680_io_s),
    .io_co(FullAdder_3680_io_co)
  );
  FullAdder FullAdder_3681 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3681_io_a),
    .io_b(FullAdder_3681_io_b),
    .io_ci(FullAdder_3681_io_ci),
    .io_s(FullAdder_3681_io_s),
    .io_co(FullAdder_3681_io_co)
  );
  FullAdder FullAdder_3682 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3682_io_a),
    .io_b(FullAdder_3682_io_b),
    .io_ci(FullAdder_3682_io_ci),
    .io_s(FullAdder_3682_io_s),
    .io_co(FullAdder_3682_io_co)
  );
  HalfAdder HalfAdder_197 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_197_io_a),
    .io_b(HalfAdder_197_io_b),
    .io_s(HalfAdder_197_io_s),
    .io_co(HalfAdder_197_io_co)
  );
  FullAdder FullAdder_3683 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3683_io_a),
    .io_b(FullAdder_3683_io_b),
    .io_ci(FullAdder_3683_io_ci),
    .io_s(FullAdder_3683_io_s),
    .io_co(FullAdder_3683_io_co)
  );
  FullAdder FullAdder_3684 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3684_io_a),
    .io_b(FullAdder_3684_io_b),
    .io_ci(FullAdder_3684_io_ci),
    .io_s(FullAdder_3684_io_s),
    .io_co(FullAdder_3684_io_co)
  );
  FullAdder FullAdder_3685 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3685_io_a),
    .io_b(FullAdder_3685_io_b),
    .io_ci(FullAdder_3685_io_ci),
    .io_s(FullAdder_3685_io_s),
    .io_co(FullAdder_3685_io_co)
  );
  FullAdder FullAdder_3686 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3686_io_a),
    .io_b(FullAdder_3686_io_b),
    .io_ci(FullAdder_3686_io_ci),
    .io_s(FullAdder_3686_io_s),
    .io_co(FullAdder_3686_io_co)
  );
  FullAdder FullAdder_3687 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3687_io_a),
    .io_b(FullAdder_3687_io_b),
    .io_ci(FullAdder_3687_io_ci),
    .io_s(FullAdder_3687_io_s),
    .io_co(FullAdder_3687_io_co)
  );
  FullAdder FullAdder_3688 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3688_io_a),
    .io_b(FullAdder_3688_io_b),
    .io_ci(FullAdder_3688_io_ci),
    .io_s(FullAdder_3688_io_s),
    .io_co(FullAdder_3688_io_co)
  );
  FullAdder FullAdder_3689 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3689_io_a),
    .io_b(FullAdder_3689_io_b),
    .io_ci(FullAdder_3689_io_ci),
    .io_s(FullAdder_3689_io_s),
    .io_co(FullAdder_3689_io_co)
  );
  FullAdder FullAdder_3690 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3690_io_a),
    .io_b(FullAdder_3690_io_b),
    .io_ci(FullAdder_3690_io_ci),
    .io_s(FullAdder_3690_io_s),
    .io_co(FullAdder_3690_io_co)
  );
  FullAdder FullAdder_3691 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3691_io_a),
    .io_b(FullAdder_3691_io_b),
    .io_ci(FullAdder_3691_io_ci),
    .io_s(FullAdder_3691_io_s),
    .io_co(FullAdder_3691_io_co)
  );
  FullAdder FullAdder_3692 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3692_io_a),
    .io_b(FullAdder_3692_io_b),
    .io_ci(FullAdder_3692_io_ci),
    .io_s(FullAdder_3692_io_s),
    .io_co(FullAdder_3692_io_co)
  );
  FullAdder FullAdder_3693 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3693_io_a),
    .io_b(FullAdder_3693_io_b),
    .io_ci(FullAdder_3693_io_ci),
    .io_s(FullAdder_3693_io_s),
    .io_co(FullAdder_3693_io_co)
  );
  FullAdder FullAdder_3694 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3694_io_a),
    .io_b(FullAdder_3694_io_b),
    .io_ci(FullAdder_3694_io_ci),
    .io_s(FullAdder_3694_io_s),
    .io_co(FullAdder_3694_io_co)
  );
  FullAdder FullAdder_3695 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3695_io_a),
    .io_b(FullAdder_3695_io_b),
    .io_ci(FullAdder_3695_io_ci),
    .io_s(FullAdder_3695_io_s),
    .io_co(FullAdder_3695_io_co)
  );
  FullAdder FullAdder_3696 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3696_io_a),
    .io_b(FullAdder_3696_io_b),
    .io_ci(FullAdder_3696_io_ci),
    .io_s(FullAdder_3696_io_s),
    .io_co(FullAdder_3696_io_co)
  );
  FullAdder FullAdder_3697 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3697_io_a),
    .io_b(FullAdder_3697_io_b),
    .io_ci(FullAdder_3697_io_ci),
    .io_s(FullAdder_3697_io_s),
    .io_co(FullAdder_3697_io_co)
  );
  FullAdder FullAdder_3698 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3698_io_a),
    .io_b(FullAdder_3698_io_b),
    .io_ci(FullAdder_3698_io_ci),
    .io_s(FullAdder_3698_io_s),
    .io_co(FullAdder_3698_io_co)
  );
  FullAdder FullAdder_3699 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3699_io_a),
    .io_b(FullAdder_3699_io_b),
    .io_ci(FullAdder_3699_io_ci),
    .io_s(FullAdder_3699_io_s),
    .io_co(FullAdder_3699_io_co)
  );
  FullAdder FullAdder_3700 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3700_io_a),
    .io_b(FullAdder_3700_io_b),
    .io_ci(FullAdder_3700_io_ci),
    .io_s(FullAdder_3700_io_s),
    .io_co(FullAdder_3700_io_co)
  );
  FullAdder FullAdder_3701 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3701_io_a),
    .io_b(FullAdder_3701_io_b),
    .io_ci(FullAdder_3701_io_ci),
    .io_s(FullAdder_3701_io_s),
    .io_co(FullAdder_3701_io_co)
  );
  FullAdder FullAdder_3702 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3702_io_a),
    .io_b(FullAdder_3702_io_b),
    .io_ci(FullAdder_3702_io_ci),
    .io_s(FullAdder_3702_io_s),
    .io_co(FullAdder_3702_io_co)
  );
  HalfAdder HalfAdder_198 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_198_io_a),
    .io_b(HalfAdder_198_io_b),
    .io_s(HalfAdder_198_io_s),
    .io_co(HalfAdder_198_io_co)
  );
  FullAdder FullAdder_3703 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3703_io_a),
    .io_b(FullAdder_3703_io_b),
    .io_ci(FullAdder_3703_io_ci),
    .io_s(FullAdder_3703_io_s),
    .io_co(FullAdder_3703_io_co)
  );
  FullAdder FullAdder_3704 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3704_io_a),
    .io_b(FullAdder_3704_io_b),
    .io_ci(FullAdder_3704_io_ci),
    .io_s(FullAdder_3704_io_s),
    .io_co(FullAdder_3704_io_co)
  );
  FullAdder FullAdder_3705 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3705_io_a),
    .io_b(FullAdder_3705_io_b),
    .io_ci(FullAdder_3705_io_ci),
    .io_s(FullAdder_3705_io_s),
    .io_co(FullAdder_3705_io_co)
  );
  FullAdder FullAdder_3706 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3706_io_a),
    .io_b(FullAdder_3706_io_b),
    .io_ci(FullAdder_3706_io_ci),
    .io_s(FullAdder_3706_io_s),
    .io_co(FullAdder_3706_io_co)
  );
  HalfAdder HalfAdder_199 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_199_io_a),
    .io_b(HalfAdder_199_io_b),
    .io_s(HalfAdder_199_io_s),
    .io_co(HalfAdder_199_io_co)
  );
  HalfAdder HalfAdder_200 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_200_io_a),
    .io_b(HalfAdder_200_io_b),
    .io_s(HalfAdder_200_io_s),
    .io_co(HalfAdder_200_io_co)
  );
  FullAdder FullAdder_3707 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3707_io_a),
    .io_b(FullAdder_3707_io_b),
    .io_ci(FullAdder_3707_io_ci),
    .io_s(FullAdder_3707_io_s),
    .io_co(FullAdder_3707_io_co)
  );
  FullAdder FullAdder_3708 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3708_io_a),
    .io_b(FullAdder_3708_io_b),
    .io_ci(FullAdder_3708_io_ci),
    .io_s(FullAdder_3708_io_s),
    .io_co(FullAdder_3708_io_co)
  );
  FullAdder FullAdder_3709 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3709_io_a),
    .io_b(FullAdder_3709_io_b),
    .io_ci(FullAdder_3709_io_ci),
    .io_s(FullAdder_3709_io_s),
    .io_co(FullAdder_3709_io_co)
  );
  HalfAdder HalfAdder_201 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_201_io_a),
    .io_b(HalfAdder_201_io_b),
    .io_s(HalfAdder_201_io_s),
    .io_co(HalfAdder_201_io_co)
  );
  FullAdder FullAdder_3710 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3710_io_a),
    .io_b(FullAdder_3710_io_b),
    .io_ci(FullAdder_3710_io_ci),
    .io_s(FullAdder_3710_io_s),
    .io_co(FullAdder_3710_io_co)
  );
  HalfAdder HalfAdder_202 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_202_io_a),
    .io_b(HalfAdder_202_io_b),
    .io_s(HalfAdder_202_io_s),
    .io_co(HalfAdder_202_io_co)
  );
  HalfAdder HalfAdder_203 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_203_io_a),
    .io_b(HalfAdder_203_io_b),
    .io_s(HalfAdder_203_io_s),
    .io_co(HalfAdder_203_io_co)
  );
  FullAdder FullAdder_3711 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3711_io_a),
    .io_b(FullAdder_3711_io_b),
    .io_ci(FullAdder_3711_io_ci),
    .io_s(FullAdder_3711_io_s),
    .io_co(FullAdder_3711_io_co)
  );
  HalfAdder HalfAdder_204 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_204_io_a),
    .io_b(HalfAdder_204_io_b),
    .io_s(HalfAdder_204_io_s),
    .io_co(HalfAdder_204_io_co)
  );
  HalfAdder HalfAdder_205 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_205_io_a),
    .io_b(HalfAdder_205_io_b),
    .io_s(HalfAdder_205_io_s),
    .io_co(HalfAdder_205_io_co)
  );
  FullAdder FullAdder_3712 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3712_io_a),
    .io_b(FullAdder_3712_io_b),
    .io_ci(FullAdder_3712_io_ci),
    .io_s(FullAdder_3712_io_s),
    .io_co(FullAdder_3712_io_co)
  );
  HalfAdder HalfAdder_206 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_206_io_a),
    .io_b(HalfAdder_206_io_b),
    .io_s(HalfAdder_206_io_s),
    .io_co(HalfAdder_206_io_co)
  );
  HalfAdder HalfAdder_207 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_207_io_a),
    .io_b(HalfAdder_207_io_b),
    .io_s(HalfAdder_207_io_s),
    .io_co(HalfAdder_207_io_co)
  );
  HalfAdder HalfAdder_208 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_208_io_a),
    .io_b(HalfAdder_208_io_b),
    .io_s(HalfAdder_208_io_s),
    .io_co(HalfAdder_208_io_co)
  );
  FullAdder FullAdder_3713 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3713_io_a),
    .io_b(FullAdder_3713_io_b),
    .io_ci(FullAdder_3713_io_ci),
    .io_s(FullAdder_3713_io_s),
    .io_co(FullAdder_3713_io_co)
  );
  HalfAdder HalfAdder_209 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_209_io_a),
    .io_b(HalfAdder_209_io_b),
    .io_s(HalfAdder_209_io_s),
    .io_co(HalfAdder_209_io_co)
  );
  FullAdder FullAdder_3714 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3714_io_a),
    .io_b(FullAdder_3714_io_b),
    .io_ci(FullAdder_3714_io_ci),
    .io_s(FullAdder_3714_io_s),
    .io_co(FullAdder_3714_io_co)
  );
  HalfAdder HalfAdder_210 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_210_io_a),
    .io_b(HalfAdder_210_io_b),
    .io_s(HalfAdder_210_io_s),
    .io_co(HalfAdder_210_io_co)
  );
  FullAdder FullAdder_3715 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3715_io_a),
    .io_b(FullAdder_3715_io_b),
    .io_ci(FullAdder_3715_io_ci),
    .io_s(FullAdder_3715_io_s),
    .io_co(FullAdder_3715_io_co)
  );
  FullAdder FullAdder_3716 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3716_io_a),
    .io_b(FullAdder_3716_io_b),
    .io_ci(FullAdder_3716_io_ci),
    .io_s(FullAdder_3716_io_s),
    .io_co(FullAdder_3716_io_co)
  );
  FullAdder FullAdder_3717 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3717_io_a),
    .io_b(FullAdder_3717_io_b),
    .io_ci(FullAdder_3717_io_ci),
    .io_s(FullAdder_3717_io_s),
    .io_co(FullAdder_3717_io_co)
  );
  FullAdder FullAdder_3718 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3718_io_a),
    .io_b(FullAdder_3718_io_b),
    .io_ci(FullAdder_3718_io_ci),
    .io_s(FullAdder_3718_io_s),
    .io_co(FullAdder_3718_io_co)
  );
  FullAdder FullAdder_3719 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3719_io_a),
    .io_b(FullAdder_3719_io_b),
    .io_ci(FullAdder_3719_io_ci),
    .io_s(FullAdder_3719_io_s),
    .io_co(FullAdder_3719_io_co)
  );
  FullAdder FullAdder_3720 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3720_io_a),
    .io_b(FullAdder_3720_io_b),
    .io_ci(FullAdder_3720_io_ci),
    .io_s(FullAdder_3720_io_s),
    .io_co(FullAdder_3720_io_co)
  );
  HalfAdder HalfAdder_211 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_211_io_a),
    .io_b(HalfAdder_211_io_b),
    .io_s(HalfAdder_211_io_s),
    .io_co(HalfAdder_211_io_co)
  );
  HalfAdder HalfAdder_212 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_212_io_a),
    .io_b(HalfAdder_212_io_b),
    .io_s(HalfAdder_212_io_s),
    .io_co(HalfAdder_212_io_co)
  );
  HalfAdder HalfAdder_213 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_213_io_a),
    .io_b(HalfAdder_213_io_b),
    .io_s(HalfAdder_213_io_s),
    .io_co(HalfAdder_213_io_co)
  );
  FullAdder FullAdder_3721 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3721_io_a),
    .io_b(FullAdder_3721_io_b),
    .io_ci(FullAdder_3721_io_ci),
    .io_s(FullAdder_3721_io_s),
    .io_co(FullAdder_3721_io_co)
  );
  FullAdder FullAdder_3722 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3722_io_a),
    .io_b(FullAdder_3722_io_b),
    .io_ci(FullAdder_3722_io_ci),
    .io_s(FullAdder_3722_io_s),
    .io_co(FullAdder_3722_io_co)
  );
  FullAdder FullAdder_3723 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3723_io_a),
    .io_b(FullAdder_3723_io_b),
    .io_ci(FullAdder_3723_io_ci),
    .io_s(FullAdder_3723_io_s),
    .io_co(FullAdder_3723_io_co)
  );
  HalfAdder HalfAdder_214 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_214_io_a),
    .io_b(HalfAdder_214_io_b),
    .io_s(HalfAdder_214_io_s),
    .io_co(HalfAdder_214_io_co)
  );
  HalfAdder HalfAdder_215 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_215_io_a),
    .io_b(HalfAdder_215_io_b),
    .io_s(HalfAdder_215_io_s),
    .io_co(HalfAdder_215_io_co)
  );
  FullAdder FullAdder_3724 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3724_io_a),
    .io_b(FullAdder_3724_io_b),
    .io_ci(FullAdder_3724_io_ci),
    .io_s(FullAdder_3724_io_s),
    .io_co(FullAdder_3724_io_co)
  );
  FullAdder FullAdder_3725 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3725_io_a),
    .io_b(FullAdder_3725_io_b),
    .io_ci(FullAdder_3725_io_ci),
    .io_s(FullAdder_3725_io_s),
    .io_co(FullAdder_3725_io_co)
  );
  FullAdder FullAdder_3726 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3726_io_a),
    .io_b(FullAdder_3726_io_b),
    .io_ci(FullAdder_3726_io_ci),
    .io_s(FullAdder_3726_io_s),
    .io_co(FullAdder_3726_io_co)
  );
  FullAdder FullAdder_3727 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3727_io_a),
    .io_b(FullAdder_3727_io_b),
    .io_ci(FullAdder_3727_io_ci),
    .io_s(FullAdder_3727_io_s),
    .io_co(FullAdder_3727_io_co)
  );
  HalfAdder HalfAdder_216 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_216_io_a),
    .io_b(HalfAdder_216_io_b),
    .io_s(HalfAdder_216_io_s),
    .io_co(HalfAdder_216_io_co)
  );
  HalfAdder HalfAdder_217 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_217_io_a),
    .io_b(HalfAdder_217_io_b),
    .io_s(HalfAdder_217_io_s),
    .io_co(HalfAdder_217_io_co)
  );
  FullAdder FullAdder_3728 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3728_io_a),
    .io_b(FullAdder_3728_io_b),
    .io_ci(FullAdder_3728_io_ci),
    .io_s(FullAdder_3728_io_s),
    .io_co(FullAdder_3728_io_co)
  );
  FullAdder FullAdder_3729 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3729_io_a),
    .io_b(FullAdder_3729_io_b),
    .io_ci(FullAdder_3729_io_ci),
    .io_s(FullAdder_3729_io_s),
    .io_co(FullAdder_3729_io_co)
  );
  FullAdder FullAdder_3730 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3730_io_a),
    .io_b(FullAdder_3730_io_b),
    .io_ci(FullAdder_3730_io_ci),
    .io_s(FullAdder_3730_io_s),
    .io_co(FullAdder_3730_io_co)
  );
  FullAdder FullAdder_3731 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3731_io_a),
    .io_b(FullAdder_3731_io_b),
    .io_ci(FullAdder_3731_io_ci),
    .io_s(FullAdder_3731_io_s),
    .io_co(FullAdder_3731_io_co)
  );
  FullAdder FullAdder_3732 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3732_io_a),
    .io_b(FullAdder_3732_io_b),
    .io_ci(FullAdder_3732_io_ci),
    .io_s(FullAdder_3732_io_s),
    .io_co(FullAdder_3732_io_co)
  );
  FullAdder FullAdder_3733 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3733_io_a),
    .io_b(FullAdder_3733_io_b),
    .io_ci(FullAdder_3733_io_ci),
    .io_s(FullAdder_3733_io_s),
    .io_co(FullAdder_3733_io_co)
  );
  FullAdder FullAdder_3734 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3734_io_a),
    .io_b(FullAdder_3734_io_b),
    .io_ci(FullAdder_3734_io_ci),
    .io_s(FullAdder_3734_io_s),
    .io_co(FullAdder_3734_io_co)
  );
  FullAdder FullAdder_3735 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3735_io_a),
    .io_b(FullAdder_3735_io_b),
    .io_ci(FullAdder_3735_io_ci),
    .io_s(FullAdder_3735_io_s),
    .io_co(FullAdder_3735_io_co)
  );
  FullAdder FullAdder_3736 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3736_io_a),
    .io_b(FullAdder_3736_io_b),
    .io_ci(FullAdder_3736_io_ci),
    .io_s(FullAdder_3736_io_s),
    .io_co(FullAdder_3736_io_co)
  );
  FullAdder FullAdder_3737 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3737_io_a),
    .io_b(FullAdder_3737_io_b),
    .io_ci(FullAdder_3737_io_ci),
    .io_s(FullAdder_3737_io_s),
    .io_co(FullAdder_3737_io_co)
  );
  FullAdder FullAdder_3738 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3738_io_a),
    .io_b(FullAdder_3738_io_b),
    .io_ci(FullAdder_3738_io_ci),
    .io_s(FullAdder_3738_io_s),
    .io_co(FullAdder_3738_io_co)
  );
  FullAdder FullAdder_3739 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3739_io_a),
    .io_b(FullAdder_3739_io_b),
    .io_ci(FullAdder_3739_io_ci),
    .io_s(FullAdder_3739_io_s),
    .io_co(FullAdder_3739_io_co)
  );
  FullAdder FullAdder_3740 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3740_io_a),
    .io_b(FullAdder_3740_io_b),
    .io_ci(FullAdder_3740_io_ci),
    .io_s(FullAdder_3740_io_s),
    .io_co(FullAdder_3740_io_co)
  );
  FullAdder FullAdder_3741 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3741_io_a),
    .io_b(FullAdder_3741_io_b),
    .io_ci(FullAdder_3741_io_ci),
    .io_s(FullAdder_3741_io_s),
    .io_co(FullAdder_3741_io_co)
  );
  FullAdder FullAdder_3742 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3742_io_a),
    .io_b(FullAdder_3742_io_b),
    .io_ci(FullAdder_3742_io_ci),
    .io_s(FullAdder_3742_io_s),
    .io_co(FullAdder_3742_io_co)
  );
  FullAdder FullAdder_3743 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3743_io_a),
    .io_b(FullAdder_3743_io_b),
    .io_ci(FullAdder_3743_io_ci),
    .io_s(FullAdder_3743_io_s),
    .io_co(FullAdder_3743_io_co)
  );
  HalfAdder HalfAdder_218 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_218_io_a),
    .io_b(HalfAdder_218_io_b),
    .io_s(HalfAdder_218_io_s),
    .io_co(HalfAdder_218_io_co)
  );
  HalfAdder HalfAdder_219 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_219_io_a),
    .io_b(HalfAdder_219_io_b),
    .io_s(HalfAdder_219_io_s),
    .io_co(HalfAdder_219_io_co)
  );
  HalfAdder HalfAdder_220 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_220_io_a),
    .io_b(HalfAdder_220_io_b),
    .io_s(HalfAdder_220_io_s),
    .io_co(HalfAdder_220_io_co)
  );
  FullAdder FullAdder_3744 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3744_io_a),
    .io_b(FullAdder_3744_io_b),
    .io_ci(FullAdder_3744_io_ci),
    .io_s(FullAdder_3744_io_s),
    .io_co(FullAdder_3744_io_co)
  );
  HalfAdder HalfAdder_221 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_221_io_a),
    .io_b(HalfAdder_221_io_b),
    .io_s(HalfAdder_221_io_s),
    .io_co(HalfAdder_221_io_co)
  );
  FullAdder FullAdder_3745 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3745_io_a),
    .io_b(FullAdder_3745_io_b),
    .io_ci(FullAdder_3745_io_ci),
    .io_s(FullAdder_3745_io_s),
    .io_co(FullAdder_3745_io_co)
  );
  FullAdder FullAdder_3746 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3746_io_a),
    .io_b(FullAdder_3746_io_b),
    .io_ci(FullAdder_3746_io_ci),
    .io_s(FullAdder_3746_io_s),
    .io_co(FullAdder_3746_io_co)
  );
  FullAdder FullAdder_3747 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3747_io_a),
    .io_b(FullAdder_3747_io_b),
    .io_ci(FullAdder_3747_io_ci),
    .io_s(FullAdder_3747_io_s),
    .io_co(FullAdder_3747_io_co)
  );
  FullAdder FullAdder_3748 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3748_io_a),
    .io_b(FullAdder_3748_io_b),
    .io_ci(FullAdder_3748_io_ci),
    .io_s(FullAdder_3748_io_s),
    .io_co(FullAdder_3748_io_co)
  );
  FullAdder FullAdder_3749 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3749_io_a),
    .io_b(FullAdder_3749_io_b),
    .io_ci(FullAdder_3749_io_ci),
    .io_s(FullAdder_3749_io_s),
    .io_co(FullAdder_3749_io_co)
  );
  FullAdder FullAdder_3750 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3750_io_a),
    .io_b(FullAdder_3750_io_b),
    .io_ci(FullAdder_3750_io_ci),
    .io_s(FullAdder_3750_io_s),
    .io_co(FullAdder_3750_io_co)
  );
  FullAdder FullAdder_3751 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3751_io_a),
    .io_b(FullAdder_3751_io_b),
    .io_ci(FullAdder_3751_io_ci),
    .io_s(FullAdder_3751_io_s),
    .io_co(FullAdder_3751_io_co)
  );
  FullAdder FullAdder_3752 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3752_io_a),
    .io_b(FullAdder_3752_io_b),
    .io_ci(FullAdder_3752_io_ci),
    .io_s(FullAdder_3752_io_s),
    .io_co(FullAdder_3752_io_co)
  );
  FullAdder FullAdder_3753 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3753_io_a),
    .io_b(FullAdder_3753_io_b),
    .io_ci(FullAdder_3753_io_ci),
    .io_s(FullAdder_3753_io_s),
    .io_co(FullAdder_3753_io_co)
  );
  FullAdder FullAdder_3754 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3754_io_a),
    .io_b(FullAdder_3754_io_b),
    .io_ci(FullAdder_3754_io_ci),
    .io_s(FullAdder_3754_io_s),
    .io_co(FullAdder_3754_io_co)
  );
  FullAdder FullAdder_3755 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3755_io_a),
    .io_b(FullAdder_3755_io_b),
    .io_ci(FullAdder_3755_io_ci),
    .io_s(FullAdder_3755_io_s),
    .io_co(FullAdder_3755_io_co)
  );
  FullAdder FullAdder_3756 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3756_io_a),
    .io_b(FullAdder_3756_io_b),
    .io_ci(FullAdder_3756_io_ci),
    .io_s(FullAdder_3756_io_s),
    .io_co(FullAdder_3756_io_co)
  );
  FullAdder FullAdder_3757 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3757_io_a),
    .io_b(FullAdder_3757_io_b),
    .io_ci(FullAdder_3757_io_ci),
    .io_s(FullAdder_3757_io_s),
    .io_co(FullAdder_3757_io_co)
  );
  FullAdder FullAdder_3758 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3758_io_a),
    .io_b(FullAdder_3758_io_b),
    .io_ci(FullAdder_3758_io_ci),
    .io_s(FullAdder_3758_io_s),
    .io_co(FullAdder_3758_io_co)
  );
  FullAdder FullAdder_3759 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3759_io_a),
    .io_b(FullAdder_3759_io_b),
    .io_ci(FullAdder_3759_io_ci),
    .io_s(FullAdder_3759_io_s),
    .io_co(FullAdder_3759_io_co)
  );
  FullAdder FullAdder_3760 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3760_io_a),
    .io_b(FullAdder_3760_io_b),
    .io_ci(FullAdder_3760_io_ci),
    .io_s(FullAdder_3760_io_s),
    .io_co(FullAdder_3760_io_co)
  );
  FullAdder FullAdder_3761 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3761_io_a),
    .io_b(FullAdder_3761_io_b),
    .io_ci(FullAdder_3761_io_ci),
    .io_s(FullAdder_3761_io_s),
    .io_co(FullAdder_3761_io_co)
  );
  FullAdder FullAdder_3762 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3762_io_a),
    .io_b(FullAdder_3762_io_b),
    .io_ci(FullAdder_3762_io_ci),
    .io_s(FullAdder_3762_io_s),
    .io_co(FullAdder_3762_io_co)
  );
  FullAdder FullAdder_3763 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3763_io_a),
    .io_b(FullAdder_3763_io_b),
    .io_ci(FullAdder_3763_io_ci),
    .io_s(FullAdder_3763_io_s),
    .io_co(FullAdder_3763_io_co)
  );
  FullAdder FullAdder_3764 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3764_io_a),
    .io_b(FullAdder_3764_io_b),
    .io_ci(FullAdder_3764_io_ci),
    .io_s(FullAdder_3764_io_s),
    .io_co(FullAdder_3764_io_co)
  );
  FullAdder FullAdder_3765 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3765_io_a),
    .io_b(FullAdder_3765_io_b),
    .io_ci(FullAdder_3765_io_ci),
    .io_s(FullAdder_3765_io_s),
    .io_co(FullAdder_3765_io_co)
  );
  FullAdder FullAdder_3766 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3766_io_a),
    .io_b(FullAdder_3766_io_b),
    .io_ci(FullAdder_3766_io_ci),
    .io_s(FullAdder_3766_io_s),
    .io_co(FullAdder_3766_io_co)
  );
  FullAdder FullAdder_3767 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3767_io_a),
    .io_b(FullAdder_3767_io_b),
    .io_ci(FullAdder_3767_io_ci),
    .io_s(FullAdder_3767_io_s),
    .io_co(FullAdder_3767_io_co)
  );
  FullAdder FullAdder_3768 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3768_io_a),
    .io_b(FullAdder_3768_io_b),
    .io_ci(FullAdder_3768_io_ci),
    .io_s(FullAdder_3768_io_s),
    .io_co(FullAdder_3768_io_co)
  );
  HalfAdder HalfAdder_222 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_222_io_a),
    .io_b(HalfAdder_222_io_b),
    .io_s(HalfAdder_222_io_s),
    .io_co(HalfAdder_222_io_co)
  );
  FullAdder FullAdder_3769 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3769_io_a),
    .io_b(FullAdder_3769_io_b),
    .io_ci(FullAdder_3769_io_ci),
    .io_s(FullAdder_3769_io_s),
    .io_co(FullAdder_3769_io_co)
  );
  FullAdder FullAdder_3770 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3770_io_a),
    .io_b(FullAdder_3770_io_b),
    .io_ci(FullAdder_3770_io_ci),
    .io_s(FullAdder_3770_io_s),
    .io_co(FullAdder_3770_io_co)
  );
  FullAdder FullAdder_3771 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3771_io_a),
    .io_b(FullAdder_3771_io_b),
    .io_ci(FullAdder_3771_io_ci),
    .io_s(FullAdder_3771_io_s),
    .io_co(FullAdder_3771_io_co)
  );
  FullAdder FullAdder_3772 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3772_io_a),
    .io_b(FullAdder_3772_io_b),
    .io_ci(FullAdder_3772_io_ci),
    .io_s(FullAdder_3772_io_s),
    .io_co(FullAdder_3772_io_co)
  );
  HalfAdder HalfAdder_223 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_223_io_a),
    .io_b(HalfAdder_223_io_b),
    .io_s(HalfAdder_223_io_s),
    .io_co(HalfAdder_223_io_co)
  );
  FullAdder FullAdder_3773 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3773_io_a),
    .io_b(FullAdder_3773_io_b),
    .io_ci(FullAdder_3773_io_ci),
    .io_s(FullAdder_3773_io_s),
    .io_co(FullAdder_3773_io_co)
  );
  HalfAdder HalfAdder_224 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_224_io_a),
    .io_b(HalfAdder_224_io_b),
    .io_s(HalfAdder_224_io_s),
    .io_co(HalfAdder_224_io_co)
  );
  FullAdder FullAdder_3774 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3774_io_a),
    .io_b(FullAdder_3774_io_b),
    .io_ci(FullAdder_3774_io_ci),
    .io_s(FullAdder_3774_io_s),
    .io_co(FullAdder_3774_io_co)
  );
  HalfAdder HalfAdder_225 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_225_io_a),
    .io_b(HalfAdder_225_io_b),
    .io_s(HalfAdder_225_io_s),
    .io_co(HalfAdder_225_io_co)
  );
  FullAdder FullAdder_3775 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3775_io_a),
    .io_b(FullAdder_3775_io_b),
    .io_ci(FullAdder_3775_io_ci),
    .io_s(FullAdder_3775_io_s),
    .io_co(FullAdder_3775_io_co)
  );
  FullAdder FullAdder_3776 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3776_io_a),
    .io_b(FullAdder_3776_io_b),
    .io_ci(FullAdder_3776_io_ci),
    .io_s(FullAdder_3776_io_s),
    .io_co(FullAdder_3776_io_co)
  );
  HalfAdder HalfAdder_226 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_226_io_a),
    .io_b(HalfAdder_226_io_b),
    .io_s(HalfAdder_226_io_s),
    .io_co(HalfAdder_226_io_co)
  );
  FullAdder FullAdder_3777 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3777_io_a),
    .io_b(FullAdder_3777_io_b),
    .io_ci(FullAdder_3777_io_ci),
    .io_s(FullAdder_3777_io_s),
    .io_co(FullAdder_3777_io_co)
  );
  FullAdder FullAdder_3778 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3778_io_a),
    .io_b(FullAdder_3778_io_b),
    .io_ci(FullAdder_3778_io_ci),
    .io_s(FullAdder_3778_io_s),
    .io_co(FullAdder_3778_io_co)
  );
  FullAdder FullAdder_3779 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3779_io_a),
    .io_b(FullAdder_3779_io_b),
    .io_ci(FullAdder_3779_io_ci),
    .io_s(FullAdder_3779_io_s),
    .io_co(FullAdder_3779_io_co)
  );
  FullAdder FullAdder_3780 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3780_io_a),
    .io_b(FullAdder_3780_io_b),
    .io_ci(FullAdder_3780_io_ci),
    .io_s(FullAdder_3780_io_s),
    .io_co(FullAdder_3780_io_co)
  );
  FullAdder FullAdder_3781 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3781_io_a),
    .io_b(FullAdder_3781_io_b),
    .io_ci(FullAdder_3781_io_ci),
    .io_s(FullAdder_3781_io_s),
    .io_co(FullAdder_3781_io_co)
  );
  HalfAdder HalfAdder_227 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_227_io_a),
    .io_b(HalfAdder_227_io_b),
    .io_s(HalfAdder_227_io_s),
    .io_co(HalfAdder_227_io_co)
  );
  FullAdder FullAdder_3782 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3782_io_a),
    .io_b(FullAdder_3782_io_b),
    .io_ci(FullAdder_3782_io_ci),
    .io_s(FullAdder_3782_io_s),
    .io_co(FullAdder_3782_io_co)
  );
  HalfAdder HalfAdder_228 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_228_io_a),
    .io_b(HalfAdder_228_io_b),
    .io_s(HalfAdder_228_io_s),
    .io_co(HalfAdder_228_io_co)
  );
  HalfAdder HalfAdder_229 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_229_io_a),
    .io_b(HalfAdder_229_io_b),
    .io_s(HalfAdder_229_io_s),
    .io_co(HalfAdder_229_io_co)
  );
  FullAdder FullAdder_3783 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3783_io_a),
    .io_b(FullAdder_3783_io_b),
    .io_ci(FullAdder_3783_io_ci),
    .io_s(FullAdder_3783_io_s),
    .io_co(FullAdder_3783_io_co)
  );
  FullAdder FullAdder_3784 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3784_io_a),
    .io_b(FullAdder_3784_io_b),
    .io_ci(FullAdder_3784_io_ci),
    .io_s(FullAdder_3784_io_s),
    .io_co(FullAdder_3784_io_co)
  );
  FullAdder FullAdder_3785 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3785_io_a),
    .io_b(FullAdder_3785_io_b),
    .io_ci(FullAdder_3785_io_ci),
    .io_s(FullAdder_3785_io_s),
    .io_co(FullAdder_3785_io_co)
  );
  FullAdder FullAdder_3786 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3786_io_a),
    .io_b(FullAdder_3786_io_b),
    .io_ci(FullAdder_3786_io_ci),
    .io_s(FullAdder_3786_io_s),
    .io_co(FullAdder_3786_io_co)
  );
  HalfAdder HalfAdder_230 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_230_io_a),
    .io_b(HalfAdder_230_io_b),
    .io_s(HalfAdder_230_io_s),
    .io_co(HalfAdder_230_io_co)
  );
  FullAdder FullAdder_3787 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3787_io_a),
    .io_b(FullAdder_3787_io_b),
    .io_ci(FullAdder_3787_io_ci),
    .io_s(FullAdder_3787_io_s),
    .io_co(FullAdder_3787_io_co)
  );
  HalfAdder HalfAdder_231 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_231_io_a),
    .io_b(HalfAdder_231_io_b),
    .io_s(HalfAdder_231_io_s),
    .io_co(HalfAdder_231_io_co)
  );
  FullAdder FullAdder_3788 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3788_io_a),
    .io_b(FullAdder_3788_io_b),
    .io_ci(FullAdder_3788_io_ci),
    .io_s(FullAdder_3788_io_s),
    .io_co(FullAdder_3788_io_co)
  );
  FullAdder FullAdder_3789 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3789_io_a),
    .io_b(FullAdder_3789_io_b),
    .io_ci(FullAdder_3789_io_ci),
    .io_s(FullAdder_3789_io_s),
    .io_co(FullAdder_3789_io_co)
  );
  FullAdder FullAdder_3790 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3790_io_a),
    .io_b(FullAdder_3790_io_b),
    .io_ci(FullAdder_3790_io_ci),
    .io_s(FullAdder_3790_io_s),
    .io_co(FullAdder_3790_io_co)
  );
  HalfAdder HalfAdder_232 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_232_io_a),
    .io_b(HalfAdder_232_io_b),
    .io_s(HalfAdder_232_io_s),
    .io_co(HalfAdder_232_io_co)
  );
  FullAdder FullAdder_3791 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3791_io_a),
    .io_b(FullAdder_3791_io_b),
    .io_ci(FullAdder_3791_io_ci),
    .io_s(FullAdder_3791_io_s),
    .io_co(FullAdder_3791_io_co)
  );
  FullAdder FullAdder_3792 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3792_io_a),
    .io_b(FullAdder_3792_io_b),
    .io_ci(FullAdder_3792_io_ci),
    .io_s(FullAdder_3792_io_s),
    .io_co(FullAdder_3792_io_co)
  );
  FullAdder FullAdder_3793 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3793_io_a),
    .io_b(FullAdder_3793_io_b),
    .io_ci(FullAdder_3793_io_ci),
    .io_s(FullAdder_3793_io_s),
    .io_co(FullAdder_3793_io_co)
  );
  HalfAdder HalfAdder_233 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_233_io_a),
    .io_b(HalfAdder_233_io_b),
    .io_s(HalfAdder_233_io_s),
    .io_co(HalfAdder_233_io_co)
  );
  FullAdder FullAdder_3794 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3794_io_a),
    .io_b(FullAdder_3794_io_b),
    .io_ci(FullAdder_3794_io_ci),
    .io_s(FullAdder_3794_io_s),
    .io_co(FullAdder_3794_io_co)
  );
  HalfAdder HalfAdder_234 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_234_io_a),
    .io_b(HalfAdder_234_io_b),
    .io_s(HalfAdder_234_io_s),
    .io_co(HalfAdder_234_io_co)
  );
  FullAdder FullAdder_3795 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3795_io_a),
    .io_b(FullAdder_3795_io_b),
    .io_ci(FullAdder_3795_io_ci),
    .io_s(FullAdder_3795_io_s),
    .io_co(FullAdder_3795_io_co)
  );
  FullAdder FullAdder_3796 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3796_io_a),
    .io_b(FullAdder_3796_io_b),
    .io_ci(FullAdder_3796_io_ci),
    .io_s(FullAdder_3796_io_s),
    .io_co(FullAdder_3796_io_co)
  );
  HalfAdder HalfAdder_235 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_235_io_a),
    .io_b(HalfAdder_235_io_b),
    .io_s(HalfAdder_235_io_s),
    .io_co(HalfAdder_235_io_co)
  );
  FullAdder FullAdder_3797 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3797_io_a),
    .io_b(FullAdder_3797_io_b),
    .io_ci(FullAdder_3797_io_ci),
    .io_s(FullAdder_3797_io_s),
    .io_co(FullAdder_3797_io_co)
  );
  FullAdder FullAdder_3798 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3798_io_a),
    .io_b(FullAdder_3798_io_b),
    .io_ci(FullAdder_3798_io_ci),
    .io_s(FullAdder_3798_io_s),
    .io_co(FullAdder_3798_io_co)
  );
  FullAdder FullAdder_3799 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3799_io_a),
    .io_b(FullAdder_3799_io_b),
    .io_ci(FullAdder_3799_io_ci),
    .io_s(FullAdder_3799_io_s),
    .io_co(FullAdder_3799_io_co)
  );
  FullAdder FullAdder_3800 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3800_io_a),
    .io_b(FullAdder_3800_io_b),
    .io_ci(FullAdder_3800_io_ci),
    .io_s(FullAdder_3800_io_s),
    .io_co(FullAdder_3800_io_co)
  );
  FullAdder FullAdder_3801 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3801_io_a),
    .io_b(FullAdder_3801_io_b),
    .io_ci(FullAdder_3801_io_ci),
    .io_s(FullAdder_3801_io_s),
    .io_co(FullAdder_3801_io_co)
  );
  FullAdder FullAdder_3802 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3802_io_a),
    .io_b(FullAdder_3802_io_b),
    .io_ci(FullAdder_3802_io_ci),
    .io_s(FullAdder_3802_io_s),
    .io_co(FullAdder_3802_io_co)
  );
  FullAdder FullAdder_3803 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3803_io_a),
    .io_b(FullAdder_3803_io_b),
    .io_ci(FullAdder_3803_io_ci),
    .io_s(FullAdder_3803_io_s),
    .io_co(FullAdder_3803_io_co)
  );
  FullAdder FullAdder_3804 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3804_io_a),
    .io_b(FullAdder_3804_io_b),
    .io_ci(FullAdder_3804_io_ci),
    .io_s(FullAdder_3804_io_s),
    .io_co(FullAdder_3804_io_co)
  );
  FullAdder FullAdder_3805 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3805_io_a),
    .io_b(FullAdder_3805_io_b),
    .io_ci(FullAdder_3805_io_ci),
    .io_s(FullAdder_3805_io_s),
    .io_co(FullAdder_3805_io_co)
  );
  FullAdder FullAdder_3806 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3806_io_a),
    .io_b(FullAdder_3806_io_b),
    .io_ci(FullAdder_3806_io_ci),
    .io_s(FullAdder_3806_io_s),
    .io_co(FullAdder_3806_io_co)
  );
  FullAdder FullAdder_3807 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3807_io_a),
    .io_b(FullAdder_3807_io_b),
    .io_ci(FullAdder_3807_io_ci),
    .io_s(FullAdder_3807_io_s),
    .io_co(FullAdder_3807_io_co)
  );
  FullAdder FullAdder_3808 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3808_io_a),
    .io_b(FullAdder_3808_io_b),
    .io_ci(FullAdder_3808_io_ci),
    .io_s(FullAdder_3808_io_s),
    .io_co(FullAdder_3808_io_co)
  );
  FullAdder FullAdder_3809 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3809_io_a),
    .io_b(FullAdder_3809_io_b),
    .io_ci(FullAdder_3809_io_ci),
    .io_s(FullAdder_3809_io_s),
    .io_co(FullAdder_3809_io_co)
  );
  FullAdder FullAdder_3810 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3810_io_a),
    .io_b(FullAdder_3810_io_b),
    .io_ci(FullAdder_3810_io_ci),
    .io_s(FullAdder_3810_io_s),
    .io_co(FullAdder_3810_io_co)
  );
  FullAdder FullAdder_3811 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3811_io_a),
    .io_b(FullAdder_3811_io_b),
    .io_ci(FullAdder_3811_io_ci),
    .io_s(FullAdder_3811_io_s),
    .io_co(FullAdder_3811_io_co)
  );
  HalfAdder HalfAdder_236 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_236_io_a),
    .io_b(HalfAdder_236_io_b),
    .io_s(HalfAdder_236_io_s),
    .io_co(HalfAdder_236_io_co)
  );
  HalfAdder HalfAdder_237 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_237_io_a),
    .io_b(HalfAdder_237_io_b),
    .io_s(HalfAdder_237_io_s),
    .io_co(HalfAdder_237_io_co)
  );
  HalfAdder HalfAdder_238 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_238_io_a),
    .io_b(HalfAdder_238_io_b),
    .io_s(HalfAdder_238_io_s),
    .io_co(HalfAdder_238_io_co)
  );
  FullAdder FullAdder_3812 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3812_io_a),
    .io_b(FullAdder_3812_io_b),
    .io_ci(FullAdder_3812_io_ci),
    .io_s(FullAdder_3812_io_s),
    .io_co(FullAdder_3812_io_co)
  );
  FullAdder FullAdder_3813 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3813_io_a),
    .io_b(FullAdder_3813_io_b),
    .io_ci(FullAdder_3813_io_ci),
    .io_s(FullAdder_3813_io_s),
    .io_co(FullAdder_3813_io_co)
  );
  FullAdder FullAdder_3814 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3814_io_a),
    .io_b(FullAdder_3814_io_b),
    .io_ci(FullAdder_3814_io_ci),
    .io_s(FullAdder_3814_io_s),
    .io_co(FullAdder_3814_io_co)
  );
  FullAdder FullAdder_3815 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3815_io_a),
    .io_b(FullAdder_3815_io_b),
    .io_ci(FullAdder_3815_io_ci),
    .io_s(FullAdder_3815_io_s),
    .io_co(FullAdder_3815_io_co)
  );
  HalfAdder HalfAdder_239 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_239_io_a),
    .io_b(HalfAdder_239_io_b),
    .io_s(HalfAdder_239_io_s),
    .io_co(HalfAdder_239_io_co)
  );
  FullAdder FullAdder_3816 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3816_io_a),
    .io_b(FullAdder_3816_io_b),
    .io_ci(FullAdder_3816_io_ci),
    .io_s(FullAdder_3816_io_s),
    .io_co(FullAdder_3816_io_co)
  );
  FullAdder FullAdder_3817 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3817_io_a),
    .io_b(FullAdder_3817_io_b),
    .io_ci(FullAdder_3817_io_ci),
    .io_s(FullAdder_3817_io_s),
    .io_co(FullAdder_3817_io_co)
  );
  FullAdder FullAdder_3818 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3818_io_a),
    .io_b(FullAdder_3818_io_b),
    .io_ci(FullAdder_3818_io_ci),
    .io_s(FullAdder_3818_io_s),
    .io_co(FullAdder_3818_io_co)
  );
  FullAdder FullAdder_3819 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3819_io_a),
    .io_b(FullAdder_3819_io_b),
    .io_ci(FullAdder_3819_io_ci),
    .io_s(FullAdder_3819_io_s),
    .io_co(FullAdder_3819_io_co)
  );
  FullAdder FullAdder_3820 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3820_io_a),
    .io_b(FullAdder_3820_io_b),
    .io_ci(FullAdder_3820_io_ci),
    .io_s(FullAdder_3820_io_s),
    .io_co(FullAdder_3820_io_co)
  );
  FullAdder FullAdder_3821 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3821_io_a),
    .io_b(FullAdder_3821_io_b),
    .io_ci(FullAdder_3821_io_ci),
    .io_s(FullAdder_3821_io_s),
    .io_co(FullAdder_3821_io_co)
  );
  FullAdder FullAdder_3822 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3822_io_a),
    .io_b(FullAdder_3822_io_b),
    .io_ci(FullAdder_3822_io_ci),
    .io_s(FullAdder_3822_io_s),
    .io_co(FullAdder_3822_io_co)
  );
  HalfAdder HalfAdder_240 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_240_io_a),
    .io_b(HalfAdder_240_io_b),
    .io_s(HalfAdder_240_io_s),
    .io_co(HalfAdder_240_io_co)
  );
  FullAdder FullAdder_3823 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3823_io_a),
    .io_b(FullAdder_3823_io_b),
    .io_ci(FullAdder_3823_io_ci),
    .io_s(FullAdder_3823_io_s),
    .io_co(FullAdder_3823_io_co)
  );
  FullAdder FullAdder_3824 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3824_io_a),
    .io_b(FullAdder_3824_io_b),
    .io_ci(FullAdder_3824_io_ci),
    .io_s(FullAdder_3824_io_s),
    .io_co(FullAdder_3824_io_co)
  );
  HalfAdder HalfAdder_241 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_241_io_a),
    .io_b(HalfAdder_241_io_b),
    .io_s(HalfAdder_241_io_s),
    .io_co(HalfAdder_241_io_co)
  );
  FullAdder FullAdder_3825 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3825_io_a),
    .io_b(FullAdder_3825_io_b),
    .io_ci(FullAdder_3825_io_ci),
    .io_s(FullAdder_3825_io_s),
    .io_co(FullAdder_3825_io_co)
  );
  FullAdder FullAdder_3826 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3826_io_a),
    .io_b(FullAdder_3826_io_b),
    .io_ci(FullAdder_3826_io_ci),
    .io_s(FullAdder_3826_io_s),
    .io_co(FullAdder_3826_io_co)
  );
  FullAdder FullAdder_3827 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3827_io_a),
    .io_b(FullAdder_3827_io_b),
    .io_ci(FullAdder_3827_io_ci),
    .io_s(FullAdder_3827_io_s),
    .io_co(FullAdder_3827_io_co)
  );
  HalfAdder HalfAdder_242 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_242_io_a),
    .io_b(HalfAdder_242_io_b),
    .io_s(HalfAdder_242_io_s),
    .io_co(HalfAdder_242_io_co)
  );
  FullAdder FullAdder_3828 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3828_io_a),
    .io_b(FullAdder_3828_io_b),
    .io_ci(FullAdder_3828_io_ci),
    .io_s(FullAdder_3828_io_s),
    .io_co(FullAdder_3828_io_co)
  );
  FullAdder FullAdder_3829 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3829_io_a),
    .io_b(FullAdder_3829_io_b),
    .io_ci(FullAdder_3829_io_ci),
    .io_s(FullAdder_3829_io_s),
    .io_co(FullAdder_3829_io_co)
  );
  HalfAdder HalfAdder_243 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_243_io_a),
    .io_b(HalfAdder_243_io_b),
    .io_s(HalfAdder_243_io_s),
    .io_co(HalfAdder_243_io_co)
  );
  FullAdder FullAdder_3830 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3830_io_a),
    .io_b(FullAdder_3830_io_b),
    .io_ci(FullAdder_3830_io_ci),
    .io_s(FullAdder_3830_io_s),
    .io_co(FullAdder_3830_io_co)
  );
  HalfAdder HalfAdder_244 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_244_io_a),
    .io_b(HalfAdder_244_io_b),
    .io_s(HalfAdder_244_io_s),
    .io_co(HalfAdder_244_io_co)
  );
  FullAdder FullAdder_3831 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3831_io_a),
    .io_b(FullAdder_3831_io_b),
    .io_ci(FullAdder_3831_io_ci),
    .io_s(FullAdder_3831_io_s),
    .io_co(FullAdder_3831_io_co)
  );
  HalfAdder HalfAdder_245 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_245_io_a),
    .io_b(HalfAdder_245_io_b),
    .io_s(HalfAdder_245_io_s),
    .io_co(HalfAdder_245_io_co)
  );
  HalfAdder HalfAdder_246 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_246_io_a),
    .io_b(HalfAdder_246_io_b),
    .io_s(HalfAdder_246_io_s),
    .io_co(HalfAdder_246_io_co)
  );
  HalfAdder HalfAdder_247 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_247_io_a),
    .io_b(HalfAdder_247_io_b),
    .io_s(HalfAdder_247_io_s),
    .io_co(HalfAdder_247_io_co)
  );
  FullAdder FullAdder_3832 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3832_io_a),
    .io_b(FullAdder_3832_io_b),
    .io_ci(FullAdder_3832_io_ci),
    .io_s(FullAdder_3832_io_s),
    .io_co(FullAdder_3832_io_co)
  );
  FullAdder FullAdder_3833 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3833_io_a),
    .io_b(FullAdder_3833_io_b),
    .io_ci(FullAdder_3833_io_ci),
    .io_s(FullAdder_3833_io_s),
    .io_co(FullAdder_3833_io_co)
  );
  HalfAdder HalfAdder_248 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_248_io_a),
    .io_b(HalfAdder_248_io_b),
    .io_s(HalfAdder_248_io_s),
    .io_co(HalfAdder_248_io_co)
  );
  FullAdder FullAdder_3834 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3834_io_a),
    .io_b(FullAdder_3834_io_b),
    .io_ci(FullAdder_3834_io_ci),
    .io_s(FullAdder_3834_io_s),
    .io_co(FullAdder_3834_io_co)
  );
  FullAdder FullAdder_3835 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3835_io_a),
    .io_b(FullAdder_3835_io_b),
    .io_ci(FullAdder_3835_io_ci),
    .io_s(FullAdder_3835_io_s),
    .io_co(FullAdder_3835_io_co)
  );
  FullAdder FullAdder_3836 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3836_io_a),
    .io_b(FullAdder_3836_io_b),
    .io_ci(FullAdder_3836_io_ci),
    .io_s(FullAdder_3836_io_s),
    .io_co(FullAdder_3836_io_co)
  );
  FullAdder FullAdder_3837 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3837_io_a),
    .io_b(FullAdder_3837_io_b),
    .io_ci(FullAdder_3837_io_ci),
    .io_s(FullAdder_3837_io_s),
    .io_co(FullAdder_3837_io_co)
  );
  FullAdder FullAdder_3838 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3838_io_a),
    .io_b(FullAdder_3838_io_b),
    .io_ci(FullAdder_3838_io_ci),
    .io_s(FullAdder_3838_io_s),
    .io_co(FullAdder_3838_io_co)
  );
  HalfAdder HalfAdder_249 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_249_io_a),
    .io_b(HalfAdder_249_io_b),
    .io_s(HalfAdder_249_io_s),
    .io_co(HalfAdder_249_io_co)
  );
  FullAdder FullAdder_3839 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3839_io_a),
    .io_b(FullAdder_3839_io_b),
    .io_ci(FullAdder_3839_io_ci),
    .io_s(FullAdder_3839_io_s),
    .io_co(FullAdder_3839_io_co)
  );
  FullAdder FullAdder_3840 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3840_io_a),
    .io_b(FullAdder_3840_io_b),
    .io_ci(FullAdder_3840_io_ci),
    .io_s(FullAdder_3840_io_s),
    .io_co(FullAdder_3840_io_co)
  );
  FullAdder FullAdder_3841 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3841_io_a),
    .io_b(FullAdder_3841_io_b),
    .io_ci(FullAdder_3841_io_ci),
    .io_s(FullAdder_3841_io_s),
    .io_co(FullAdder_3841_io_co)
  );
  HalfAdder HalfAdder_250 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_250_io_a),
    .io_b(HalfAdder_250_io_b),
    .io_s(HalfAdder_250_io_s),
    .io_co(HalfAdder_250_io_co)
  );
  FullAdder FullAdder_3842 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3842_io_a),
    .io_b(FullAdder_3842_io_b),
    .io_ci(FullAdder_3842_io_ci),
    .io_s(FullAdder_3842_io_s),
    .io_co(FullAdder_3842_io_co)
  );
  FullAdder FullAdder_3843 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3843_io_a),
    .io_b(FullAdder_3843_io_b),
    .io_ci(FullAdder_3843_io_ci),
    .io_s(FullAdder_3843_io_s),
    .io_co(FullAdder_3843_io_co)
  );
  FullAdder FullAdder_3844 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3844_io_a),
    .io_b(FullAdder_3844_io_b),
    .io_ci(FullAdder_3844_io_ci),
    .io_s(FullAdder_3844_io_s),
    .io_co(FullAdder_3844_io_co)
  );
  HalfAdder HalfAdder_251 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_251_io_a),
    .io_b(HalfAdder_251_io_b),
    .io_s(HalfAdder_251_io_s),
    .io_co(HalfAdder_251_io_co)
  );
  HalfAdder HalfAdder_252 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_252_io_a),
    .io_b(HalfAdder_252_io_b),
    .io_s(HalfAdder_252_io_s),
    .io_co(HalfAdder_252_io_co)
  );
  FullAdder FullAdder_3845 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3845_io_a),
    .io_b(FullAdder_3845_io_b),
    .io_ci(FullAdder_3845_io_ci),
    .io_s(FullAdder_3845_io_s),
    .io_co(FullAdder_3845_io_co)
  );
  HalfAdder HalfAdder_253 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_253_io_a),
    .io_b(HalfAdder_253_io_b),
    .io_s(HalfAdder_253_io_s),
    .io_co(HalfAdder_253_io_co)
  );
  FullAdder FullAdder_3846 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3846_io_a),
    .io_b(FullAdder_3846_io_b),
    .io_ci(FullAdder_3846_io_ci),
    .io_s(FullAdder_3846_io_s),
    .io_co(FullAdder_3846_io_co)
  );
  FullAdder FullAdder_3847 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3847_io_a),
    .io_b(FullAdder_3847_io_b),
    .io_ci(FullAdder_3847_io_ci),
    .io_s(FullAdder_3847_io_s),
    .io_co(FullAdder_3847_io_co)
  );
  HalfAdder HalfAdder_254 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_254_io_a),
    .io_b(HalfAdder_254_io_b),
    .io_s(HalfAdder_254_io_s),
    .io_co(HalfAdder_254_io_co)
  );
  FullAdder FullAdder_3848 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3848_io_a),
    .io_b(FullAdder_3848_io_b),
    .io_ci(FullAdder_3848_io_ci),
    .io_s(FullAdder_3848_io_s),
    .io_co(FullAdder_3848_io_co)
  );
  FullAdder FullAdder_3849 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3849_io_a),
    .io_b(FullAdder_3849_io_b),
    .io_ci(FullAdder_3849_io_ci),
    .io_s(FullAdder_3849_io_s),
    .io_co(FullAdder_3849_io_co)
  );
  HalfAdder HalfAdder_255 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_255_io_a),
    .io_b(HalfAdder_255_io_b),
    .io_s(HalfAdder_255_io_s),
    .io_co(HalfAdder_255_io_co)
  );
  HalfAdder HalfAdder_256 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_256_io_a),
    .io_b(HalfAdder_256_io_b),
    .io_s(HalfAdder_256_io_s),
    .io_co(HalfAdder_256_io_co)
  );
  FullAdder FullAdder_3850 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3850_io_a),
    .io_b(FullAdder_3850_io_b),
    .io_ci(FullAdder_3850_io_ci),
    .io_s(FullAdder_3850_io_s),
    .io_co(FullAdder_3850_io_co)
  );
  FullAdder FullAdder_3851 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3851_io_a),
    .io_b(FullAdder_3851_io_b),
    .io_ci(FullAdder_3851_io_ci),
    .io_s(FullAdder_3851_io_s),
    .io_co(FullAdder_3851_io_co)
  );
  FullAdder FullAdder_3852 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3852_io_a),
    .io_b(FullAdder_3852_io_b),
    .io_ci(FullAdder_3852_io_ci),
    .io_s(FullAdder_3852_io_s),
    .io_co(FullAdder_3852_io_co)
  );
  HalfAdder HalfAdder_257 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_257_io_a),
    .io_b(HalfAdder_257_io_b),
    .io_s(HalfAdder_257_io_s),
    .io_co(HalfAdder_257_io_co)
  );
  HalfAdder HalfAdder_258 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_258_io_a),
    .io_b(HalfAdder_258_io_b),
    .io_s(HalfAdder_258_io_s),
    .io_co(HalfAdder_258_io_co)
  );
  HalfAdder HalfAdder_259 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_259_io_a),
    .io_b(HalfAdder_259_io_b),
    .io_s(HalfAdder_259_io_s),
    .io_co(HalfAdder_259_io_co)
  );
  HalfAdder HalfAdder_260 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_260_io_a),
    .io_b(HalfAdder_260_io_b),
    .io_s(HalfAdder_260_io_s),
    .io_co(HalfAdder_260_io_co)
  );
  HalfAdder HalfAdder_261 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_261_io_a),
    .io_b(HalfAdder_261_io_b),
    .io_s(HalfAdder_261_io_s),
    .io_co(HalfAdder_261_io_co)
  );
  FullAdder FullAdder_3853 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3853_io_a),
    .io_b(FullAdder_3853_io_b),
    .io_ci(FullAdder_3853_io_ci),
    .io_s(FullAdder_3853_io_s),
    .io_co(FullAdder_3853_io_co)
  );
  FullAdder FullAdder_3854 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3854_io_a),
    .io_b(FullAdder_3854_io_b),
    .io_ci(FullAdder_3854_io_ci),
    .io_s(FullAdder_3854_io_s),
    .io_co(FullAdder_3854_io_co)
  );
  FullAdder FullAdder_3855 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3855_io_a),
    .io_b(FullAdder_3855_io_b),
    .io_ci(FullAdder_3855_io_ci),
    .io_s(FullAdder_3855_io_s),
    .io_co(FullAdder_3855_io_co)
  );
  FullAdder FullAdder_3856 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3856_io_a),
    .io_b(FullAdder_3856_io_b),
    .io_ci(FullAdder_3856_io_ci),
    .io_s(FullAdder_3856_io_s),
    .io_co(FullAdder_3856_io_co)
  );
  FullAdder FullAdder_3857 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3857_io_a),
    .io_b(FullAdder_3857_io_b),
    .io_ci(FullAdder_3857_io_ci),
    .io_s(FullAdder_3857_io_s),
    .io_co(FullAdder_3857_io_co)
  );
  FullAdder FullAdder_3858 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3858_io_a),
    .io_b(FullAdder_3858_io_b),
    .io_ci(FullAdder_3858_io_ci),
    .io_s(FullAdder_3858_io_s),
    .io_co(FullAdder_3858_io_co)
  );
  FullAdder FullAdder_3859 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3859_io_a),
    .io_b(FullAdder_3859_io_b),
    .io_ci(FullAdder_3859_io_ci),
    .io_s(FullAdder_3859_io_s),
    .io_co(FullAdder_3859_io_co)
  );
  FullAdder FullAdder_3860 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3860_io_a),
    .io_b(FullAdder_3860_io_b),
    .io_ci(FullAdder_3860_io_ci),
    .io_s(FullAdder_3860_io_s),
    .io_co(FullAdder_3860_io_co)
  );
  FullAdder FullAdder_3861 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3861_io_a),
    .io_b(FullAdder_3861_io_b),
    .io_ci(FullAdder_3861_io_ci),
    .io_s(FullAdder_3861_io_s),
    .io_co(FullAdder_3861_io_co)
  );
  FullAdder FullAdder_3862 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3862_io_a),
    .io_b(FullAdder_3862_io_b),
    .io_ci(FullAdder_3862_io_ci),
    .io_s(FullAdder_3862_io_s),
    .io_co(FullAdder_3862_io_co)
  );
  HalfAdder HalfAdder_262 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_262_io_a),
    .io_b(HalfAdder_262_io_b),
    .io_s(HalfAdder_262_io_s),
    .io_co(HalfAdder_262_io_co)
  );
  FullAdder FullAdder_3863 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3863_io_a),
    .io_b(FullAdder_3863_io_b),
    .io_ci(FullAdder_3863_io_ci),
    .io_s(FullAdder_3863_io_s),
    .io_co(FullAdder_3863_io_co)
  );
  FullAdder FullAdder_3864 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3864_io_a),
    .io_b(FullAdder_3864_io_b),
    .io_ci(FullAdder_3864_io_ci),
    .io_s(FullAdder_3864_io_s),
    .io_co(FullAdder_3864_io_co)
  );
  FullAdder FullAdder_3865 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3865_io_a),
    .io_b(FullAdder_3865_io_b),
    .io_ci(FullAdder_3865_io_ci),
    .io_s(FullAdder_3865_io_s),
    .io_co(FullAdder_3865_io_co)
  );
  HalfAdder HalfAdder_263 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_263_io_a),
    .io_b(HalfAdder_263_io_b),
    .io_s(HalfAdder_263_io_s),
    .io_co(HalfAdder_263_io_co)
  );
  FullAdder FullAdder_3866 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3866_io_a),
    .io_b(FullAdder_3866_io_b),
    .io_ci(FullAdder_3866_io_ci),
    .io_s(FullAdder_3866_io_s),
    .io_co(FullAdder_3866_io_co)
  );
  FullAdder FullAdder_3867 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3867_io_a),
    .io_b(FullAdder_3867_io_b),
    .io_ci(FullAdder_3867_io_ci),
    .io_s(FullAdder_3867_io_s),
    .io_co(FullAdder_3867_io_co)
  );
  FullAdder FullAdder_3868 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3868_io_a),
    .io_b(FullAdder_3868_io_b),
    .io_ci(FullAdder_3868_io_ci),
    .io_s(FullAdder_3868_io_s),
    .io_co(FullAdder_3868_io_co)
  );
  HalfAdder HalfAdder_264 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_264_io_a),
    .io_b(HalfAdder_264_io_b),
    .io_s(HalfAdder_264_io_s),
    .io_co(HalfAdder_264_io_co)
  );
  HalfAdder HalfAdder_265 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_265_io_a),
    .io_b(HalfAdder_265_io_b),
    .io_s(HalfAdder_265_io_s),
    .io_co(HalfAdder_265_io_co)
  );
  HalfAdder HalfAdder_266 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_266_io_a),
    .io_b(HalfAdder_266_io_b),
    .io_s(HalfAdder_266_io_s),
    .io_co(HalfAdder_266_io_co)
  );
  FullAdder FullAdder_3869 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3869_io_a),
    .io_b(FullAdder_3869_io_b),
    .io_ci(FullAdder_3869_io_ci),
    .io_s(FullAdder_3869_io_s),
    .io_co(FullAdder_3869_io_co)
  );
  FullAdder FullAdder_3870 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3870_io_a),
    .io_b(FullAdder_3870_io_b),
    .io_ci(FullAdder_3870_io_ci),
    .io_s(FullAdder_3870_io_s),
    .io_co(FullAdder_3870_io_co)
  );
  FullAdder FullAdder_3871 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3871_io_a),
    .io_b(FullAdder_3871_io_b),
    .io_ci(FullAdder_3871_io_ci),
    .io_s(FullAdder_3871_io_s),
    .io_co(FullAdder_3871_io_co)
  );
  HalfAdder HalfAdder_267 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_267_io_a),
    .io_b(HalfAdder_267_io_b),
    .io_s(HalfAdder_267_io_s),
    .io_co(HalfAdder_267_io_co)
  );
  FullAdder FullAdder_3872 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3872_io_a),
    .io_b(FullAdder_3872_io_b),
    .io_ci(FullAdder_3872_io_ci),
    .io_s(FullAdder_3872_io_s),
    .io_co(FullAdder_3872_io_co)
  );
  FullAdder FullAdder_3873 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3873_io_a),
    .io_b(FullAdder_3873_io_b),
    .io_ci(FullAdder_3873_io_ci),
    .io_s(FullAdder_3873_io_s),
    .io_co(FullAdder_3873_io_co)
  );
  HalfAdder HalfAdder_268 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_268_io_a),
    .io_b(HalfAdder_268_io_b),
    .io_s(HalfAdder_268_io_s),
    .io_co(HalfAdder_268_io_co)
  );
  HalfAdder HalfAdder_269 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_269_io_a),
    .io_b(HalfAdder_269_io_b),
    .io_s(HalfAdder_269_io_s),
    .io_co(HalfAdder_269_io_co)
  );
  FullAdder FullAdder_3874 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3874_io_a),
    .io_b(FullAdder_3874_io_b),
    .io_ci(FullAdder_3874_io_ci),
    .io_s(FullAdder_3874_io_s),
    .io_co(FullAdder_3874_io_co)
  );
  FullAdder FullAdder_3875 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3875_io_a),
    .io_b(FullAdder_3875_io_b),
    .io_ci(FullAdder_3875_io_ci),
    .io_s(FullAdder_3875_io_s),
    .io_co(FullAdder_3875_io_co)
  );
  FullAdder FullAdder_3876 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3876_io_a),
    .io_b(FullAdder_3876_io_b),
    .io_ci(FullAdder_3876_io_ci),
    .io_s(FullAdder_3876_io_s),
    .io_co(FullAdder_3876_io_co)
  );
  HalfAdder HalfAdder_270 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_270_io_a),
    .io_b(HalfAdder_270_io_b),
    .io_s(HalfAdder_270_io_s),
    .io_co(HalfAdder_270_io_co)
  );
  FullAdder FullAdder_3877 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3877_io_a),
    .io_b(FullAdder_3877_io_b),
    .io_ci(FullAdder_3877_io_ci),
    .io_s(FullAdder_3877_io_s),
    .io_co(FullAdder_3877_io_co)
  );
  HalfAdder HalfAdder_271 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_271_io_a),
    .io_b(HalfAdder_271_io_b),
    .io_s(HalfAdder_271_io_s),
    .io_co(HalfAdder_271_io_co)
  );
  FullAdder FullAdder_3878 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3878_io_a),
    .io_b(FullAdder_3878_io_b),
    .io_ci(FullAdder_3878_io_ci),
    .io_s(FullAdder_3878_io_s),
    .io_co(FullAdder_3878_io_co)
  );
  FullAdder FullAdder_3879 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3879_io_a),
    .io_b(FullAdder_3879_io_b),
    .io_ci(FullAdder_3879_io_ci),
    .io_s(FullAdder_3879_io_s),
    .io_co(FullAdder_3879_io_co)
  );
  HalfAdder HalfAdder_272 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_272_io_a),
    .io_b(HalfAdder_272_io_b),
    .io_s(HalfAdder_272_io_s),
    .io_co(HalfAdder_272_io_co)
  );
  FullAdder FullAdder_3880 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3880_io_a),
    .io_b(FullAdder_3880_io_b),
    .io_ci(FullAdder_3880_io_ci),
    .io_s(FullAdder_3880_io_s),
    .io_co(FullAdder_3880_io_co)
  );
  FullAdder FullAdder_3881 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3881_io_a),
    .io_b(FullAdder_3881_io_b),
    .io_ci(FullAdder_3881_io_ci),
    .io_s(FullAdder_3881_io_s),
    .io_co(FullAdder_3881_io_co)
  );
  FullAdder FullAdder_3882 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3882_io_a),
    .io_b(FullAdder_3882_io_b),
    .io_ci(FullAdder_3882_io_ci),
    .io_s(FullAdder_3882_io_s),
    .io_co(FullAdder_3882_io_co)
  );
  HalfAdder HalfAdder_273 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_273_io_a),
    .io_b(HalfAdder_273_io_b),
    .io_s(HalfAdder_273_io_s),
    .io_co(HalfAdder_273_io_co)
  );
  FullAdder FullAdder_3883 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3883_io_a),
    .io_b(FullAdder_3883_io_b),
    .io_ci(FullAdder_3883_io_ci),
    .io_s(FullAdder_3883_io_s),
    .io_co(FullAdder_3883_io_co)
  );
  FullAdder FullAdder_3884 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3884_io_a),
    .io_b(FullAdder_3884_io_b),
    .io_ci(FullAdder_3884_io_ci),
    .io_s(FullAdder_3884_io_s),
    .io_co(FullAdder_3884_io_co)
  );
  FullAdder FullAdder_3885 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3885_io_a),
    .io_b(FullAdder_3885_io_b),
    .io_ci(FullAdder_3885_io_ci),
    .io_s(FullAdder_3885_io_s),
    .io_co(FullAdder_3885_io_co)
  );
  FullAdder FullAdder_3886 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3886_io_a),
    .io_b(FullAdder_3886_io_b),
    .io_ci(FullAdder_3886_io_ci),
    .io_s(FullAdder_3886_io_s),
    .io_co(FullAdder_3886_io_co)
  );
  FullAdder FullAdder_3887 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3887_io_a),
    .io_b(FullAdder_3887_io_b),
    .io_ci(FullAdder_3887_io_ci),
    .io_s(FullAdder_3887_io_s),
    .io_co(FullAdder_3887_io_co)
  );
  FullAdder FullAdder_3888 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3888_io_a),
    .io_b(FullAdder_3888_io_b),
    .io_ci(FullAdder_3888_io_ci),
    .io_s(FullAdder_3888_io_s),
    .io_co(FullAdder_3888_io_co)
  );
  HalfAdder HalfAdder_274 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_274_io_a),
    .io_b(HalfAdder_274_io_b),
    .io_s(HalfAdder_274_io_s),
    .io_co(HalfAdder_274_io_co)
  );
  HalfAdder HalfAdder_275 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_275_io_a),
    .io_b(HalfAdder_275_io_b),
    .io_s(HalfAdder_275_io_s),
    .io_co(HalfAdder_275_io_co)
  );
  FullAdder FullAdder_3889 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3889_io_a),
    .io_b(FullAdder_3889_io_b),
    .io_ci(FullAdder_3889_io_ci),
    .io_s(FullAdder_3889_io_s),
    .io_co(FullAdder_3889_io_co)
  );
  FullAdder FullAdder_3890 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3890_io_a),
    .io_b(FullAdder_3890_io_b),
    .io_ci(FullAdder_3890_io_ci),
    .io_s(FullAdder_3890_io_s),
    .io_co(FullAdder_3890_io_co)
  );
  FullAdder FullAdder_3891 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3891_io_a),
    .io_b(FullAdder_3891_io_b),
    .io_ci(FullAdder_3891_io_ci),
    .io_s(FullAdder_3891_io_s),
    .io_co(FullAdder_3891_io_co)
  );
  HalfAdder HalfAdder_276 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_276_io_a),
    .io_b(HalfAdder_276_io_b),
    .io_s(HalfAdder_276_io_s),
    .io_co(HalfAdder_276_io_co)
  );
  FullAdder FullAdder_3892 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3892_io_a),
    .io_b(FullAdder_3892_io_b),
    .io_ci(FullAdder_3892_io_ci),
    .io_s(FullAdder_3892_io_s),
    .io_co(FullAdder_3892_io_co)
  );
  HalfAdder HalfAdder_277 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_277_io_a),
    .io_b(HalfAdder_277_io_b),
    .io_s(HalfAdder_277_io_s),
    .io_co(HalfAdder_277_io_co)
  );
  HalfAdder HalfAdder_278 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_278_io_a),
    .io_b(HalfAdder_278_io_b),
    .io_s(HalfAdder_278_io_s),
    .io_co(HalfAdder_278_io_co)
  );
  HalfAdder HalfAdder_279 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_279_io_a),
    .io_b(HalfAdder_279_io_b),
    .io_s(HalfAdder_279_io_s),
    .io_co(HalfAdder_279_io_co)
  );
  HalfAdder HalfAdder_280 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_280_io_a),
    .io_b(HalfAdder_280_io_b),
    .io_s(HalfAdder_280_io_s),
    .io_co(HalfAdder_280_io_co)
  );
  FullAdder FullAdder_3893 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3893_io_a),
    .io_b(FullAdder_3893_io_b),
    .io_ci(FullAdder_3893_io_ci),
    .io_s(FullAdder_3893_io_s),
    .io_co(FullAdder_3893_io_co)
  );
  FullAdder FullAdder_3894 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3894_io_a),
    .io_b(FullAdder_3894_io_b),
    .io_ci(FullAdder_3894_io_ci),
    .io_s(FullAdder_3894_io_s),
    .io_co(FullAdder_3894_io_co)
  );
  HalfAdder HalfAdder_281 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_281_io_a),
    .io_b(HalfAdder_281_io_b),
    .io_s(HalfAdder_281_io_s),
    .io_co(HalfAdder_281_io_co)
  );
  FullAdder FullAdder_3895 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3895_io_a),
    .io_b(FullAdder_3895_io_b),
    .io_ci(FullAdder_3895_io_ci),
    .io_s(FullAdder_3895_io_s),
    .io_co(FullAdder_3895_io_co)
  );
  FullAdder FullAdder_3896 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3896_io_a),
    .io_b(FullAdder_3896_io_b),
    .io_ci(FullAdder_3896_io_ci),
    .io_s(FullAdder_3896_io_s),
    .io_co(FullAdder_3896_io_co)
  );
  HalfAdder HalfAdder_282 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_282_io_a),
    .io_b(HalfAdder_282_io_b),
    .io_s(HalfAdder_282_io_s),
    .io_co(HalfAdder_282_io_co)
  );
  FullAdder FullAdder_3897 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3897_io_a),
    .io_b(FullAdder_3897_io_b),
    .io_ci(FullAdder_3897_io_ci),
    .io_s(FullAdder_3897_io_s),
    .io_co(FullAdder_3897_io_co)
  );
  FullAdder FullAdder_3898 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3898_io_a),
    .io_b(FullAdder_3898_io_b),
    .io_ci(FullAdder_3898_io_ci),
    .io_s(FullAdder_3898_io_s),
    .io_co(FullAdder_3898_io_co)
  );
  HalfAdder HalfAdder_283 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_283_io_a),
    .io_b(HalfAdder_283_io_b),
    .io_s(HalfAdder_283_io_s),
    .io_co(HalfAdder_283_io_co)
  );
  FullAdder FullAdder_3899 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3899_io_a),
    .io_b(FullAdder_3899_io_b),
    .io_ci(FullAdder_3899_io_ci),
    .io_s(FullAdder_3899_io_s),
    .io_co(FullAdder_3899_io_co)
  );
  HalfAdder HalfAdder_284 ( // @[wallace.scala 57:25]
    .io_a(HalfAdder_284_io_a),
    .io_b(HalfAdder_284_io_b),
    .io_s(HalfAdder_284_io_s),
    .io_co(HalfAdder_284_io_co)
  );
  FullAdder FullAdder_3900 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3900_io_a),
    .io_b(FullAdder_3900_io_b),
    .io_ci(FullAdder_3900_io_ci),
    .io_s(FullAdder_3900_io_s),
    .io_co(FullAdder_3900_io_co)
  );
  FullAdder FullAdder_3901 ( // @[wallace.scala 67:25]
    .io_a(FullAdder_3901_io_a),
    .io_b(FullAdder_3901_io_b),
    .io_ci(FullAdder_3901_io_ci),
    .io_s(FullAdder_3901_io_s),
    .io_co(FullAdder_3901_io_co)
  );
  assign io_augend = {{1'd0}, _T_4221}; // @[wallace.scala 90:13]
  assign io_addend = {{1'd0}, _T_4347}; // @[wallace.scala 91:13]
  assign HalfAdder_io_a = io_pp_62[63]; // @[wallace.scala 59:18]
  assign HalfAdder_io_b = io_pp_63[62]; // @[wallace.scala 60:18]
  assign FullAdder_io_a = io_pp_61[63]; // @[wallace.scala 69:18]
  assign FullAdder_io_b = io_pp_62[62]; // @[wallace.scala 70:18]
  assign FullAdder_io_ci = io_pp_63[61]; // @[wallace.scala 71:19]
  assign FullAdder_1_io_a = io_pp_60[63]; // @[wallace.scala 69:18]
  assign FullAdder_1_io_b = io_pp_61[62]; // @[wallace.scala 70:18]
  assign FullAdder_1_io_ci = io_pp_62[61]; // @[wallace.scala 71:19]
  assign FullAdder_2_io_a = io_pp_59[63]; // @[wallace.scala 69:18]
  assign FullAdder_2_io_b = io_pp_60[62]; // @[wallace.scala 70:18]
  assign FullAdder_2_io_ci = io_pp_61[61]; // @[wallace.scala 71:19]
  assign HalfAdder_1_io_a = io_pp_62[60]; // @[wallace.scala 59:18]
  assign HalfAdder_1_io_b = io_pp_63[59]; // @[wallace.scala 60:18]
  assign FullAdder_3_io_a = io_pp_58[63]; // @[wallace.scala 69:18]
  assign FullAdder_3_io_b = io_pp_59[62]; // @[wallace.scala 70:18]
  assign FullAdder_3_io_ci = io_pp_60[61]; // @[wallace.scala 71:19]
  assign FullAdder_4_io_a = io_pp_61[60]; // @[wallace.scala 69:18]
  assign FullAdder_4_io_b = io_pp_62[59]; // @[wallace.scala 70:18]
  assign FullAdder_4_io_ci = io_pp_63[58]; // @[wallace.scala 71:19]
  assign FullAdder_5_io_a = io_pp_57[63]; // @[wallace.scala 69:18]
  assign FullAdder_5_io_b = io_pp_58[62]; // @[wallace.scala 70:18]
  assign FullAdder_5_io_ci = io_pp_59[61]; // @[wallace.scala 71:19]
  assign FullAdder_6_io_a = io_pp_60[60]; // @[wallace.scala 69:18]
  assign FullAdder_6_io_b = io_pp_61[59]; // @[wallace.scala 70:18]
  assign FullAdder_6_io_ci = io_pp_62[58]; // @[wallace.scala 71:19]
  assign FullAdder_7_io_a = io_pp_56[63]; // @[wallace.scala 69:18]
  assign FullAdder_7_io_b = io_pp_57[62]; // @[wallace.scala 70:18]
  assign FullAdder_7_io_ci = io_pp_58[61]; // @[wallace.scala 71:19]
  assign FullAdder_8_io_a = io_pp_59[60]; // @[wallace.scala 69:18]
  assign FullAdder_8_io_b = io_pp_60[59]; // @[wallace.scala 70:18]
  assign FullAdder_8_io_ci = io_pp_61[58]; // @[wallace.scala 71:19]
  assign HalfAdder_2_io_a = io_pp_62[57]; // @[wallace.scala 59:18]
  assign HalfAdder_2_io_b = io_pp_63[56]; // @[wallace.scala 60:18]
  assign FullAdder_9_io_a = io_pp_55[63]; // @[wallace.scala 69:18]
  assign FullAdder_9_io_b = io_pp_56[62]; // @[wallace.scala 70:18]
  assign FullAdder_9_io_ci = io_pp_57[61]; // @[wallace.scala 71:19]
  assign FullAdder_10_io_a = io_pp_58[60]; // @[wallace.scala 69:18]
  assign FullAdder_10_io_b = io_pp_59[59]; // @[wallace.scala 70:18]
  assign FullAdder_10_io_ci = io_pp_60[58]; // @[wallace.scala 71:19]
  assign FullAdder_11_io_a = io_pp_61[57]; // @[wallace.scala 69:18]
  assign FullAdder_11_io_b = io_pp_62[56]; // @[wallace.scala 70:18]
  assign FullAdder_11_io_ci = io_pp_63[55]; // @[wallace.scala 71:19]
  assign FullAdder_12_io_a = io_pp_54[63]; // @[wallace.scala 69:18]
  assign FullAdder_12_io_b = io_pp_55[62]; // @[wallace.scala 70:18]
  assign FullAdder_12_io_ci = io_pp_56[61]; // @[wallace.scala 71:19]
  assign FullAdder_13_io_a = io_pp_57[60]; // @[wallace.scala 69:18]
  assign FullAdder_13_io_b = io_pp_58[59]; // @[wallace.scala 70:18]
  assign FullAdder_13_io_ci = io_pp_59[58]; // @[wallace.scala 71:19]
  assign FullAdder_14_io_a = io_pp_60[57]; // @[wallace.scala 69:18]
  assign FullAdder_14_io_b = io_pp_61[56]; // @[wallace.scala 70:18]
  assign FullAdder_14_io_ci = io_pp_62[55]; // @[wallace.scala 71:19]
  assign FullAdder_15_io_a = io_pp_53[63]; // @[wallace.scala 69:18]
  assign FullAdder_15_io_b = io_pp_54[62]; // @[wallace.scala 70:18]
  assign FullAdder_15_io_ci = io_pp_55[61]; // @[wallace.scala 71:19]
  assign FullAdder_16_io_a = io_pp_56[60]; // @[wallace.scala 69:18]
  assign FullAdder_16_io_b = io_pp_57[59]; // @[wallace.scala 70:18]
  assign FullAdder_16_io_ci = io_pp_58[58]; // @[wallace.scala 71:19]
  assign FullAdder_17_io_a = io_pp_59[57]; // @[wallace.scala 69:18]
  assign FullAdder_17_io_b = io_pp_60[56]; // @[wallace.scala 70:18]
  assign FullAdder_17_io_ci = io_pp_61[55]; // @[wallace.scala 71:19]
  assign HalfAdder_3_io_a = io_pp_62[54]; // @[wallace.scala 59:18]
  assign HalfAdder_3_io_b = io_pp_63[53]; // @[wallace.scala 60:18]
  assign FullAdder_18_io_a = io_pp_52[63]; // @[wallace.scala 69:18]
  assign FullAdder_18_io_b = io_pp_53[62]; // @[wallace.scala 70:18]
  assign FullAdder_18_io_ci = io_pp_54[61]; // @[wallace.scala 71:19]
  assign FullAdder_19_io_a = io_pp_55[60]; // @[wallace.scala 69:18]
  assign FullAdder_19_io_b = io_pp_56[59]; // @[wallace.scala 70:18]
  assign FullAdder_19_io_ci = io_pp_57[58]; // @[wallace.scala 71:19]
  assign FullAdder_20_io_a = io_pp_58[57]; // @[wallace.scala 69:18]
  assign FullAdder_20_io_b = io_pp_59[56]; // @[wallace.scala 70:18]
  assign FullAdder_20_io_ci = io_pp_60[55]; // @[wallace.scala 71:19]
  assign FullAdder_21_io_a = io_pp_61[54]; // @[wallace.scala 69:18]
  assign FullAdder_21_io_b = io_pp_62[53]; // @[wallace.scala 70:18]
  assign FullAdder_21_io_ci = io_pp_63[52]; // @[wallace.scala 71:19]
  assign FullAdder_22_io_a = io_pp_51[63]; // @[wallace.scala 69:18]
  assign FullAdder_22_io_b = io_pp_52[62]; // @[wallace.scala 70:18]
  assign FullAdder_22_io_ci = io_pp_53[61]; // @[wallace.scala 71:19]
  assign FullAdder_23_io_a = io_pp_54[60]; // @[wallace.scala 69:18]
  assign FullAdder_23_io_b = io_pp_55[59]; // @[wallace.scala 70:18]
  assign FullAdder_23_io_ci = io_pp_56[58]; // @[wallace.scala 71:19]
  assign FullAdder_24_io_a = io_pp_57[57]; // @[wallace.scala 69:18]
  assign FullAdder_24_io_b = io_pp_58[56]; // @[wallace.scala 70:18]
  assign FullAdder_24_io_ci = io_pp_59[55]; // @[wallace.scala 71:19]
  assign FullAdder_25_io_a = io_pp_60[54]; // @[wallace.scala 69:18]
  assign FullAdder_25_io_b = io_pp_61[53]; // @[wallace.scala 70:18]
  assign FullAdder_25_io_ci = io_pp_62[52]; // @[wallace.scala 71:19]
  assign FullAdder_26_io_a = io_pp_50[63]; // @[wallace.scala 69:18]
  assign FullAdder_26_io_b = io_pp_51[62]; // @[wallace.scala 70:18]
  assign FullAdder_26_io_ci = io_pp_52[61]; // @[wallace.scala 71:19]
  assign FullAdder_27_io_a = io_pp_53[60]; // @[wallace.scala 69:18]
  assign FullAdder_27_io_b = io_pp_54[59]; // @[wallace.scala 70:18]
  assign FullAdder_27_io_ci = io_pp_55[58]; // @[wallace.scala 71:19]
  assign FullAdder_28_io_a = io_pp_56[57]; // @[wallace.scala 69:18]
  assign FullAdder_28_io_b = io_pp_57[56]; // @[wallace.scala 70:18]
  assign FullAdder_28_io_ci = io_pp_58[55]; // @[wallace.scala 71:19]
  assign FullAdder_29_io_a = io_pp_59[54]; // @[wallace.scala 69:18]
  assign FullAdder_29_io_b = io_pp_60[53]; // @[wallace.scala 70:18]
  assign FullAdder_29_io_ci = io_pp_61[52]; // @[wallace.scala 71:19]
  assign FullAdder_30_io_a = io_pp_49[63]; // @[wallace.scala 69:18]
  assign FullAdder_30_io_b = io_pp_50[62]; // @[wallace.scala 70:18]
  assign FullAdder_30_io_ci = io_pp_51[61]; // @[wallace.scala 71:19]
  assign FullAdder_31_io_a = io_pp_52[60]; // @[wallace.scala 69:18]
  assign FullAdder_31_io_b = io_pp_53[59]; // @[wallace.scala 70:18]
  assign FullAdder_31_io_ci = io_pp_54[58]; // @[wallace.scala 71:19]
  assign FullAdder_32_io_a = io_pp_55[57]; // @[wallace.scala 69:18]
  assign FullAdder_32_io_b = io_pp_56[56]; // @[wallace.scala 70:18]
  assign FullAdder_32_io_ci = io_pp_57[55]; // @[wallace.scala 71:19]
  assign FullAdder_33_io_a = io_pp_58[54]; // @[wallace.scala 69:18]
  assign FullAdder_33_io_b = io_pp_59[53]; // @[wallace.scala 70:18]
  assign FullAdder_33_io_ci = io_pp_60[52]; // @[wallace.scala 71:19]
  assign FullAdder_34_io_a = io_pp_61[51]; // @[wallace.scala 69:18]
  assign FullAdder_34_io_b = io_pp_62[50]; // @[wallace.scala 70:18]
  assign FullAdder_34_io_ci = io_pp_63[49]; // @[wallace.scala 71:19]
  assign FullAdder_35_io_a = io_pp_48[63]; // @[wallace.scala 69:18]
  assign FullAdder_35_io_b = io_pp_49[62]; // @[wallace.scala 70:18]
  assign FullAdder_35_io_ci = io_pp_50[61]; // @[wallace.scala 71:19]
  assign FullAdder_36_io_a = io_pp_51[60]; // @[wallace.scala 69:18]
  assign FullAdder_36_io_b = io_pp_52[59]; // @[wallace.scala 70:18]
  assign FullAdder_36_io_ci = io_pp_53[58]; // @[wallace.scala 71:19]
  assign FullAdder_37_io_a = io_pp_54[57]; // @[wallace.scala 69:18]
  assign FullAdder_37_io_b = io_pp_55[56]; // @[wallace.scala 70:18]
  assign FullAdder_37_io_ci = io_pp_56[55]; // @[wallace.scala 71:19]
  assign FullAdder_38_io_a = io_pp_57[54]; // @[wallace.scala 69:18]
  assign FullAdder_38_io_b = io_pp_58[53]; // @[wallace.scala 70:18]
  assign FullAdder_38_io_ci = io_pp_59[52]; // @[wallace.scala 71:19]
  assign FullAdder_39_io_a = io_pp_60[51]; // @[wallace.scala 69:18]
  assign FullAdder_39_io_b = io_pp_61[50]; // @[wallace.scala 70:18]
  assign FullAdder_39_io_ci = io_pp_62[49]; // @[wallace.scala 71:19]
  assign FullAdder_40_io_a = io_pp_47[63]; // @[wallace.scala 69:18]
  assign FullAdder_40_io_b = io_pp_48[62]; // @[wallace.scala 70:18]
  assign FullAdder_40_io_ci = io_pp_49[61]; // @[wallace.scala 71:19]
  assign FullAdder_41_io_a = io_pp_50[60]; // @[wallace.scala 69:18]
  assign FullAdder_41_io_b = io_pp_51[59]; // @[wallace.scala 70:18]
  assign FullAdder_41_io_ci = io_pp_52[58]; // @[wallace.scala 71:19]
  assign FullAdder_42_io_a = io_pp_53[57]; // @[wallace.scala 69:18]
  assign FullAdder_42_io_b = io_pp_54[56]; // @[wallace.scala 70:18]
  assign FullAdder_42_io_ci = io_pp_55[55]; // @[wallace.scala 71:19]
  assign FullAdder_43_io_a = io_pp_56[54]; // @[wallace.scala 69:18]
  assign FullAdder_43_io_b = io_pp_57[53]; // @[wallace.scala 70:18]
  assign FullAdder_43_io_ci = io_pp_58[52]; // @[wallace.scala 71:19]
  assign FullAdder_44_io_a = io_pp_59[51]; // @[wallace.scala 69:18]
  assign FullAdder_44_io_b = io_pp_60[50]; // @[wallace.scala 70:18]
  assign FullAdder_44_io_ci = io_pp_61[49]; // @[wallace.scala 71:19]
  assign HalfAdder_4_io_a = io_pp_62[48]; // @[wallace.scala 59:18]
  assign HalfAdder_4_io_b = io_pp_63[47]; // @[wallace.scala 60:18]
  assign FullAdder_45_io_a = io_pp_46[63]; // @[wallace.scala 69:18]
  assign FullAdder_45_io_b = io_pp_47[62]; // @[wallace.scala 70:18]
  assign FullAdder_45_io_ci = io_pp_48[61]; // @[wallace.scala 71:19]
  assign FullAdder_46_io_a = io_pp_49[60]; // @[wallace.scala 69:18]
  assign FullAdder_46_io_b = io_pp_50[59]; // @[wallace.scala 70:18]
  assign FullAdder_46_io_ci = io_pp_51[58]; // @[wallace.scala 71:19]
  assign FullAdder_47_io_a = io_pp_52[57]; // @[wallace.scala 69:18]
  assign FullAdder_47_io_b = io_pp_53[56]; // @[wallace.scala 70:18]
  assign FullAdder_47_io_ci = io_pp_54[55]; // @[wallace.scala 71:19]
  assign FullAdder_48_io_a = io_pp_55[54]; // @[wallace.scala 69:18]
  assign FullAdder_48_io_b = io_pp_56[53]; // @[wallace.scala 70:18]
  assign FullAdder_48_io_ci = io_pp_57[52]; // @[wallace.scala 71:19]
  assign FullAdder_49_io_a = io_pp_58[51]; // @[wallace.scala 69:18]
  assign FullAdder_49_io_b = io_pp_59[50]; // @[wallace.scala 70:18]
  assign FullAdder_49_io_ci = io_pp_60[49]; // @[wallace.scala 71:19]
  assign FullAdder_50_io_a = io_pp_61[48]; // @[wallace.scala 69:18]
  assign FullAdder_50_io_b = io_pp_62[47]; // @[wallace.scala 70:18]
  assign FullAdder_50_io_ci = io_pp_63[46]; // @[wallace.scala 71:19]
  assign FullAdder_51_io_a = io_pp_45[63]; // @[wallace.scala 69:18]
  assign FullAdder_51_io_b = io_pp_46[62]; // @[wallace.scala 70:18]
  assign FullAdder_51_io_ci = io_pp_47[61]; // @[wallace.scala 71:19]
  assign FullAdder_52_io_a = io_pp_48[60]; // @[wallace.scala 69:18]
  assign FullAdder_52_io_b = io_pp_49[59]; // @[wallace.scala 70:18]
  assign FullAdder_52_io_ci = io_pp_50[58]; // @[wallace.scala 71:19]
  assign FullAdder_53_io_a = io_pp_51[57]; // @[wallace.scala 69:18]
  assign FullAdder_53_io_b = io_pp_52[56]; // @[wallace.scala 70:18]
  assign FullAdder_53_io_ci = io_pp_53[55]; // @[wallace.scala 71:19]
  assign FullAdder_54_io_a = io_pp_54[54]; // @[wallace.scala 69:18]
  assign FullAdder_54_io_b = io_pp_55[53]; // @[wallace.scala 70:18]
  assign FullAdder_54_io_ci = io_pp_56[52]; // @[wallace.scala 71:19]
  assign FullAdder_55_io_a = io_pp_57[51]; // @[wallace.scala 69:18]
  assign FullAdder_55_io_b = io_pp_58[50]; // @[wallace.scala 70:18]
  assign FullAdder_55_io_ci = io_pp_59[49]; // @[wallace.scala 71:19]
  assign FullAdder_56_io_a = io_pp_60[48]; // @[wallace.scala 69:18]
  assign FullAdder_56_io_b = io_pp_61[47]; // @[wallace.scala 70:18]
  assign FullAdder_56_io_ci = io_pp_62[46]; // @[wallace.scala 71:19]
  assign FullAdder_57_io_a = io_pp_44[63]; // @[wallace.scala 69:18]
  assign FullAdder_57_io_b = io_pp_45[62]; // @[wallace.scala 70:18]
  assign FullAdder_57_io_ci = io_pp_46[61]; // @[wallace.scala 71:19]
  assign FullAdder_58_io_a = io_pp_47[60]; // @[wallace.scala 69:18]
  assign FullAdder_58_io_b = io_pp_48[59]; // @[wallace.scala 70:18]
  assign FullAdder_58_io_ci = io_pp_49[58]; // @[wallace.scala 71:19]
  assign FullAdder_59_io_a = io_pp_50[57]; // @[wallace.scala 69:18]
  assign FullAdder_59_io_b = io_pp_51[56]; // @[wallace.scala 70:18]
  assign FullAdder_59_io_ci = io_pp_52[55]; // @[wallace.scala 71:19]
  assign FullAdder_60_io_a = io_pp_53[54]; // @[wallace.scala 69:18]
  assign FullAdder_60_io_b = io_pp_54[53]; // @[wallace.scala 70:18]
  assign FullAdder_60_io_ci = io_pp_55[52]; // @[wallace.scala 71:19]
  assign FullAdder_61_io_a = io_pp_56[51]; // @[wallace.scala 69:18]
  assign FullAdder_61_io_b = io_pp_57[50]; // @[wallace.scala 70:18]
  assign FullAdder_61_io_ci = io_pp_58[49]; // @[wallace.scala 71:19]
  assign FullAdder_62_io_a = io_pp_59[48]; // @[wallace.scala 69:18]
  assign FullAdder_62_io_b = io_pp_60[47]; // @[wallace.scala 70:18]
  assign FullAdder_62_io_ci = io_pp_61[46]; // @[wallace.scala 71:19]
  assign HalfAdder_5_io_a = io_pp_62[45]; // @[wallace.scala 59:18]
  assign HalfAdder_5_io_b = io_pp_63[44]; // @[wallace.scala 60:18]
  assign FullAdder_63_io_a = io_pp_43[63]; // @[wallace.scala 69:18]
  assign FullAdder_63_io_b = io_pp_44[62]; // @[wallace.scala 70:18]
  assign FullAdder_63_io_ci = io_pp_45[61]; // @[wallace.scala 71:19]
  assign FullAdder_64_io_a = io_pp_46[60]; // @[wallace.scala 69:18]
  assign FullAdder_64_io_b = io_pp_47[59]; // @[wallace.scala 70:18]
  assign FullAdder_64_io_ci = io_pp_48[58]; // @[wallace.scala 71:19]
  assign FullAdder_65_io_a = io_pp_49[57]; // @[wallace.scala 69:18]
  assign FullAdder_65_io_b = io_pp_50[56]; // @[wallace.scala 70:18]
  assign FullAdder_65_io_ci = io_pp_51[55]; // @[wallace.scala 71:19]
  assign FullAdder_66_io_a = io_pp_52[54]; // @[wallace.scala 69:18]
  assign FullAdder_66_io_b = io_pp_53[53]; // @[wallace.scala 70:18]
  assign FullAdder_66_io_ci = io_pp_54[52]; // @[wallace.scala 71:19]
  assign FullAdder_67_io_a = io_pp_55[51]; // @[wallace.scala 69:18]
  assign FullAdder_67_io_b = io_pp_56[50]; // @[wallace.scala 70:18]
  assign FullAdder_67_io_ci = io_pp_57[49]; // @[wallace.scala 71:19]
  assign FullAdder_68_io_a = io_pp_58[48]; // @[wallace.scala 69:18]
  assign FullAdder_68_io_b = io_pp_59[47]; // @[wallace.scala 70:18]
  assign FullAdder_68_io_ci = io_pp_60[46]; // @[wallace.scala 71:19]
  assign FullAdder_69_io_a = io_pp_61[45]; // @[wallace.scala 69:18]
  assign FullAdder_69_io_b = io_pp_62[44]; // @[wallace.scala 70:18]
  assign FullAdder_69_io_ci = io_pp_63[43]; // @[wallace.scala 71:19]
  assign FullAdder_70_io_a = io_pp_42[63]; // @[wallace.scala 69:18]
  assign FullAdder_70_io_b = io_pp_43[62]; // @[wallace.scala 70:18]
  assign FullAdder_70_io_ci = io_pp_44[61]; // @[wallace.scala 71:19]
  assign FullAdder_71_io_a = io_pp_45[60]; // @[wallace.scala 69:18]
  assign FullAdder_71_io_b = io_pp_46[59]; // @[wallace.scala 70:18]
  assign FullAdder_71_io_ci = io_pp_47[58]; // @[wallace.scala 71:19]
  assign FullAdder_72_io_a = io_pp_48[57]; // @[wallace.scala 69:18]
  assign FullAdder_72_io_b = io_pp_49[56]; // @[wallace.scala 70:18]
  assign FullAdder_72_io_ci = io_pp_50[55]; // @[wallace.scala 71:19]
  assign FullAdder_73_io_a = io_pp_51[54]; // @[wallace.scala 69:18]
  assign FullAdder_73_io_b = io_pp_52[53]; // @[wallace.scala 70:18]
  assign FullAdder_73_io_ci = io_pp_53[52]; // @[wallace.scala 71:19]
  assign FullAdder_74_io_a = io_pp_54[51]; // @[wallace.scala 69:18]
  assign FullAdder_74_io_b = io_pp_55[50]; // @[wallace.scala 70:18]
  assign FullAdder_74_io_ci = io_pp_56[49]; // @[wallace.scala 71:19]
  assign FullAdder_75_io_a = io_pp_57[48]; // @[wallace.scala 69:18]
  assign FullAdder_75_io_b = io_pp_58[47]; // @[wallace.scala 70:18]
  assign FullAdder_75_io_ci = io_pp_59[46]; // @[wallace.scala 71:19]
  assign FullAdder_76_io_a = io_pp_60[45]; // @[wallace.scala 69:18]
  assign FullAdder_76_io_b = io_pp_61[44]; // @[wallace.scala 70:18]
  assign FullAdder_76_io_ci = io_pp_62[43]; // @[wallace.scala 71:19]
  assign FullAdder_77_io_a = io_pp_41[63]; // @[wallace.scala 69:18]
  assign FullAdder_77_io_b = io_pp_42[62]; // @[wallace.scala 70:18]
  assign FullAdder_77_io_ci = io_pp_43[61]; // @[wallace.scala 71:19]
  assign FullAdder_78_io_a = io_pp_44[60]; // @[wallace.scala 69:18]
  assign FullAdder_78_io_b = io_pp_45[59]; // @[wallace.scala 70:18]
  assign FullAdder_78_io_ci = io_pp_46[58]; // @[wallace.scala 71:19]
  assign FullAdder_79_io_a = io_pp_47[57]; // @[wallace.scala 69:18]
  assign FullAdder_79_io_b = io_pp_48[56]; // @[wallace.scala 70:18]
  assign FullAdder_79_io_ci = io_pp_49[55]; // @[wallace.scala 71:19]
  assign FullAdder_80_io_a = io_pp_50[54]; // @[wallace.scala 69:18]
  assign FullAdder_80_io_b = io_pp_51[53]; // @[wallace.scala 70:18]
  assign FullAdder_80_io_ci = io_pp_52[52]; // @[wallace.scala 71:19]
  assign FullAdder_81_io_a = io_pp_53[51]; // @[wallace.scala 69:18]
  assign FullAdder_81_io_b = io_pp_54[50]; // @[wallace.scala 70:18]
  assign FullAdder_81_io_ci = io_pp_55[49]; // @[wallace.scala 71:19]
  assign FullAdder_82_io_a = io_pp_56[48]; // @[wallace.scala 69:18]
  assign FullAdder_82_io_b = io_pp_57[47]; // @[wallace.scala 70:18]
  assign FullAdder_82_io_ci = io_pp_58[46]; // @[wallace.scala 71:19]
  assign FullAdder_83_io_a = io_pp_59[45]; // @[wallace.scala 69:18]
  assign FullAdder_83_io_b = io_pp_60[44]; // @[wallace.scala 70:18]
  assign FullAdder_83_io_ci = io_pp_61[43]; // @[wallace.scala 71:19]
  assign HalfAdder_6_io_a = io_pp_62[42]; // @[wallace.scala 59:18]
  assign HalfAdder_6_io_b = io_pp_63[41]; // @[wallace.scala 60:18]
  assign FullAdder_84_io_a = io_pp_40[63]; // @[wallace.scala 69:18]
  assign FullAdder_84_io_b = io_pp_41[62]; // @[wallace.scala 70:18]
  assign FullAdder_84_io_ci = io_pp_42[61]; // @[wallace.scala 71:19]
  assign FullAdder_85_io_a = io_pp_43[60]; // @[wallace.scala 69:18]
  assign FullAdder_85_io_b = io_pp_44[59]; // @[wallace.scala 70:18]
  assign FullAdder_85_io_ci = io_pp_45[58]; // @[wallace.scala 71:19]
  assign FullAdder_86_io_a = io_pp_46[57]; // @[wallace.scala 69:18]
  assign FullAdder_86_io_b = io_pp_47[56]; // @[wallace.scala 70:18]
  assign FullAdder_86_io_ci = io_pp_48[55]; // @[wallace.scala 71:19]
  assign FullAdder_87_io_a = io_pp_49[54]; // @[wallace.scala 69:18]
  assign FullAdder_87_io_b = io_pp_50[53]; // @[wallace.scala 70:18]
  assign FullAdder_87_io_ci = io_pp_51[52]; // @[wallace.scala 71:19]
  assign FullAdder_88_io_a = io_pp_52[51]; // @[wallace.scala 69:18]
  assign FullAdder_88_io_b = io_pp_53[50]; // @[wallace.scala 70:18]
  assign FullAdder_88_io_ci = io_pp_54[49]; // @[wallace.scala 71:19]
  assign FullAdder_89_io_a = io_pp_55[48]; // @[wallace.scala 69:18]
  assign FullAdder_89_io_b = io_pp_56[47]; // @[wallace.scala 70:18]
  assign FullAdder_89_io_ci = io_pp_57[46]; // @[wallace.scala 71:19]
  assign FullAdder_90_io_a = io_pp_58[45]; // @[wallace.scala 69:18]
  assign FullAdder_90_io_b = io_pp_59[44]; // @[wallace.scala 70:18]
  assign FullAdder_90_io_ci = io_pp_60[43]; // @[wallace.scala 71:19]
  assign FullAdder_91_io_a = io_pp_61[42]; // @[wallace.scala 69:18]
  assign FullAdder_91_io_b = io_pp_62[41]; // @[wallace.scala 70:18]
  assign FullAdder_91_io_ci = io_pp_63[40]; // @[wallace.scala 71:19]
  assign FullAdder_92_io_a = io_pp_39[63]; // @[wallace.scala 69:18]
  assign FullAdder_92_io_b = io_pp_40[62]; // @[wallace.scala 70:18]
  assign FullAdder_92_io_ci = io_pp_41[61]; // @[wallace.scala 71:19]
  assign FullAdder_93_io_a = io_pp_42[60]; // @[wallace.scala 69:18]
  assign FullAdder_93_io_b = io_pp_43[59]; // @[wallace.scala 70:18]
  assign FullAdder_93_io_ci = io_pp_44[58]; // @[wallace.scala 71:19]
  assign FullAdder_94_io_a = io_pp_45[57]; // @[wallace.scala 69:18]
  assign FullAdder_94_io_b = io_pp_46[56]; // @[wallace.scala 70:18]
  assign FullAdder_94_io_ci = io_pp_47[55]; // @[wallace.scala 71:19]
  assign FullAdder_95_io_a = io_pp_48[54]; // @[wallace.scala 69:18]
  assign FullAdder_95_io_b = io_pp_49[53]; // @[wallace.scala 70:18]
  assign FullAdder_95_io_ci = io_pp_50[52]; // @[wallace.scala 71:19]
  assign FullAdder_96_io_a = io_pp_51[51]; // @[wallace.scala 69:18]
  assign FullAdder_96_io_b = io_pp_52[50]; // @[wallace.scala 70:18]
  assign FullAdder_96_io_ci = io_pp_53[49]; // @[wallace.scala 71:19]
  assign FullAdder_97_io_a = io_pp_54[48]; // @[wallace.scala 69:18]
  assign FullAdder_97_io_b = io_pp_55[47]; // @[wallace.scala 70:18]
  assign FullAdder_97_io_ci = io_pp_56[46]; // @[wallace.scala 71:19]
  assign FullAdder_98_io_a = io_pp_57[45]; // @[wallace.scala 69:18]
  assign FullAdder_98_io_b = io_pp_58[44]; // @[wallace.scala 70:18]
  assign FullAdder_98_io_ci = io_pp_59[43]; // @[wallace.scala 71:19]
  assign FullAdder_99_io_a = io_pp_60[42]; // @[wallace.scala 69:18]
  assign FullAdder_99_io_b = io_pp_61[41]; // @[wallace.scala 70:18]
  assign FullAdder_99_io_ci = io_pp_62[40]; // @[wallace.scala 71:19]
  assign FullAdder_100_io_a = io_pp_38[63]; // @[wallace.scala 69:18]
  assign FullAdder_100_io_b = io_pp_39[62]; // @[wallace.scala 70:18]
  assign FullAdder_100_io_ci = io_pp_40[61]; // @[wallace.scala 71:19]
  assign FullAdder_101_io_a = io_pp_41[60]; // @[wallace.scala 69:18]
  assign FullAdder_101_io_b = io_pp_42[59]; // @[wallace.scala 70:18]
  assign FullAdder_101_io_ci = io_pp_43[58]; // @[wallace.scala 71:19]
  assign FullAdder_102_io_a = io_pp_44[57]; // @[wallace.scala 69:18]
  assign FullAdder_102_io_b = io_pp_45[56]; // @[wallace.scala 70:18]
  assign FullAdder_102_io_ci = io_pp_46[55]; // @[wallace.scala 71:19]
  assign FullAdder_103_io_a = io_pp_47[54]; // @[wallace.scala 69:18]
  assign FullAdder_103_io_b = io_pp_48[53]; // @[wallace.scala 70:18]
  assign FullAdder_103_io_ci = io_pp_49[52]; // @[wallace.scala 71:19]
  assign FullAdder_104_io_a = io_pp_50[51]; // @[wallace.scala 69:18]
  assign FullAdder_104_io_b = io_pp_51[50]; // @[wallace.scala 70:18]
  assign FullAdder_104_io_ci = io_pp_52[49]; // @[wallace.scala 71:19]
  assign FullAdder_105_io_a = io_pp_53[48]; // @[wallace.scala 69:18]
  assign FullAdder_105_io_b = io_pp_54[47]; // @[wallace.scala 70:18]
  assign FullAdder_105_io_ci = io_pp_55[46]; // @[wallace.scala 71:19]
  assign FullAdder_106_io_a = io_pp_56[45]; // @[wallace.scala 69:18]
  assign FullAdder_106_io_b = io_pp_57[44]; // @[wallace.scala 70:18]
  assign FullAdder_106_io_ci = io_pp_58[43]; // @[wallace.scala 71:19]
  assign FullAdder_107_io_a = io_pp_59[42]; // @[wallace.scala 69:18]
  assign FullAdder_107_io_b = io_pp_60[41]; // @[wallace.scala 70:18]
  assign FullAdder_107_io_ci = io_pp_61[40]; // @[wallace.scala 71:19]
  assign FullAdder_108_io_a = io_pp_37[63]; // @[wallace.scala 69:18]
  assign FullAdder_108_io_b = io_pp_38[62]; // @[wallace.scala 70:18]
  assign FullAdder_108_io_ci = io_pp_39[61]; // @[wallace.scala 71:19]
  assign FullAdder_109_io_a = io_pp_40[60]; // @[wallace.scala 69:18]
  assign FullAdder_109_io_b = io_pp_41[59]; // @[wallace.scala 70:18]
  assign FullAdder_109_io_ci = io_pp_42[58]; // @[wallace.scala 71:19]
  assign FullAdder_110_io_a = io_pp_43[57]; // @[wallace.scala 69:18]
  assign FullAdder_110_io_b = io_pp_44[56]; // @[wallace.scala 70:18]
  assign FullAdder_110_io_ci = io_pp_45[55]; // @[wallace.scala 71:19]
  assign FullAdder_111_io_a = io_pp_46[54]; // @[wallace.scala 69:18]
  assign FullAdder_111_io_b = io_pp_47[53]; // @[wallace.scala 70:18]
  assign FullAdder_111_io_ci = io_pp_48[52]; // @[wallace.scala 71:19]
  assign FullAdder_112_io_a = io_pp_49[51]; // @[wallace.scala 69:18]
  assign FullAdder_112_io_b = io_pp_50[50]; // @[wallace.scala 70:18]
  assign FullAdder_112_io_ci = io_pp_51[49]; // @[wallace.scala 71:19]
  assign FullAdder_113_io_a = io_pp_52[48]; // @[wallace.scala 69:18]
  assign FullAdder_113_io_b = io_pp_53[47]; // @[wallace.scala 70:18]
  assign FullAdder_113_io_ci = io_pp_54[46]; // @[wallace.scala 71:19]
  assign FullAdder_114_io_a = io_pp_55[45]; // @[wallace.scala 69:18]
  assign FullAdder_114_io_b = io_pp_56[44]; // @[wallace.scala 70:18]
  assign FullAdder_114_io_ci = io_pp_57[43]; // @[wallace.scala 71:19]
  assign FullAdder_115_io_a = io_pp_58[42]; // @[wallace.scala 69:18]
  assign FullAdder_115_io_b = io_pp_59[41]; // @[wallace.scala 70:18]
  assign FullAdder_115_io_ci = io_pp_60[40]; // @[wallace.scala 71:19]
  assign FullAdder_116_io_a = io_pp_61[39]; // @[wallace.scala 69:18]
  assign FullAdder_116_io_b = io_pp_62[38]; // @[wallace.scala 70:18]
  assign FullAdder_116_io_ci = io_pp_63[37]; // @[wallace.scala 71:19]
  assign FullAdder_117_io_a = io_pp_36[63]; // @[wallace.scala 69:18]
  assign FullAdder_117_io_b = io_pp_37[62]; // @[wallace.scala 70:18]
  assign FullAdder_117_io_ci = io_pp_38[61]; // @[wallace.scala 71:19]
  assign FullAdder_118_io_a = io_pp_39[60]; // @[wallace.scala 69:18]
  assign FullAdder_118_io_b = io_pp_40[59]; // @[wallace.scala 70:18]
  assign FullAdder_118_io_ci = io_pp_41[58]; // @[wallace.scala 71:19]
  assign FullAdder_119_io_a = io_pp_42[57]; // @[wallace.scala 69:18]
  assign FullAdder_119_io_b = io_pp_43[56]; // @[wallace.scala 70:18]
  assign FullAdder_119_io_ci = io_pp_44[55]; // @[wallace.scala 71:19]
  assign FullAdder_120_io_a = io_pp_45[54]; // @[wallace.scala 69:18]
  assign FullAdder_120_io_b = io_pp_46[53]; // @[wallace.scala 70:18]
  assign FullAdder_120_io_ci = io_pp_47[52]; // @[wallace.scala 71:19]
  assign FullAdder_121_io_a = io_pp_48[51]; // @[wallace.scala 69:18]
  assign FullAdder_121_io_b = io_pp_49[50]; // @[wallace.scala 70:18]
  assign FullAdder_121_io_ci = io_pp_50[49]; // @[wallace.scala 71:19]
  assign FullAdder_122_io_a = io_pp_51[48]; // @[wallace.scala 69:18]
  assign FullAdder_122_io_b = io_pp_52[47]; // @[wallace.scala 70:18]
  assign FullAdder_122_io_ci = io_pp_53[46]; // @[wallace.scala 71:19]
  assign FullAdder_123_io_a = io_pp_54[45]; // @[wallace.scala 69:18]
  assign FullAdder_123_io_b = io_pp_55[44]; // @[wallace.scala 70:18]
  assign FullAdder_123_io_ci = io_pp_56[43]; // @[wallace.scala 71:19]
  assign FullAdder_124_io_a = io_pp_57[42]; // @[wallace.scala 69:18]
  assign FullAdder_124_io_b = io_pp_58[41]; // @[wallace.scala 70:18]
  assign FullAdder_124_io_ci = io_pp_59[40]; // @[wallace.scala 71:19]
  assign FullAdder_125_io_a = io_pp_60[39]; // @[wallace.scala 69:18]
  assign FullAdder_125_io_b = io_pp_61[38]; // @[wallace.scala 70:18]
  assign FullAdder_125_io_ci = io_pp_62[37]; // @[wallace.scala 71:19]
  assign FullAdder_126_io_a = io_pp_35[63]; // @[wallace.scala 69:18]
  assign FullAdder_126_io_b = io_pp_36[62]; // @[wallace.scala 70:18]
  assign FullAdder_126_io_ci = io_pp_37[61]; // @[wallace.scala 71:19]
  assign FullAdder_127_io_a = io_pp_38[60]; // @[wallace.scala 69:18]
  assign FullAdder_127_io_b = io_pp_39[59]; // @[wallace.scala 70:18]
  assign FullAdder_127_io_ci = io_pp_40[58]; // @[wallace.scala 71:19]
  assign FullAdder_128_io_a = io_pp_41[57]; // @[wallace.scala 69:18]
  assign FullAdder_128_io_b = io_pp_42[56]; // @[wallace.scala 70:18]
  assign FullAdder_128_io_ci = io_pp_43[55]; // @[wallace.scala 71:19]
  assign FullAdder_129_io_a = io_pp_44[54]; // @[wallace.scala 69:18]
  assign FullAdder_129_io_b = io_pp_45[53]; // @[wallace.scala 70:18]
  assign FullAdder_129_io_ci = io_pp_46[52]; // @[wallace.scala 71:19]
  assign FullAdder_130_io_a = io_pp_47[51]; // @[wallace.scala 69:18]
  assign FullAdder_130_io_b = io_pp_48[50]; // @[wallace.scala 70:18]
  assign FullAdder_130_io_ci = io_pp_49[49]; // @[wallace.scala 71:19]
  assign FullAdder_131_io_a = io_pp_50[48]; // @[wallace.scala 69:18]
  assign FullAdder_131_io_b = io_pp_51[47]; // @[wallace.scala 70:18]
  assign FullAdder_131_io_ci = io_pp_52[46]; // @[wallace.scala 71:19]
  assign FullAdder_132_io_a = io_pp_53[45]; // @[wallace.scala 69:18]
  assign FullAdder_132_io_b = io_pp_54[44]; // @[wallace.scala 70:18]
  assign FullAdder_132_io_ci = io_pp_55[43]; // @[wallace.scala 71:19]
  assign FullAdder_133_io_a = io_pp_56[42]; // @[wallace.scala 69:18]
  assign FullAdder_133_io_b = io_pp_57[41]; // @[wallace.scala 70:18]
  assign FullAdder_133_io_ci = io_pp_58[40]; // @[wallace.scala 71:19]
  assign FullAdder_134_io_a = io_pp_59[39]; // @[wallace.scala 69:18]
  assign FullAdder_134_io_b = io_pp_60[38]; // @[wallace.scala 70:18]
  assign FullAdder_134_io_ci = io_pp_61[37]; // @[wallace.scala 71:19]
  assign FullAdder_135_io_a = io_pp_34[63]; // @[wallace.scala 69:18]
  assign FullAdder_135_io_b = io_pp_35[62]; // @[wallace.scala 70:18]
  assign FullAdder_135_io_ci = io_pp_36[61]; // @[wallace.scala 71:19]
  assign FullAdder_136_io_a = io_pp_37[60]; // @[wallace.scala 69:18]
  assign FullAdder_136_io_b = io_pp_38[59]; // @[wallace.scala 70:18]
  assign FullAdder_136_io_ci = io_pp_39[58]; // @[wallace.scala 71:19]
  assign FullAdder_137_io_a = io_pp_40[57]; // @[wallace.scala 69:18]
  assign FullAdder_137_io_b = io_pp_41[56]; // @[wallace.scala 70:18]
  assign FullAdder_137_io_ci = io_pp_42[55]; // @[wallace.scala 71:19]
  assign FullAdder_138_io_a = io_pp_43[54]; // @[wallace.scala 69:18]
  assign FullAdder_138_io_b = io_pp_44[53]; // @[wallace.scala 70:18]
  assign FullAdder_138_io_ci = io_pp_45[52]; // @[wallace.scala 71:19]
  assign FullAdder_139_io_a = io_pp_46[51]; // @[wallace.scala 69:18]
  assign FullAdder_139_io_b = io_pp_47[50]; // @[wallace.scala 70:18]
  assign FullAdder_139_io_ci = io_pp_48[49]; // @[wallace.scala 71:19]
  assign FullAdder_140_io_a = io_pp_49[48]; // @[wallace.scala 69:18]
  assign FullAdder_140_io_b = io_pp_50[47]; // @[wallace.scala 70:18]
  assign FullAdder_140_io_ci = io_pp_51[46]; // @[wallace.scala 71:19]
  assign FullAdder_141_io_a = io_pp_52[45]; // @[wallace.scala 69:18]
  assign FullAdder_141_io_b = io_pp_53[44]; // @[wallace.scala 70:18]
  assign FullAdder_141_io_ci = io_pp_54[43]; // @[wallace.scala 71:19]
  assign FullAdder_142_io_a = io_pp_55[42]; // @[wallace.scala 69:18]
  assign FullAdder_142_io_b = io_pp_56[41]; // @[wallace.scala 70:18]
  assign FullAdder_142_io_ci = io_pp_57[40]; // @[wallace.scala 71:19]
  assign FullAdder_143_io_a = io_pp_58[39]; // @[wallace.scala 69:18]
  assign FullAdder_143_io_b = io_pp_59[38]; // @[wallace.scala 70:18]
  assign FullAdder_143_io_ci = io_pp_60[37]; // @[wallace.scala 71:19]
  assign FullAdder_144_io_a = io_pp_61[36]; // @[wallace.scala 69:18]
  assign FullAdder_144_io_b = io_pp_62[35]; // @[wallace.scala 70:18]
  assign FullAdder_144_io_ci = io_pp_63[34]; // @[wallace.scala 71:19]
  assign FullAdder_145_io_a = io_pp_33[63]; // @[wallace.scala 69:18]
  assign FullAdder_145_io_b = io_pp_34[62]; // @[wallace.scala 70:18]
  assign FullAdder_145_io_ci = io_pp_35[61]; // @[wallace.scala 71:19]
  assign FullAdder_146_io_a = io_pp_36[60]; // @[wallace.scala 69:18]
  assign FullAdder_146_io_b = io_pp_37[59]; // @[wallace.scala 70:18]
  assign FullAdder_146_io_ci = io_pp_38[58]; // @[wallace.scala 71:19]
  assign FullAdder_147_io_a = io_pp_39[57]; // @[wallace.scala 69:18]
  assign FullAdder_147_io_b = io_pp_40[56]; // @[wallace.scala 70:18]
  assign FullAdder_147_io_ci = io_pp_41[55]; // @[wallace.scala 71:19]
  assign FullAdder_148_io_a = io_pp_42[54]; // @[wallace.scala 69:18]
  assign FullAdder_148_io_b = io_pp_43[53]; // @[wallace.scala 70:18]
  assign FullAdder_148_io_ci = io_pp_44[52]; // @[wallace.scala 71:19]
  assign FullAdder_149_io_a = io_pp_45[51]; // @[wallace.scala 69:18]
  assign FullAdder_149_io_b = io_pp_46[50]; // @[wallace.scala 70:18]
  assign FullAdder_149_io_ci = io_pp_47[49]; // @[wallace.scala 71:19]
  assign FullAdder_150_io_a = io_pp_48[48]; // @[wallace.scala 69:18]
  assign FullAdder_150_io_b = io_pp_49[47]; // @[wallace.scala 70:18]
  assign FullAdder_150_io_ci = io_pp_50[46]; // @[wallace.scala 71:19]
  assign FullAdder_151_io_a = io_pp_51[45]; // @[wallace.scala 69:18]
  assign FullAdder_151_io_b = io_pp_52[44]; // @[wallace.scala 70:18]
  assign FullAdder_151_io_ci = io_pp_53[43]; // @[wallace.scala 71:19]
  assign FullAdder_152_io_a = io_pp_54[42]; // @[wallace.scala 69:18]
  assign FullAdder_152_io_b = io_pp_55[41]; // @[wallace.scala 70:18]
  assign FullAdder_152_io_ci = io_pp_56[40]; // @[wallace.scala 71:19]
  assign FullAdder_153_io_a = io_pp_57[39]; // @[wallace.scala 69:18]
  assign FullAdder_153_io_b = io_pp_58[38]; // @[wallace.scala 70:18]
  assign FullAdder_153_io_ci = io_pp_59[37]; // @[wallace.scala 71:19]
  assign FullAdder_154_io_a = io_pp_60[36]; // @[wallace.scala 69:18]
  assign FullAdder_154_io_b = io_pp_61[35]; // @[wallace.scala 70:18]
  assign FullAdder_154_io_ci = io_pp_62[34]; // @[wallace.scala 71:19]
  assign FullAdder_155_io_a = io_pp_32[63]; // @[wallace.scala 69:18]
  assign FullAdder_155_io_b = io_pp_33[62]; // @[wallace.scala 70:18]
  assign FullAdder_155_io_ci = io_pp_34[61]; // @[wallace.scala 71:19]
  assign FullAdder_156_io_a = io_pp_35[60]; // @[wallace.scala 69:18]
  assign FullAdder_156_io_b = io_pp_36[59]; // @[wallace.scala 70:18]
  assign FullAdder_156_io_ci = io_pp_37[58]; // @[wallace.scala 71:19]
  assign FullAdder_157_io_a = io_pp_38[57]; // @[wallace.scala 69:18]
  assign FullAdder_157_io_b = io_pp_39[56]; // @[wallace.scala 70:18]
  assign FullAdder_157_io_ci = io_pp_40[55]; // @[wallace.scala 71:19]
  assign FullAdder_158_io_a = io_pp_41[54]; // @[wallace.scala 69:18]
  assign FullAdder_158_io_b = io_pp_42[53]; // @[wallace.scala 70:18]
  assign FullAdder_158_io_ci = io_pp_43[52]; // @[wallace.scala 71:19]
  assign FullAdder_159_io_a = io_pp_44[51]; // @[wallace.scala 69:18]
  assign FullAdder_159_io_b = io_pp_45[50]; // @[wallace.scala 70:18]
  assign FullAdder_159_io_ci = io_pp_46[49]; // @[wallace.scala 71:19]
  assign FullAdder_160_io_a = io_pp_47[48]; // @[wallace.scala 69:18]
  assign FullAdder_160_io_b = io_pp_48[47]; // @[wallace.scala 70:18]
  assign FullAdder_160_io_ci = io_pp_49[46]; // @[wallace.scala 71:19]
  assign FullAdder_161_io_a = io_pp_50[45]; // @[wallace.scala 69:18]
  assign FullAdder_161_io_b = io_pp_51[44]; // @[wallace.scala 70:18]
  assign FullAdder_161_io_ci = io_pp_52[43]; // @[wallace.scala 71:19]
  assign FullAdder_162_io_a = io_pp_53[42]; // @[wallace.scala 69:18]
  assign FullAdder_162_io_b = io_pp_54[41]; // @[wallace.scala 70:18]
  assign FullAdder_162_io_ci = io_pp_55[40]; // @[wallace.scala 71:19]
  assign FullAdder_163_io_a = io_pp_56[39]; // @[wallace.scala 69:18]
  assign FullAdder_163_io_b = io_pp_57[38]; // @[wallace.scala 70:18]
  assign FullAdder_163_io_ci = io_pp_58[37]; // @[wallace.scala 71:19]
  assign FullAdder_164_io_a = io_pp_59[36]; // @[wallace.scala 69:18]
  assign FullAdder_164_io_b = io_pp_60[35]; // @[wallace.scala 70:18]
  assign FullAdder_164_io_ci = io_pp_61[34]; // @[wallace.scala 71:19]
  assign HalfAdder_7_io_a = io_pp_62[33]; // @[wallace.scala 59:18]
  assign HalfAdder_7_io_b = io_pp_63[32]; // @[wallace.scala 60:18]
  assign FullAdder_165_io_a = io_pp_31[63]; // @[wallace.scala 69:18]
  assign FullAdder_165_io_b = io_pp_32[62]; // @[wallace.scala 70:18]
  assign FullAdder_165_io_ci = io_pp_33[61]; // @[wallace.scala 71:19]
  assign FullAdder_166_io_a = io_pp_34[60]; // @[wallace.scala 69:18]
  assign FullAdder_166_io_b = io_pp_35[59]; // @[wallace.scala 70:18]
  assign FullAdder_166_io_ci = io_pp_36[58]; // @[wallace.scala 71:19]
  assign FullAdder_167_io_a = io_pp_37[57]; // @[wallace.scala 69:18]
  assign FullAdder_167_io_b = io_pp_38[56]; // @[wallace.scala 70:18]
  assign FullAdder_167_io_ci = io_pp_39[55]; // @[wallace.scala 71:19]
  assign FullAdder_168_io_a = io_pp_40[54]; // @[wallace.scala 69:18]
  assign FullAdder_168_io_b = io_pp_41[53]; // @[wallace.scala 70:18]
  assign FullAdder_168_io_ci = io_pp_42[52]; // @[wallace.scala 71:19]
  assign FullAdder_169_io_a = io_pp_43[51]; // @[wallace.scala 69:18]
  assign FullAdder_169_io_b = io_pp_44[50]; // @[wallace.scala 70:18]
  assign FullAdder_169_io_ci = io_pp_45[49]; // @[wallace.scala 71:19]
  assign FullAdder_170_io_a = io_pp_46[48]; // @[wallace.scala 69:18]
  assign FullAdder_170_io_b = io_pp_47[47]; // @[wallace.scala 70:18]
  assign FullAdder_170_io_ci = io_pp_48[46]; // @[wallace.scala 71:19]
  assign FullAdder_171_io_a = io_pp_49[45]; // @[wallace.scala 69:18]
  assign FullAdder_171_io_b = io_pp_50[44]; // @[wallace.scala 70:18]
  assign FullAdder_171_io_ci = io_pp_51[43]; // @[wallace.scala 71:19]
  assign FullAdder_172_io_a = io_pp_52[42]; // @[wallace.scala 69:18]
  assign FullAdder_172_io_b = io_pp_53[41]; // @[wallace.scala 70:18]
  assign FullAdder_172_io_ci = io_pp_54[40]; // @[wallace.scala 71:19]
  assign FullAdder_173_io_a = io_pp_55[39]; // @[wallace.scala 69:18]
  assign FullAdder_173_io_b = io_pp_56[38]; // @[wallace.scala 70:18]
  assign FullAdder_173_io_ci = io_pp_57[37]; // @[wallace.scala 71:19]
  assign FullAdder_174_io_a = io_pp_58[36]; // @[wallace.scala 69:18]
  assign FullAdder_174_io_b = io_pp_59[35]; // @[wallace.scala 70:18]
  assign FullAdder_174_io_ci = io_pp_60[34]; // @[wallace.scala 71:19]
  assign FullAdder_175_io_a = io_pp_61[33]; // @[wallace.scala 69:18]
  assign FullAdder_175_io_b = io_pp_62[32]; // @[wallace.scala 70:18]
  assign FullAdder_175_io_ci = io_pp_63[31]; // @[wallace.scala 71:19]
  assign FullAdder_176_io_a = io_pp_30[63]; // @[wallace.scala 69:18]
  assign FullAdder_176_io_b = io_pp_31[62]; // @[wallace.scala 70:18]
  assign FullAdder_176_io_ci = io_pp_32[61]; // @[wallace.scala 71:19]
  assign FullAdder_177_io_a = io_pp_33[60]; // @[wallace.scala 69:18]
  assign FullAdder_177_io_b = io_pp_34[59]; // @[wallace.scala 70:18]
  assign FullAdder_177_io_ci = io_pp_35[58]; // @[wallace.scala 71:19]
  assign FullAdder_178_io_a = io_pp_36[57]; // @[wallace.scala 69:18]
  assign FullAdder_178_io_b = io_pp_37[56]; // @[wallace.scala 70:18]
  assign FullAdder_178_io_ci = io_pp_38[55]; // @[wallace.scala 71:19]
  assign FullAdder_179_io_a = io_pp_39[54]; // @[wallace.scala 69:18]
  assign FullAdder_179_io_b = io_pp_40[53]; // @[wallace.scala 70:18]
  assign FullAdder_179_io_ci = io_pp_41[52]; // @[wallace.scala 71:19]
  assign FullAdder_180_io_a = io_pp_42[51]; // @[wallace.scala 69:18]
  assign FullAdder_180_io_b = io_pp_43[50]; // @[wallace.scala 70:18]
  assign FullAdder_180_io_ci = io_pp_44[49]; // @[wallace.scala 71:19]
  assign FullAdder_181_io_a = io_pp_45[48]; // @[wallace.scala 69:18]
  assign FullAdder_181_io_b = io_pp_46[47]; // @[wallace.scala 70:18]
  assign FullAdder_181_io_ci = io_pp_47[46]; // @[wallace.scala 71:19]
  assign FullAdder_182_io_a = io_pp_48[45]; // @[wallace.scala 69:18]
  assign FullAdder_182_io_b = io_pp_49[44]; // @[wallace.scala 70:18]
  assign FullAdder_182_io_ci = io_pp_50[43]; // @[wallace.scala 71:19]
  assign FullAdder_183_io_a = io_pp_51[42]; // @[wallace.scala 69:18]
  assign FullAdder_183_io_b = io_pp_52[41]; // @[wallace.scala 70:18]
  assign FullAdder_183_io_ci = io_pp_53[40]; // @[wallace.scala 71:19]
  assign FullAdder_184_io_a = io_pp_54[39]; // @[wallace.scala 69:18]
  assign FullAdder_184_io_b = io_pp_55[38]; // @[wallace.scala 70:18]
  assign FullAdder_184_io_ci = io_pp_56[37]; // @[wallace.scala 71:19]
  assign FullAdder_185_io_a = io_pp_57[36]; // @[wallace.scala 69:18]
  assign FullAdder_185_io_b = io_pp_58[35]; // @[wallace.scala 70:18]
  assign FullAdder_185_io_ci = io_pp_59[34]; // @[wallace.scala 71:19]
  assign FullAdder_186_io_a = io_pp_60[33]; // @[wallace.scala 69:18]
  assign FullAdder_186_io_b = io_pp_61[32]; // @[wallace.scala 70:18]
  assign FullAdder_186_io_ci = io_pp_62[31]; // @[wallace.scala 71:19]
  assign FullAdder_187_io_a = io_pp_29[63]; // @[wallace.scala 69:18]
  assign FullAdder_187_io_b = io_pp_30[62]; // @[wallace.scala 70:18]
  assign FullAdder_187_io_ci = io_pp_31[61]; // @[wallace.scala 71:19]
  assign FullAdder_188_io_a = io_pp_32[60]; // @[wallace.scala 69:18]
  assign FullAdder_188_io_b = io_pp_33[59]; // @[wallace.scala 70:18]
  assign FullAdder_188_io_ci = io_pp_34[58]; // @[wallace.scala 71:19]
  assign FullAdder_189_io_a = io_pp_35[57]; // @[wallace.scala 69:18]
  assign FullAdder_189_io_b = io_pp_36[56]; // @[wallace.scala 70:18]
  assign FullAdder_189_io_ci = io_pp_37[55]; // @[wallace.scala 71:19]
  assign FullAdder_190_io_a = io_pp_38[54]; // @[wallace.scala 69:18]
  assign FullAdder_190_io_b = io_pp_39[53]; // @[wallace.scala 70:18]
  assign FullAdder_190_io_ci = io_pp_40[52]; // @[wallace.scala 71:19]
  assign FullAdder_191_io_a = io_pp_41[51]; // @[wallace.scala 69:18]
  assign FullAdder_191_io_b = io_pp_42[50]; // @[wallace.scala 70:18]
  assign FullAdder_191_io_ci = io_pp_43[49]; // @[wallace.scala 71:19]
  assign FullAdder_192_io_a = io_pp_44[48]; // @[wallace.scala 69:18]
  assign FullAdder_192_io_b = io_pp_45[47]; // @[wallace.scala 70:18]
  assign FullAdder_192_io_ci = io_pp_46[46]; // @[wallace.scala 71:19]
  assign FullAdder_193_io_a = io_pp_47[45]; // @[wallace.scala 69:18]
  assign FullAdder_193_io_b = io_pp_48[44]; // @[wallace.scala 70:18]
  assign FullAdder_193_io_ci = io_pp_49[43]; // @[wallace.scala 71:19]
  assign FullAdder_194_io_a = io_pp_50[42]; // @[wallace.scala 69:18]
  assign FullAdder_194_io_b = io_pp_51[41]; // @[wallace.scala 70:18]
  assign FullAdder_194_io_ci = io_pp_52[40]; // @[wallace.scala 71:19]
  assign FullAdder_195_io_a = io_pp_53[39]; // @[wallace.scala 69:18]
  assign FullAdder_195_io_b = io_pp_54[38]; // @[wallace.scala 70:18]
  assign FullAdder_195_io_ci = io_pp_55[37]; // @[wallace.scala 71:19]
  assign FullAdder_196_io_a = io_pp_56[36]; // @[wallace.scala 69:18]
  assign FullAdder_196_io_b = io_pp_57[35]; // @[wallace.scala 70:18]
  assign FullAdder_196_io_ci = io_pp_58[34]; // @[wallace.scala 71:19]
  assign FullAdder_197_io_a = io_pp_59[33]; // @[wallace.scala 69:18]
  assign FullAdder_197_io_b = io_pp_60[32]; // @[wallace.scala 70:18]
  assign FullAdder_197_io_ci = io_pp_61[31]; // @[wallace.scala 71:19]
  assign HalfAdder_8_io_a = io_pp_62[30]; // @[wallace.scala 59:18]
  assign HalfAdder_8_io_b = io_pp_63[29]; // @[wallace.scala 60:18]
  assign FullAdder_198_io_a = io_pp_28[63]; // @[wallace.scala 69:18]
  assign FullAdder_198_io_b = io_pp_29[62]; // @[wallace.scala 70:18]
  assign FullAdder_198_io_ci = io_pp_30[61]; // @[wallace.scala 71:19]
  assign FullAdder_199_io_a = io_pp_31[60]; // @[wallace.scala 69:18]
  assign FullAdder_199_io_b = io_pp_32[59]; // @[wallace.scala 70:18]
  assign FullAdder_199_io_ci = io_pp_33[58]; // @[wallace.scala 71:19]
  assign FullAdder_200_io_a = io_pp_34[57]; // @[wallace.scala 69:18]
  assign FullAdder_200_io_b = io_pp_35[56]; // @[wallace.scala 70:18]
  assign FullAdder_200_io_ci = io_pp_36[55]; // @[wallace.scala 71:19]
  assign FullAdder_201_io_a = io_pp_37[54]; // @[wallace.scala 69:18]
  assign FullAdder_201_io_b = io_pp_38[53]; // @[wallace.scala 70:18]
  assign FullAdder_201_io_ci = io_pp_39[52]; // @[wallace.scala 71:19]
  assign FullAdder_202_io_a = io_pp_40[51]; // @[wallace.scala 69:18]
  assign FullAdder_202_io_b = io_pp_41[50]; // @[wallace.scala 70:18]
  assign FullAdder_202_io_ci = io_pp_42[49]; // @[wallace.scala 71:19]
  assign FullAdder_203_io_a = io_pp_43[48]; // @[wallace.scala 69:18]
  assign FullAdder_203_io_b = io_pp_44[47]; // @[wallace.scala 70:18]
  assign FullAdder_203_io_ci = io_pp_45[46]; // @[wallace.scala 71:19]
  assign FullAdder_204_io_a = io_pp_46[45]; // @[wallace.scala 69:18]
  assign FullAdder_204_io_b = io_pp_47[44]; // @[wallace.scala 70:18]
  assign FullAdder_204_io_ci = io_pp_48[43]; // @[wallace.scala 71:19]
  assign FullAdder_205_io_a = io_pp_49[42]; // @[wallace.scala 69:18]
  assign FullAdder_205_io_b = io_pp_50[41]; // @[wallace.scala 70:18]
  assign FullAdder_205_io_ci = io_pp_51[40]; // @[wallace.scala 71:19]
  assign FullAdder_206_io_a = io_pp_52[39]; // @[wallace.scala 69:18]
  assign FullAdder_206_io_b = io_pp_53[38]; // @[wallace.scala 70:18]
  assign FullAdder_206_io_ci = io_pp_54[37]; // @[wallace.scala 71:19]
  assign FullAdder_207_io_a = io_pp_55[36]; // @[wallace.scala 69:18]
  assign FullAdder_207_io_b = io_pp_56[35]; // @[wallace.scala 70:18]
  assign FullAdder_207_io_ci = io_pp_57[34]; // @[wallace.scala 71:19]
  assign FullAdder_208_io_a = io_pp_58[33]; // @[wallace.scala 69:18]
  assign FullAdder_208_io_b = io_pp_59[32]; // @[wallace.scala 70:18]
  assign FullAdder_208_io_ci = io_pp_60[31]; // @[wallace.scala 71:19]
  assign FullAdder_209_io_a = io_pp_61[30]; // @[wallace.scala 69:18]
  assign FullAdder_209_io_b = io_pp_62[29]; // @[wallace.scala 70:18]
  assign FullAdder_209_io_ci = io_pp_63[28]; // @[wallace.scala 71:19]
  assign FullAdder_210_io_a = io_pp_27[63]; // @[wallace.scala 69:18]
  assign FullAdder_210_io_b = io_pp_28[62]; // @[wallace.scala 70:18]
  assign FullAdder_210_io_ci = io_pp_29[61]; // @[wallace.scala 71:19]
  assign FullAdder_211_io_a = io_pp_30[60]; // @[wallace.scala 69:18]
  assign FullAdder_211_io_b = io_pp_31[59]; // @[wallace.scala 70:18]
  assign FullAdder_211_io_ci = io_pp_32[58]; // @[wallace.scala 71:19]
  assign FullAdder_212_io_a = io_pp_33[57]; // @[wallace.scala 69:18]
  assign FullAdder_212_io_b = io_pp_34[56]; // @[wallace.scala 70:18]
  assign FullAdder_212_io_ci = io_pp_35[55]; // @[wallace.scala 71:19]
  assign FullAdder_213_io_a = io_pp_36[54]; // @[wallace.scala 69:18]
  assign FullAdder_213_io_b = io_pp_37[53]; // @[wallace.scala 70:18]
  assign FullAdder_213_io_ci = io_pp_38[52]; // @[wallace.scala 71:19]
  assign FullAdder_214_io_a = io_pp_39[51]; // @[wallace.scala 69:18]
  assign FullAdder_214_io_b = io_pp_40[50]; // @[wallace.scala 70:18]
  assign FullAdder_214_io_ci = io_pp_41[49]; // @[wallace.scala 71:19]
  assign FullAdder_215_io_a = io_pp_42[48]; // @[wallace.scala 69:18]
  assign FullAdder_215_io_b = io_pp_43[47]; // @[wallace.scala 70:18]
  assign FullAdder_215_io_ci = io_pp_44[46]; // @[wallace.scala 71:19]
  assign FullAdder_216_io_a = io_pp_45[45]; // @[wallace.scala 69:18]
  assign FullAdder_216_io_b = io_pp_46[44]; // @[wallace.scala 70:18]
  assign FullAdder_216_io_ci = io_pp_47[43]; // @[wallace.scala 71:19]
  assign FullAdder_217_io_a = io_pp_48[42]; // @[wallace.scala 69:18]
  assign FullAdder_217_io_b = io_pp_49[41]; // @[wallace.scala 70:18]
  assign FullAdder_217_io_ci = io_pp_50[40]; // @[wallace.scala 71:19]
  assign FullAdder_218_io_a = io_pp_51[39]; // @[wallace.scala 69:18]
  assign FullAdder_218_io_b = io_pp_52[38]; // @[wallace.scala 70:18]
  assign FullAdder_218_io_ci = io_pp_53[37]; // @[wallace.scala 71:19]
  assign FullAdder_219_io_a = io_pp_54[36]; // @[wallace.scala 69:18]
  assign FullAdder_219_io_b = io_pp_55[35]; // @[wallace.scala 70:18]
  assign FullAdder_219_io_ci = io_pp_56[34]; // @[wallace.scala 71:19]
  assign FullAdder_220_io_a = io_pp_57[33]; // @[wallace.scala 69:18]
  assign FullAdder_220_io_b = io_pp_58[32]; // @[wallace.scala 70:18]
  assign FullAdder_220_io_ci = io_pp_59[31]; // @[wallace.scala 71:19]
  assign FullAdder_221_io_a = io_pp_60[30]; // @[wallace.scala 69:18]
  assign FullAdder_221_io_b = io_pp_61[29]; // @[wallace.scala 70:18]
  assign FullAdder_221_io_ci = io_pp_62[28]; // @[wallace.scala 71:19]
  assign FullAdder_222_io_a = io_pp_26[63]; // @[wallace.scala 69:18]
  assign FullAdder_222_io_b = io_pp_27[62]; // @[wallace.scala 70:18]
  assign FullAdder_222_io_ci = io_pp_28[61]; // @[wallace.scala 71:19]
  assign FullAdder_223_io_a = io_pp_29[60]; // @[wallace.scala 69:18]
  assign FullAdder_223_io_b = io_pp_30[59]; // @[wallace.scala 70:18]
  assign FullAdder_223_io_ci = io_pp_31[58]; // @[wallace.scala 71:19]
  assign FullAdder_224_io_a = io_pp_32[57]; // @[wallace.scala 69:18]
  assign FullAdder_224_io_b = io_pp_33[56]; // @[wallace.scala 70:18]
  assign FullAdder_224_io_ci = io_pp_34[55]; // @[wallace.scala 71:19]
  assign FullAdder_225_io_a = io_pp_35[54]; // @[wallace.scala 69:18]
  assign FullAdder_225_io_b = io_pp_36[53]; // @[wallace.scala 70:18]
  assign FullAdder_225_io_ci = io_pp_37[52]; // @[wallace.scala 71:19]
  assign FullAdder_226_io_a = io_pp_38[51]; // @[wallace.scala 69:18]
  assign FullAdder_226_io_b = io_pp_39[50]; // @[wallace.scala 70:18]
  assign FullAdder_226_io_ci = io_pp_40[49]; // @[wallace.scala 71:19]
  assign FullAdder_227_io_a = io_pp_41[48]; // @[wallace.scala 69:18]
  assign FullAdder_227_io_b = io_pp_42[47]; // @[wallace.scala 70:18]
  assign FullAdder_227_io_ci = io_pp_43[46]; // @[wallace.scala 71:19]
  assign FullAdder_228_io_a = io_pp_44[45]; // @[wallace.scala 69:18]
  assign FullAdder_228_io_b = io_pp_45[44]; // @[wallace.scala 70:18]
  assign FullAdder_228_io_ci = io_pp_46[43]; // @[wallace.scala 71:19]
  assign FullAdder_229_io_a = io_pp_47[42]; // @[wallace.scala 69:18]
  assign FullAdder_229_io_b = io_pp_48[41]; // @[wallace.scala 70:18]
  assign FullAdder_229_io_ci = io_pp_49[40]; // @[wallace.scala 71:19]
  assign FullAdder_230_io_a = io_pp_50[39]; // @[wallace.scala 69:18]
  assign FullAdder_230_io_b = io_pp_51[38]; // @[wallace.scala 70:18]
  assign FullAdder_230_io_ci = io_pp_52[37]; // @[wallace.scala 71:19]
  assign FullAdder_231_io_a = io_pp_53[36]; // @[wallace.scala 69:18]
  assign FullAdder_231_io_b = io_pp_54[35]; // @[wallace.scala 70:18]
  assign FullAdder_231_io_ci = io_pp_55[34]; // @[wallace.scala 71:19]
  assign FullAdder_232_io_a = io_pp_56[33]; // @[wallace.scala 69:18]
  assign FullAdder_232_io_b = io_pp_57[32]; // @[wallace.scala 70:18]
  assign FullAdder_232_io_ci = io_pp_58[31]; // @[wallace.scala 71:19]
  assign FullAdder_233_io_a = io_pp_59[30]; // @[wallace.scala 69:18]
  assign FullAdder_233_io_b = io_pp_60[29]; // @[wallace.scala 70:18]
  assign FullAdder_233_io_ci = io_pp_61[28]; // @[wallace.scala 71:19]
  assign HalfAdder_9_io_a = io_pp_62[27]; // @[wallace.scala 59:18]
  assign HalfAdder_9_io_b = io_pp_63[26]; // @[wallace.scala 60:18]
  assign FullAdder_234_io_a = io_pp_25[63]; // @[wallace.scala 69:18]
  assign FullAdder_234_io_b = io_pp_26[62]; // @[wallace.scala 70:18]
  assign FullAdder_234_io_ci = io_pp_27[61]; // @[wallace.scala 71:19]
  assign FullAdder_235_io_a = io_pp_28[60]; // @[wallace.scala 69:18]
  assign FullAdder_235_io_b = io_pp_29[59]; // @[wallace.scala 70:18]
  assign FullAdder_235_io_ci = io_pp_30[58]; // @[wallace.scala 71:19]
  assign FullAdder_236_io_a = io_pp_31[57]; // @[wallace.scala 69:18]
  assign FullAdder_236_io_b = io_pp_32[56]; // @[wallace.scala 70:18]
  assign FullAdder_236_io_ci = io_pp_33[55]; // @[wallace.scala 71:19]
  assign FullAdder_237_io_a = io_pp_34[54]; // @[wallace.scala 69:18]
  assign FullAdder_237_io_b = io_pp_35[53]; // @[wallace.scala 70:18]
  assign FullAdder_237_io_ci = io_pp_36[52]; // @[wallace.scala 71:19]
  assign FullAdder_238_io_a = io_pp_37[51]; // @[wallace.scala 69:18]
  assign FullAdder_238_io_b = io_pp_38[50]; // @[wallace.scala 70:18]
  assign FullAdder_238_io_ci = io_pp_39[49]; // @[wallace.scala 71:19]
  assign FullAdder_239_io_a = io_pp_40[48]; // @[wallace.scala 69:18]
  assign FullAdder_239_io_b = io_pp_41[47]; // @[wallace.scala 70:18]
  assign FullAdder_239_io_ci = io_pp_42[46]; // @[wallace.scala 71:19]
  assign FullAdder_240_io_a = io_pp_43[45]; // @[wallace.scala 69:18]
  assign FullAdder_240_io_b = io_pp_44[44]; // @[wallace.scala 70:18]
  assign FullAdder_240_io_ci = io_pp_45[43]; // @[wallace.scala 71:19]
  assign FullAdder_241_io_a = io_pp_46[42]; // @[wallace.scala 69:18]
  assign FullAdder_241_io_b = io_pp_47[41]; // @[wallace.scala 70:18]
  assign FullAdder_241_io_ci = io_pp_48[40]; // @[wallace.scala 71:19]
  assign FullAdder_242_io_a = io_pp_49[39]; // @[wallace.scala 69:18]
  assign FullAdder_242_io_b = io_pp_50[38]; // @[wallace.scala 70:18]
  assign FullAdder_242_io_ci = io_pp_51[37]; // @[wallace.scala 71:19]
  assign FullAdder_243_io_a = io_pp_52[36]; // @[wallace.scala 69:18]
  assign FullAdder_243_io_b = io_pp_53[35]; // @[wallace.scala 70:18]
  assign FullAdder_243_io_ci = io_pp_54[34]; // @[wallace.scala 71:19]
  assign FullAdder_244_io_a = io_pp_55[33]; // @[wallace.scala 69:18]
  assign FullAdder_244_io_b = io_pp_56[32]; // @[wallace.scala 70:18]
  assign FullAdder_244_io_ci = io_pp_57[31]; // @[wallace.scala 71:19]
  assign FullAdder_245_io_a = io_pp_58[30]; // @[wallace.scala 69:18]
  assign FullAdder_245_io_b = io_pp_59[29]; // @[wallace.scala 70:18]
  assign FullAdder_245_io_ci = io_pp_60[28]; // @[wallace.scala 71:19]
  assign FullAdder_246_io_a = io_pp_61[27]; // @[wallace.scala 69:18]
  assign FullAdder_246_io_b = io_pp_62[26]; // @[wallace.scala 70:18]
  assign FullAdder_246_io_ci = io_pp_63[25]; // @[wallace.scala 71:19]
  assign FullAdder_247_io_a = io_pp_24[63]; // @[wallace.scala 69:18]
  assign FullAdder_247_io_b = io_pp_25[62]; // @[wallace.scala 70:18]
  assign FullAdder_247_io_ci = io_pp_26[61]; // @[wallace.scala 71:19]
  assign FullAdder_248_io_a = io_pp_27[60]; // @[wallace.scala 69:18]
  assign FullAdder_248_io_b = io_pp_28[59]; // @[wallace.scala 70:18]
  assign FullAdder_248_io_ci = io_pp_29[58]; // @[wallace.scala 71:19]
  assign FullAdder_249_io_a = io_pp_30[57]; // @[wallace.scala 69:18]
  assign FullAdder_249_io_b = io_pp_31[56]; // @[wallace.scala 70:18]
  assign FullAdder_249_io_ci = io_pp_32[55]; // @[wallace.scala 71:19]
  assign FullAdder_250_io_a = io_pp_33[54]; // @[wallace.scala 69:18]
  assign FullAdder_250_io_b = io_pp_34[53]; // @[wallace.scala 70:18]
  assign FullAdder_250_io_ci = io_pp_35[52]; // @[wallace.scala 71:19]
  assign FullAdder_251_io_a = io_pp_36[51]; // @[wallace.scala 69:18]
  assign FullAdder_251_io_b = io_pp_37[50]; // @[wallace.scala 70:18]
  assign FullAdder_251_io_ci = io_pp_38[49]; // @[wallace.scala 71:19]
  assign FullAdder_252_io_a = io_pp_39[48]; // @[wallace.scala 69:18]
  assign FullAdder_252_io_b = io_pp_40[47]; // @[wallace.scala 70:18]
  assign FullAdder_252_io_ci = io_pp_41[46]; // @[wallace.scala 71:19]
  assign FullAdder_253_io_a = io_pp_42[45]; // @[wallace.scala 69:18]
  assign FullAdder_253_io_b = io_pp_43[44]; // @[wallace.scala 70:18]
  assign FullAdder_253_io_ci = io_pp_44[43]; // @[wallace.scala 71:19]
  assign FullAdder_254_io_a = io_pp_45[42]; // @[wallace.scala 69:18]
  assign FullAdder_254_io_b = io_pp_46[41]; // @[wallace.scala 70:18]
  assign FullAdder_254_io_ci = io_pp_47[40]; // @[wallace.scala 71:19]
  assign FullAdder_255_io_a = io_pp_48[39]; // @[wallace.scala 69:18]
  assign FullAdder_255_io_b = io_pp_49[38]; // @[wallace.scala 70:18]
  assign FullAdder_255_io_ci = io_pp_50[37]; // @[wallace.scala 71:19]
  assign FullAdder_256_io_a = io_pp_51[36]; // @[wallace.scala 69:18]
  assign FullAdder_256_io_b = io_pp_52[35]; // @[wallace.scala 70:18]
  assign FullAdder_256_io_ci = io_pp_53[34]; // @[wallace.scala 71:19]
  assign FullAdder_257_io_a = io_pp_54[33]; // @[wallace.scala 69:18]
  assign FullAdder_257_io_b = io_pp_55[32]; // @[wallace.scala 70:18]
  assign FullAdder_257_io_ci = io_pp_56[31]; // @[wallace.scala 71:19]
  assign FullAdder_258_io_a = io_pp_57[30]; // @[wallace.scala 69:18]
  assign FullAdder_258_io_b = io_pp_58[29]; // @[wallace.scala 70:18]
  assign FullAdder_258_io_ci = io_pp_59[28]; // @[wallace.scala 71:19]
  assign FullAdder_259_io_a = io_pp_60[27]; // @[wallace.scala 69:18]
  assign FullAdder_259_io_b = io_pp_61[26]; // @[wallace.scala 70:18]
  assign FullAdder_259_io_ci = io_pp_62[25]; // @[wallace.scala 71:19]
  assign FullAdder_260_io_a = io_pp_23[63]; // @[wallace.scala 69:18]
  assign FullAdder_260_io_b = io_pp_24[62]; // @[wallace.scala 70:18]
  assign FullAdder_260_io_ci = io_pp_25[61]; // @[wallace.scala 71:19]
  assign FullAdder_261_io_a = io_pp_26[60]; // @[wallace.scala 69:18]
  assign FullAdder_261_io_b = io_pp_27[59]; // @[wallace.scala 70:18]
  assign FullAdder_261_io_ci = io_pp_28[58]; // @[wallace.scala 71:19]
  assign FullAdder_262_io_a = io_pp_29[57]; // @[wallace.scala 69:18]
  assign FullAdder_262_io_b = io_pp_30[56]; // @[wallace.scala 70:18]
  assign FullAdder_262_io_ci = io_pp_31[55]; // @[wallace.scala 71:19]
  assign FullAdder_263_io_a = io_pp_32[54]; // @[wallace.scala 69:18]
  assign FullAdder_263_io_b = io_pp_33[53]; // @[wallace.scala 70:18]
  assign FullAdder_263_io_ci = io_pp_34[52]; // @[wallace.scala 71:19]
  assign FullAdder_264_io_a = io_pp_35[51]; // @[wallace.scala 69:18]
  assign FullAdder_264_io_b = io_pp_36[50]; // @[wallace.scala 70:18]
  assign FullAdder_264_io_ci = io_pp_37[49]; // @[wallace.scala 71:19]
  assign FullAdder_265_io_a = io_pp_38[48]; // @[wallace.scala 69:18]
  assign FullAdder_265_io_b = io_pp_39[47]; // @[wallace.scala 70:18]
  assign FullAdder_265_io_ci = io_pp_40[46]; // @[wallace.scala 71:19]
  assign FullAdder_266_io_a = io_pp_41[45]; // @[wallace.scala 69:18]
  assign FullAdder_266_io_b = io_pp_42[44]; // @[wallace.scala 70:18]
  assign FullAdder_266_io_ci = io_pp_43[43]; // @[wallace.scala 71:19]
  assign FullAdder_267_io_a = io_pp_44[42]; // @[wallace.scala 69:18]
  assign FullAdder_267_io_b = io_pp_45[41]; // @[wallace.scala 70:18]
  assign FullAdder_267_io_ci = io_pp_46[40]; // @[wallace.scala 71:19]
  assign FullAdder_268_io_a = io_pp_47[39]; // @[wallace.scala 69:18]
  assign FullAdder_268_io_b = io_pp_48[38]; // @[wallace.scala 70:18]
  assign FullAdder_268_io_ci = io_pp_49[37]; // @[wallace.scala 71:19]
  assign FullAdder_269_io_a = io_pp_50[36]; // @[wallace.scala 69:18]
  assign FullAdder_269_io_b = io_pp_51[35]; // @[wallace.scala 70:18]
  assign FullAdder_269_io_ci = io_pp_52[34]; // @[wallace.scala 71:19]
  assign FullAdder_270_io_a = io_pp_53[33]; // @[wallace.scala 69:18]
  assign FullAdder_270_io_b = io_pp_54[32]; // @[wallace.scala 70:18]
  assign FullAdder_270_io_ci = io_pp_55[31]; // @[wallace.scala 71:19]
  assign FullAdder_271_io_a = io_pp_56[30]; // @[wallace.scala 69:18]
  assign FullAdder_271_io_b = io_pp_57[29]; // @[wallace.scala 70:18]
  assign FullAdder_271_io_ci = io_pp_58[28]; // @[wallace.scala 71:19]
  assign FullAdder_272_io_a = io_pp_59[27]; // @[wallace.scala 69:18]
  assign FullAdder_272_io_b = io_pp_60[26]; // @[wallace.scala 70:18]
  assign FullAdder_272_io_ci = io_pp_61[25]; // @[wallace.scala 71:19]
  assign HalfAdder_10_io_a = io_pp_62[24]; // @[wallace.scala 59:18]
  assign HalfAdder_10_io_b = io_pp_63[23]; // @[wallace.scala 60:18]
  assign FullAdder_273_io_a = io_pp_22[63]; // @[wallace.scala 69:18]
  assign FullAdder_273_io_b = io_pp_23[62]; // @[wallace.scala 70:18]
  assign FullAdder_273_io_ci = io_pp_24[61]; // @[wallace.scala 71:19]
  assign FullAdder_274_io_a = io_pp_25[60]; // @[wallace.scala 69:18]
  assign FullAdder_274_io_b = io_pp_26[59]; // @[wallace.scala 70:18]
  assign FullAdder_274_io_ci = io_pp_27[58]; // @[wallace.scala 71:19]
  assign FullAdder_275_io_a = io_pp_28[57]; // @[wallace.scala 69:18]
  assign FullAdder_275_io_b = io_pp_29[56]; // @[wallace.scala 70:18]
  assign FullAdder_275_io_ci = io_pp_30[55]; // @[wallace.scala 71:19]
  assign FullAdder_276_io_a = io_pp_31[54]; // @[wallace.scala 69:18]
  assign FullAdder_276_io_b = io_pp_32[53]; // @[wallace.scala 70:18]
  assign FullAdder_276_io_ci = io_pp_33[52]; // @[wallace.scala 71:19]
  assign FullAdder_277_io_a = io_pp_34[51]; // @[wallace.scala 69:18]
  assign FullAdder_277_io_b = io_pp_35[50]; // @[wallace.scala 70:18]
  assign FullAdder_277_io_ci = io_pp_36[49]; // @[wallace.scala 71:19]
  assign FullAdder_278_io_a = io_pp_37[48]; // @[wallace.scala 69:18]
  assign FullAdder_278_io_b = io_pp_38[47]; // @[wallace.scala 70:18]
  assign FullAdder_278_io_ci = io_pp_39[46]; // @[wallace.scala 71:19]
  assign FullAdder_279_io_a = io_pp_40[45]; // @[wallace.scala 69:18]
  assign FullAdder_279_io_b = io_pp_41[44]; // @[wallace.scala 70:18]
  assign FullAdder_279_io_ci = io_pp_42[43]; // @[wallace.scala 71:19]
  assign FullAdder_280_io_a = io_pp_43[42]; // @[wallace.scala 69:18]
  assign FullAdder_280_io_b = io_pp_44[41]; // @[wallace.scala 70:18]
  assign FullAdder_280_io_ci = io_pp_45[40]; // @[wallace.scala 71:19]
  assign FullAdder_281_io_a = io_pp_46[39]; // @[wallace.scala 69:18]
  assign FullAdder_281_io_b = io_pp_47[38]; // @[wallace.scala 70:18]
  assign FullAdder_281_io_ci = io_pp_48[37]; // @[wallace.scala 71:19]
  assign FullAdder_282_io_a = io_pp_49[36]; // @[wallace.scala 69:18]
  assign FullAdder_282_io_b = io_pp_50[35]; // @[wallace.scala 70:18]
  assign FullAdder_282_io_ci = io_pp_51[34]; // @[wallace.scala 71:19]
  assign FullAdder_283_io_a = io_pp_52[33]; // @[wallace.scala 69:18]
  assign FullAdder_283_io_b = io_pp_53[32]; // @[wallace.scala 70:18]
  assign FullAdder_283_io_ci = io_pp_54[31]; // @[wallace.scala 71:19]
  assign FullAdder_284_io_a = io_pp_55[30]; // @[wallace.scala 69:18]
  assign FullAdder_284_io_b = io_pp_56[29]; // @[wallace.scala 70:18]
  assign FullAdder_284_io_ci = io_pp_57[28]; // @[wallace.scala 71:19]
  assign FullAdder_285_io_a = io_pp_58[27]; // @[wallace.scala 69:18]
  assign FullAdder_285_io_b = io_pp_59[26]; // @[wallace.scala 70:18]
  assign FullAdder_285_io_ci = io_pp_60[25]; // @[wallace.scala 71:19]
  assign FullAdder_286_io_a = io_pp_61[24]; // @[wallace.scala 69:18]
  assign FullAdder_286_io_b = io_pp_62[23]; // @[wallace.scala 70:18]
  assign FullAdder_286_io_ci = io_pp_63[22]; // @[wallace.scala 71:19]
  assign FullAdder_287_io_a = io_pp_21[63]; // @[wallace.scala 69:18]
  assign FullAdder_287_io_b = io_pp_22[62]; // @[wallace.scala 70:18]
  assign FullAdder_287_io_ci = io_pp_23[61]; // @[wallace.scala 71:19]
  assign FullAdder_288_io_a = io_pp_24[60]; // @[wallace.scala 69:18]
  assign FullAdder_288_io_b = io_pp_25[59]; // @[wallace.scala 70:18]
  assign FullAdder_288_io_ci = io_pp_26[58]; // @[wallace.scala 71:19]
  assign FullAdder_289_io_a = io_pp_27[57]; // @[wallace.scala 69:18]
  assign FullAdder_289_io_b = io_pp_28[56]; // @[wallace.scala 70:18]
  assign FullAdder_289_io_ci = io_pp_29[55]; // @[wallace.scala 71:19]
  assign FullAdder_290_io_a = io_pp_30[54]; // @[wallace.scala 69:18]
  assign FullAdder_290_io_b = io_pp_31[53]; // @[wallace.scala 70:18]
  assign FullAdder_290_io_ci = io_pp_32[52]; // @[wallace.scala 71:19]
  assign FullAdder_291_io_a = io_pp_33[51]; // @[wallace.scala 69:18]
  assign FullAdder_291_io_b = io_pp_34[50]; // @[wallace.scala 70:18]
  assign FullAdder_291_io_ci = io_pp_35[49]; // @[wallace.scala 71:19]
  assign FullAdder_292_io_a = io_pp_36[48]; // @[wallace.scala 69:18]
  assign FullAdder_292_io_b = io_pp_37[47]; // @[wallace.scala 70:18]
  assign FullAdder_292_io_ci = io_pp_38[46]; // @[wallace.scala 71:19]
  assign FullAdder_293_io_a = io_pp_39[45]; // @[wallace.scala 69:18]
  assign FullAdder_293_io_b = io_pp_40[44]; // @[wallace.scala 70:18]
  assign FullAdder_293_io_ci = io_pp_41[43]; // @[wallace.scala 71:19]
  assign FullAdder_294_io_a = io_pp_42[42]; // @[wallace.scala 69:18]
  assign FullAdder_294_io_b = io_pp_43[41]; // @[wallace.scala 70:18]
  assign FullAdder_294_io_ci = io_pp_44[40]; // @[wallace.scala 71:19]
  assign FullAdder_295_io_a = io_pp_45[39]; // @[wallace.scala 69:18]
  assign FullAdder_295_io_b = io_pp_46[38]; // @[wallace.scala 70:18]
  assign FullAdder_295_io_ci = io_pp_47[37]; // @[wallace.scala 71:19]
  assign FullAdder_296_io_a = io_pp_48[36]; // @[wallace.scala 69:18]
  assign FullAdder_296_io_b = io_pp_49[35]; // @[wallace.scala 70:18]
  assign FullAdder_296_io_ci = io_pp_50[34]; // @[wallace.scala 71:19]
  assign FullAdder_297_io_a = io_pp_51[33]; // @[wallace.scala 69:18]
  assign FullAdder_297_io_b = io_pp_52[32]; // @[wallace.scala 70:18]
  assign FullAdder_297_io_ci = io_pp_53[31]; // @[wallace.scala 71:19]
  assign FullAdder_298_io_a = io_pp_54[30]; // @[wallace.scala 69:18]
  assign FullAdder_298_io_b = io_pp_55[29]; // @[wallace.scala 70:18]
  assign FullAdder_298_io_ci = io_pp_56[28]; // @[wallace.scala 71:19]
  assign FullAdder_299_io_a = io_pp_57[27]; // @[wallace.scala 69:18]
  assign FullAdder_299_io_b = io_pp_58[26]; // @[wallace.scala 70:18]
  assign FullAdder_299_io_ci = io_pp_59[25]; // @[wallace.scala 71:19]
  assign FullAdder_300_io_a = io_pp_60[24]; // @[wallace.scala 69:18]
  assign FullAdder_300_io_b = io_pp_61[23]; // @[wallace.scala 70:18]
  assign FullAdder_300_io_ci = io_pp_62[22]; // @[wallace.scala 71:19]
  assign FullAdder_301_io_a = io_pp_20[63]; // @[wallace.scala 69:18]
  assign FullAdder_301_io_b = io_pp_21[62]; // @[wallace.scala 70:18]
  assign FullAdder_301_io_ci = io_pp_22[61]; // @[wallace.scala 71:19]
  assign FullAdder_302_io_a = io_pp_23[60]; // @[wallace.scala 69:18]
  assign FullAdder_302_io_b = io_pp_24[59]; // @[wallace.scala 70:18]
  assign FullAdder_302_io_ci = io_pp_25[58]; // @[wallace.scala 71:19]
  assign FullAdder_303_io_a = io_pp_26[57]; // @[wallace.scala 69:18]
  assign FullAdder_303_io_b = io_pp_27[56]; // @[wallace.scala 70:18]
  assign FullAdder_303_io_ci = io_pp_28[55]; // @[wallace.scala 71:19]
  assign FullAdder_304_io_a = io_pp_29[54]; // @[wallace.scala 69:18]
  assign FullAdder_304_io_b = io_pp_30[53]; // @[wallace.scala 70:18]
  assign FullAdder_304_io_ci = io_pp_31[52]; // @[wallace.scala 71:19]
  assign FullAdder_305_io_a = io_pp_32[51]; // @[wallace.scala 69:18]
  assign FullAdder_305_io_b = io_pp_33[50]; // @[wallace.scala 70:18]
  assign FullAdder_305_io_ci = io_pp_34[49]; // @[wallace.scala 71:19]
  assign FullAdder_306_io_a = io_pp_35[48]; // @[wallace.scala 69:18]
  assign FullAdder_306_io_b = io_pp_36[47]; // @[wallace.scala 70:18]
  assign FullAdder_306_io_ci = io_pp_37[46]; // @[wallace.scala 71:19]
  assign FullAdder_307_io_a = io_pp_38[45]; // @[wallace.scala 69:18]
  assign FullAdder_307_io_b = io_pp_39[44]; // @[wallace.scala 70:18]
  assign FullAdder_307_io_ci = io_pp_40[43]; // @[wallace.scala 71:19]
  assign FullAdder_308_io_a = io_pp_41[42]; // @[wallace.scala 69:18]
  assign FullAdder_308_io_b = io_pp_42[41]; // @[wallace.scala 70:18]
  assign FullAdder_308_io_ci = io_pp_43[40]; // @[wallace.scala 71:19]
  assign FullAdder_309_io_a = io_pp_44[39]; // @[wallace.scala 69:18]
  assign FullAdder_309_io_b = io_pp_45[38]; // @[wallace.scala 70:18]
  assign FullAdder_309_io_ci = io_pp_46[37]; // @[wallace.scala 71:19]
  assign FullAdder_310_io_a = io_pp_47[36]; // @[wallace.scala 69:18]
  assign FullAdder_310_io_b = io_pp_48[35]; // @[wallace.scala 70:18]
  assign FullAdder_310_io_ci = io_pp_49[34]; // @[wallace.scala 71:19]
  assign FullAdder_311_io_a = io_pp_50[33]; // @[wallace.scala 69:18]
  assign FullAdder_311_io_b = io_pp_51[32]; // @[wallace.scala 70:18]
  assign FullAdder_311_io_ci = io_pp_52[31]; // @[wallace.scala 71:19]
  assign FullAdder_312_io_a = io_pp_53[30]; // @[wallace.scala 69:18]
  assign FullAdder_312_io_b = io_pp_54[29]; // @[wallace.scala 70:18]
  assign FullAdder_312_io_ci = io_pp_55[28]; // @[wallace.scala 71:19]
  assign FullAdder_313_io_a = io_pp_56[27]; // @[wallace.scala 69:18]
  assign FullAdder_313_io_b = io_pp_57[26]; // @[wallace.scala 70:18]
  assign FullAdder_313_io_ci = io_pp_58[25]; // @[wallace.scala 71:19]
  assign FullAdder_314_io_a = io_pp_59[24]; // @[wallace.scala 69:18]
  assign FullAdder_314_io_b = io_pp_60[23]; // @[wallace.scala 70:18]
  assign FullAdder_314_io_ci = io_pp_61[22]; // @[wallace.scala 71:19]
  assign HalfAdder_11_io_a = io_pp_62[21]; // @[wallace.scala 59:18]
  assign HalfAdder_11_io_b = io_pp_63[20]; // @[wallace.scala 60:18]
  assign FullAdder_315_io_a = io_pp_19[63]; // @[wallace.scala 69:18]
  assign FullAdder_315_io_b = io_pp_20[62]; // @[wallace.scala 70:18]
  assign FullAdder_315_io_ci = io_pp_21[61]; // @[wallace.scala 71:19]
  assign FullAdder_316_io_a = io_pp_22[60]; // @[wallace.scala 69:18]
  assign FullAdder_316_io_b = io_pp_23[59]; // @[wallace.scala 70:18]
  assign FullAdder_316_io_ci = io_pp_24[58]; // @[wallace.scala 71:19]
  assign FullAdder_317_io_a = io_pp_25[57]; // @[wallace.scala 69:18]
  assign FullAdder_317_io_b = io_pp_26[56]; // @[wallace.scala 70:18]
  assign FullAdder_317_io_ci = io_pp_27[55]; // @[wallace.scala 71:19]
  assign FullAdder_318_io_a = io_pp_28[54]; // @[wallace.scala 69:18]
  assign FullAdder_318_io_b = io_pp_29[53]; // @[wallace.scala 70:18]
  assign FullAdder_318_io_ci = io_pp_30[52]; // @[wallace.scala 71:19]
  assign FullAdder_319_io_a = io_pp_31[51]; // @[wallace.scala 69:18]
  assign FullAdder_319_io_b = io_pp_32[50]; // @[wallace.scala 70:18]
  assign FullAdder_319_io_ci = io_pp_33[49]; // @[wallace.scala 71:19]
  assign FullAdder_320_io_a = io_pp_34[48]; // @[wallace.scala 69:18]
  assign FullAdder_320_io_b = io_pp_35[47]; // @[wallace.scala 70:18]
  assign FullAdder_320_io_ci = io_pp_36[46]; // @[wallace.scala 71:19]
  assign FullAdder_321_io_a = io_pp_37[45]; // @[wallace.scala 69:18]
  assign FullAdder_321_io_b = io_pp_38[44]; // @[wallace.scala 70:18]
  assign FullAdder_321_io_ci = io_pp_39[43]; // @[wallace.scala 71:19]
  assign FullAdder_322_io_a = io_pp_40[42]; // @[wallace.scala 69:18]
  assign FullAdder_322_io_b = io_pp_41[41]; // @[wallace.scala 70:18]
  assign FullAdder_322_io_ci = io_pp_42[40]; // @[wallace.scala 71:19]
  assign FullAdder_323_io_a = io_pp_43[39]; // @[wallace.scala 69:18]
  assign FullAdder_323_io_b = io_pp_44[38]; // @[wallace.scala 70:18]
  assign FullAdder_323_io_ci = io_pp_45[37]; // @[wallace.scala 71:19]
  assign FullAdder_324_io_a = io_pp_46[36]; // @[wallace.scala 69:18]
  assign FullAdder_324_io_b = io_pp_47[35]; // @[wallace.scala 70:18]
  assign FullAdder_324_io_ci = io_pp_48[34]; // @[wallace.scala 71:19]
  assign FullAdder_325_io_a = io_pp_49[33]; // @[wallace.scala 69:18]
  assign FullAdder_325_io_b = io_pp_50[32]; // @[wallace.scala 70:18]
  assign FullAdder_325_io_ci = io_pp_51[31]; // @[wallace.scala 71:19]
  assign FullAdder_326_io_a = io_pp_52[30]; // @[wallace.scala 69:18]
  assign FullAdder_326_io_b = io_pp_53[29]; // @[wallace.scala 70:18]
  assign FullAdder_326_io_ci = io_pp_54[28]; // @[wallace.scala 71:19]
  assign FullAdder_327_io_a = io_pp_55[27]; // @[wallace.scala 69:18]
  assign FullAdder_327_io_b = io_pp_56[26]; // @[wallace.scala 70:18]
  assign FullAdder_327_io_ci = io_pp_57[25]; // @[wallace.scala 71:19]
  assign FullAdder_328_io_a = io_pp_58[24]; // @[wallace.scala 69:18]
  assign FullAdder_328_io_b = io_pp_59[23]; // @[wallace.scala 70:18]
  assign FullAdder_328_io_ci = io_pp_60[22]; // @[wallace.scala 71:19]
  assign FullAdder_329_io_a = io_pp_61[21]; // @[wallace.scala 69:18]
  assign FullAdder_329_io_b = io_pp_62[20]; // @[wallace.scala 70:18]
  assign FullAdder_329_io_ci = io_pp_63[19]; // @[wallace.scala 71:19]
  assign FullAdder_330_io_a = io_pp_18[63]; // @[wallace.scala 69:18]
  assign FullAdder_330_io_b = io_pp_19[62]; // @[wallace.scala 70:18]
  assign FullAdder_330_io_ci = io_pp_20[61]; // @[wallace.scala 71:19]
  assign FullAdder_331_io_a = io_pp_21[60]; // @[wallace.scala 69:18]
  assign FullAdder_331_io_b = io_pp_22[59]; // @[wallace.scala 70:18]
  assign FullAdder_331_io_ci = io_pp_23[58]; // @[wallace.scala 71:19]
  assign FullAdder_332_io_a = io_pp_24[57]; // @[wallace.scala 69:18]
  assign FullAdder_332_io_b = io_pp_25[56]; // @[wallace.scala 70:18]
  assign FullAdder_332_io_ci = io_pp_26[55]; // @[wallace.scala 71:19]
  assign FullAdder_333_io_a = io_pp_27[54]; // @[wallace.scala 69:18]
  assign FullAdder_333_io_b = io_pp_28[53]; // @[wallace.scala 70:18]
  assign FullAdder_333_io_ci = io_pp_29[52]; // @[wallace.scala 71:19]
  assign FullAdder_334_io_a = io_pp_30[51]; // @[wallace.scala 69:18]
  assign FullAdder_334_io_b = io_pp_31[50]; // @[wallace.scala 70:18]
  assign FullAdder_334_io_ci = io_pp_32[49]; // @[wallace.scala 71:19]
  assign FullAdder_335_io_a = io_pp_33[48]; // @[wallace.scala 69:18]
  assign FullAdder_335_io_b = io_pp_34[47]; // @[wallace.scala 70:18]
  assign FullAdder_335_io_ci = io_pp_35[46]; // @[wallace.scala 71:19]
  assign FullAdder_336_io_a = io_pp_36[45]; // @[wallace.scala 69:18]
  assign FullAdder_336_io_b = io_pp_37[44]; // @[wallace.scala 70:18]
  assign FullAdder_336_io_ci = io_pp_38[43]; // @[wallace.scala 71:19]
  assign FullAdder_337_io_a = io_pp_39[42]; // @[wallace.scala 69:18]
  assign FullAdder_337_io_b = io_pp_40[41]; // @[wallace.scala 70:18]
  assign FullAdder_337_io_ci = io_pp_41[40]; // @[wallace.scala 71:19]
  assign FullAdder_338_io_a = io_pp_42[39]; // @[wallace.scala 69:18]
  assign FullAdder_338_io_b = io_pp_43[38]; // @[wallace.scala 70:18]
  assign FullAdder_338_io_ci = io_pp_44[37]; // @[wallace.scala 71:19]
  assign FullAdder_339_io_a = io_pp_45[36]; // @[wallace.scala 69:18]
  assign FullAdder_339_io_b = io_pp_46[35]; // @[wallace.scala 70:18]
  assign FullAdder_339_io_ci = io_pp_47[34]; // @[wallace.scala 71:19]
  assign FullAdder_340_io_a = io_pp_48[33]; // @[wallace.scala 69:18]
  assign FullAdder_340_io_b = io_pp_49[32]; // @[wallace.scala 70:18]
  assign FullAdder_340_io_ci = io_pp_50[31]; // @[wallace.scala 71:19]
  assign FullAdder_341_io_a = io_pp_51[30]; // @[wallace.scala 69:18]
  assign FullAdder_341_io_b = io_pp_52[29]; // @[wallace.scala 70:18]
  assign FullAdder_341_io_ci = io_pp_53[28]; // @[wallace.scala 71:19]
  assign FullAdder_342_io_a = io_pp_54[27]; // @[wallace.scala 69:18]
  assign FullAdder_342_io_b = io_pp_55[26]; // @[wallace.scala 70:18]
  assign FullAdder_342_io_ci = io_pp_56[25]; // @[wallace.scala 71:19]
  assign FullAdder_343_io_a = io_pp_57[24]; // @[wallace.scala 69:18]
  assign FullAdder_343_io_b = io_pp_58[23]; // @[wallace.scala 70:18]
  assign FullAdder_343_io_ci = io_pp_59[22]; // @[wallace.scala 71:19]
  assign FullAdder_344_io_a = io_pp_60[21]; // @[wallace.scala 69:18]
  assign FullAdder_344_io_b = io_pp_61[20]; // @[wallace.scala 70:18]
  assign FullAdder_344_io_ci = io_pp_62[19]; // @[wallace.scala 71:19]
  assign FullAdder_345_io_a = io_pp_17[63]; // @[wallace.scala 69:18]
  assign FullAdder_345_io_b = io_pp_18[62]; // @[wallace.scala 70:18]
  assign FullAdder_345_io_ci = io_pp_19[61]; // @[wallace.scala 71:19]
  assign FullAdder_346_io_a = io_pp_20[60]; // @[wallace.scala 69:18]
  assign FullAdder_346_io_b = io_pp_21[59]; // @[wallace.scala 70:18]
  assign FullAdder_346_io_ci = io_pp_22[58]; // @[wallace.scala 71:19]
  assign FullAdder_347_io_a = io_pp_23[57]; // @[wallace.scala 69:18]
  assign FullAdder_347_io_b = io_pp_24[56]; // @[wallace.scala 70:18]
  assign FullAdder_347_io_ci = io_pp_25[55]; // @[wallace.scala 71:19]
  assign FullAdder_348_io_a = io_pp_26[54]; // @[wallace.scala 69:18]
  assign FullAdder_348_io_b = io_pp_27[53]; // @[wallace.scala 70:18]
  assign FullAdder_348_io_ci = io_pp_28[52]; // @[wallace.scala 71:19]
  assign FullAdder_349_io_a = io_pp_29[51]; // @[wallace.scala 69:18]
  assign FullAdder_349_io_b = io_pp_30[50]; // @[wallace.scala 70:18]
  assign FullAdder_349_io_ci = io_pp_31[49]; // @[wallace.scala 71:19]
  assign FullAdder_350_io_a = io_pp_32[48]; // @[wallace.scala 69:18]
  assign FullAdder_350_io_b = io_pp_33[47]; // @[wallace.scala 70:18]
  assign FullAdder_350_io_ci = io_pp_34[46]; // @[wallace.scala 71:19]
  assign FullAdder_351_io_a = io_pp_35[45]; // @[wallace.scala 69:18]
  assign FullAdder_351_io_b = io_pp_36[44]; // @[wallace.scala 70:18]
  assign FullAdder_351_io_ci = io_pp_37[43]; // @[wallace.scala 71:19]
  assign FullAdder_352_io_a = io_pp_38[42]; // @[wallace.scala 69:18]
  assign FullAdder_352_io_b = io_pp_39[41]; // @[wallace.scala 70:18]
  assign FullAdder_352_io_ci = io_pp_40[40]; // @[wallace.scala 71:19]
  assign FullAdder_353_io_a = io_pp_41[39]; // @[wallace.scala 69:18]
  assign FullAdder_353_io_b = io_pp_42[38]; // @[wallace.scala 70:18]
  assign FullAdder_353_io_ci = io_pp_43[37]; // @[wallace.scala 71:19]
  assign FullAdder_354_io_a = io_pp_44[36]; // @[wallace.scala 69:18]
  assign FullAdder_354_io_b = io_pp_45[35]; // @[wallace.scala 70:18]
  assign FullAdder_354_io_ci = io_pp_46[34]; // @[wallace.scala 71:19]
  assign FullAdder_355_io_a = io_pp_47[33]; // @[wallace.scala 69:18]
  assign FullAdder_355_io_b = io_pp_48[32]; // @[wallace.scala 70:18]
  assign FullAdder_355_io_ci = io_pp_49[31]; // @[wallace.scala 71:19]
  assign FullAdder_356_io_a = io_pp_50[30]; // @[wallace.scala 69:18]
  assign FullAdder_356_io_b = io_pp_51[29]; // @[wallace.scala 70:18]
  assign FullAdder_356_io_ci = io_pp_52[28]; // @[wallace.scala 71:19]
  assign FullAdder_357_io_a = io_pp_53[27]; // @[wallace.scala 69:18]
  assign FullAdder_357_io_b = io_pp_54[26]; // @[wallace.scala 70:18]
  assign FullAdder_357_io_ci = io_pp_55[25]; // @[wallace.scala 71:19]
  assign FullAdder_358_io_a = io_pp_56[24]; // @[wallace.scala 69:18]
  assign FullAdder_358_io_b = io_pp_57[23]; // @[wallace.scala 70:18]
  assign FullAdder_358_io_ci = io_pp_58[22]; // @[wallace.scala 71:19]
  assign FullAdder_359_io_a = io_pp_59[21]; // @[wallace.scala 69:18]
  assign FullAdder_359_io_b = io_pp_60[20]; // @[wallace.scala 70:18]
  assign FullAdder_359_io_ci = io_pp_61[19]; // @[wallace.scala 71:19]
  assign HalfAdder_12_io_a = io_pp_62[18]; // @[wallace.scala 59:18]
  assign HalfAdder_12_io_b = io_pp_63[17]; // @[wallace.scala 60:18]
  assign FullAdder_360_io_a = io_pp_16[63]; // @[wallace.scala 69:18]
  assign FullAdder_360_io_b = io_pp_17[62]; // @[wallace.scala 70:18]
  assign FullAdder_360_io_ci = io_pp_18[61]; // @[wallace.scala 71:19]
  assign FullAdder_361_io_a = io_pp_19[60]; // @[wallace.scala 69:18]
  assign FullAdder_361_io_b = io_pp_20[59]; // @[wallace.scala 70:18]
  assign FullAdder_361_io_ci = io_pp_21[58]; // @[wallace.scala 71:19]
  assign FullAdder_362_io_a = io_pp_22[57]; // @[wallace.scala 69:18]
  assign FullAdder_362_io_b = io_pp_23[56]; // @[wallace.scala 70:18]
  assign FullAdder_362_io_ci = io_pp_24[55]; // @[wallace.scala 71:19]
  assign FullAdder_363_io_a = io_pp_25[54]; // @[wallace.scala 69:18]
  assign FullAdder_363_io_b = io_pp_26[53]; // @[wallace.scala 70:18]
  assign FullAdder_363_io_ci = io_pp_27[52]; // @[wallace.scala 71:19]
  assign FullAdder_364_io_a = io_pp_28[51]; // @[wallace.scala 69:18]
  assign FullAdder_364_io_b = io_pp_29[50]; // @[wallace.scala 70:18]
  assign FullAdder_364_io_ci = io_pp_30[49]; // @[wallace.scala 71:19]
  assign FullAdder_365_io_a = io_pp_31[48]; // @[wallace.scala 69:18]
  assign FullAdder_365_io_b = io_pp_32[47]; // @[wallace.scala 70:18]
  assign FullAdder_365_io_ci = io_pp_33[46]; // @[wallace.scala 71:19]
  assign FullAdder_366_io_a = io_pp_34[45]; // @[wallace.scala 69:18]
  assign FullAdder_366_io_b = io_pp_35[44]; // @[wallace.scala 70:18]
  assign FullAdder_366_io_ci = io_pp_36[43]; // @[wallace.scala 71:19]
  assign FullAdder_367_io_a = io_pp_37[42]; // @[wallace.scala 69:18]
  assign FullAdder_367_io_b = io_pp_38[41]; // @[wallace.scala 70:18]
  assign FullAdder_367_io_ci = io_pp_39[40]; // @[wallace.scala 71:19]
  assign FullAdder_368_io_a = io_pp_40[39]; // @[wallace.scala 69:18]
  assign FullAdder_368_io_b = io_pp_41[38]; // @[wallace.scala 70:18]
  assign FullAdder_368_io_ci = io_pp_42[37]; // @[wallace.scala 71:19]
  assign FullAdder_369_io_a = io_pp_43[36]; // @[wallace.scala 69:18]
  assign FullAdder_369_io_b = io_pp_44[35]; // @[wallace.scala 70:18]
  assign FullAdder_369_io_ci = io_pp_45[34]; // @[wallace.scala 71:19]
  assign FullAdder_370_io_a = io_pp_46[33]; // @[wallace.scala 69:18]
  assign FullAdder_370_io_b = io_pp_47[32]; // @[wallace.scala 70:18]
  assign FullAdder_370_io_ci = io_pp_48[31]; // @[wallace.scala 71:19]
  assign FullAdder_371_io_a = io_pp_49[30]; // @[wallace.scala 69:18]
  assign FullAdder_371_io_b = io_pp_50[29]; // @[wallace.scala 70:18]
  assign FullAdder_371_io_ci = io_pp_51[28]; // @[wallace.scala 71:19]
  assign FullAdder_372_io_a = io_pp_52[27]; // @[wallace.scala 69:18]
  assign FullAdder_372_io_b = io_pp_53[26]; // @[wallace.scala 70:18]
  assign FullAdder_372_io_ci = io_pp_54[25]; // @[wallace.scala 71:19]
  assign FullAdder_373_io_a = io_pp_55[24]; // @[wallace.scala 69:18]
  assign FullAdder_373_io_b = io_pp_56[23]; // @[wallace.scala 70:18]
  assign FullAdder_373_io_ci = io_pp_57[22]; // @[wallace.scala 71:19]
  assign FullAdder_374_io_a = io_pp_58[21]; // @[wallace.scala 69:18]
  assign FullAdder_374_io_b = io_pp_59[20]; // @[wallace.scala 70:18]
  assign FullAdder_374_io_ci = io_pp_60[19]; // @[wallace.scala 71:19]
  assign FullAdder_375_io_a = io_pp_61[18]; // @[wallace.scala 69:18]
  assign FullAdder_375_io_b = io_pp_62[17]; // @[wallace.scala 70:18]
  assign FullAdder_375_io_ci = io_pp_63[16]; // @[wallace.scala 71:19]
  assign FullAdder_376_io_a = io_pp_15[63]; // @[wallace.scala 69:18]
  assign FullAdder_376_io_b = io_pp_16[62]; // @[wallace.scala 70:18]
  assign FullAdder_376_io_ci = io_pp_17[61]; // @[wallace.scala 71:19]
  assign FullAdder_377_io_a = io_pp_18[60]; // @[wallace.scala 69:18]
  assign FullAdder_377_io_b = io_pp_19[59]; // @[wallace.scala 70:18]
  assign FullAdder_377_io_ci = io_pp_20[58]; // @[wallace.scala 71:19]
  assign FullAdder_378_io_a = io_pp_21[57]; // @[wallace.scala 69:18]
  assign FullAdder_378_io_b = io_pp_22[56]; // @[wallace.scala 70:18]
  assign FullAdder_378_io_ci = io_pp_23[55]; // @[wallace.scala 71:19]
  assign FullAdder_379_io_a = io_pp_24[54]; // @[wallace.scala 69:18]
  assign FullAdder_379_io_b = io_pp_25[53]; // @[wallace.scala 70:18]
  assign FullAdder_379_io_ci = io_pp_26[52]; // @[wallace.scala 71:19]
  assign FullAdder_380_io_a = io_pp_27[51]; // @[wallace.scala 69:18]
  assign FullAdder_380_io_b = io_pp_28[50]; // @[wallace.scala 70:18]
  assign FullAdder_380_io_ci = io_pp_29[49]; // @[wallace.scala 71:19]
  assign FullAdder_381_io_a = io_pp_30[48]; // @[wallace.scala 69:18]
  assign FullAdder_381_io_b = io_pp_31[47]; // @[wallace.scala 70:18]
  assign FullAdder_381_io_ci = io_pp_32[46]; // @[wallace.scala 71:19]
  assign FullAdder_382_io_a = io_pp_33[45]; // @[wallace.scala 69:18]
  assign FullAdder_382_io_b = io_pp_34[44]; // @[wallace.scala 70:18]
  assign FullAdder_382_io_ci = io_pp_35[43]; // @[wallace.scala 71:19]
  assign FullAdder_383_io_a = io_pp_36[42]; // @[wallace.scala 69:18]
  assign FullAdder_383_io_b = io_pp_37[41]; // @[wallace.scala 70:18]
  assign FullAdder_383_io_ci = io_pp_38[40]; // @[wallace.scala 71:19]
  assign FullAdder_384_io_a = io_pp_39[39]; // @[wallace.scala 69:18]
  assign FullAdder_384_io_b = io_pp_40[38]; // @[wallace.scala 70:18]
  assign FullAdder_384_io_ci = io_pp_41[37]; // @[wallace.scala 71:19]
  assign FullAdder_385_io_a = io_pp_42[36]; // @[wallace.scala 69:18]
  assign FullAdder_385_io_b = io_pp_43[35]; // @[wallace.scala 70:18]
  assign FullAdder_385_io_ci = io_pp_44[34]; // @[wallace.scala 71:19]
  assign FullAdder_386_io_a = io_pp_45[33]; // @[wallace.scala 69:18]
  assign FullAdder_386_io_b = io_pp_46[32]; // @[wallace.scala 70:18]
  assign FullAdder_386_io_ci = io_pp_47[31]; // @[wallace.scala 71:19]
  assign FullAdder_387_io_a = io_pp_48[30]; // @[wallace.scala 69:18]
  assign FullAdder_387_io_b = io_pp_49[29]; // @[wallace.scala 70:18]
  assign FullAdder_387_io_ci = io_pp_50[28]; // @[wallace.scala 71:19]
  assign FullAdder_388_io_a = io_pp_51[27]; // @[wallace.scala 69:18]
  assign FullAdder_388_io_b = io_pp_52[26]; // @[wallace.scala 70:18]
  assign FullAdder_388_io_ci = io_pp_53[25]; // @[wallace.scala 71:19]
  assign FullAdder_389_io_a = io_pp_54[24]; // @[wallace.scala 69:18]
  assign FullAdder_389_io_b = io_pp_55[23]; // @[wallace.scala 70:18]
  assign FullAdder_389_io_ci = io_pp_56[22]; // @[wallace.scala 71:19]
  assign FullAdder_390_io_a = io_pp_57[21]; // @[wallace.scala 69:18]
  assign FullAdder_390_io_b = io_pp_58[20]; // @[wallace.scala 70:18]
  assign FullAdder_390_io_ci = io_pp_59[19]; // @[wallace.scala 71:19]
  assign FullAdder_391_io_a = io_pp_60[18]; // @[wallace.scala 69:18]
  assign FullAdder_391_io_b = io_pp_61[17]; // @[wallace.scala 70:18]
  assign FullAdder_391_io_ci = io_pp_62[16]; // @[wallace.scala 71:19]
  assign FullAdder_392_io_a = io_pp_14[63]; // @[wallace.scala 69:18]
  assign FullAdder_392_io_b = io_pp_15[62]; // @[wallace.scala 70:18]
  assign FullAdder_392_io_ci = io_pp_16[61]; // @[wallace.scala 71:19]
  assign FullAdder_393_io_a = io_pp_17[60]; // @[wallace.scala 69:18]
  assign FullAdder_393_io_b = io_pp_18[59]; // @[wallace.scala 70:18]
  assign FullAdder_393_io_ci = io_pp_19[58]; // @[wallace.scala 71:19]
  assign FullAdder_394_io_a = io_pp_20[57]; // @[wallace.scala 69:18]
  assign FullAdder_394_io_b = io_pp_21[56]; // @[wallace.scala 70:18]
  assign FullAdder_394_io_ci = io_pp_22[55]; // @[wallace.scala 71:19]
  assign FullAdder_395_io_a = io_pp_23[54]; // @[wallace.scala 69:18]
  assign FullAdder_395_io_b = io_pp_24[53]; // @[wallace.scala 70:18]
  assign FullAdder_395_io_ci = io_pp_25[52]; // @[wallace.scala 71:19]
  assign FullAdder_396_io_a = io_pp_26[51]; // @[wallace.scala 69:18]
  assign FullAdder_396_io_b = io_pp_27[50]; // @[wallace.scala 70:18]
  assign FullAdder_396_io_ci = io_pp_28[49]; // @[wallace.scala 71:19]
  assign FullAdder_397_io_a = io_pp_29[48]; // @[wallace.scala 69:18]
  assign FullAdder_397_io_b = io_pp_30[47]; // @[wallace.scala 70:18]
  assign FullAdder_397_io_ci = io_pp_31[46]; // @[wallace.scala 71:19]
  assign FullAdder_398_io_a = io_pp_32[45]; // @[wallace.scala 69:18]
  assign FullAdder_398_io_b = io_pp_33[44]; // @[wallace.scala 70:18]
  assign FullAdder_398_io_ci = io_pp_34[43]; // @[wallace.scala 71:19]
  assign FullAdder_399_io_a = io_pp_35[42]; // @[wallace.scala 69:18]
  assign FullAdder_399_io_b = io_pp_36[41]; // @[wallace.scala 70:18]
  assign FullAdder_399_io_ci = io_pp_37[40]; // @[wallace.scala 71:19]
  assign FullAdder_400_io_a = io_pp_38[39]; // @[wallace.scala 69:18]
  assign FullAdder_400_io_b = io_pp_39[38]; // @[wallace.scala 70:18]
  assign FullAdder_400_io_ci = io_pp_40[37]; // @[wallace.scala 71:19]
  assign FullAdder_401_io_a = io_pp_41[36]; // @[wallace.scala 69:18]
  assign FullAdder_401_io_b = io_pp_42[35]; // @[wallace.scala 70:18]
  assign FullAdder_401_io_ci = io_pp_43[34]; // @[wallace.scala 71:19]
  assign FullAdder_402_io_a = io_pp_44[33]; // @[wallace.scala 69:18]
  assign FullAdder_402_io_b = io_pp_45[32]; // @[wallace.scala 70:18]
  assign FullAdder_402_io_ci = io_pp_46[31]; // @[wallace.scala 71:19]
  assign FullAdder_403_io_a = io_pp_47[30]; // @[wallace.scala 69:18]
  assign FullAdder_403_io_b = io_pp_48[29]; // @[wallace.scala 70:18]
  assign FullAdder_403_io_ci = io_pp_49[28]; // @[wallace.scala 71:19]
  assign FullAdder_404_io_a = io_pp_50[27]; // @[wallace.scala 69:18]
  assign FullAdder_404_io_b = io_pp_51[26]; // @[wallace.scala 70:18]
  assign FullAdder_404_io_ci = io_pp_52[25]; // @[wallace.scala 71:19]
  assign FullAdder_405_io_a = io_pp_53[24]; // @[wallace.scala 69:18]
  assign FullAdder_405_io_b = io_pp_54[23]; // @[wallace.scala 70:18]
  assign FullAdder_405_io_ci = io_pp_55[22]; // @[wallace.scala 71:19]
  assign FullAdder_406_io_a = io_pp_56[21]; // @[wallace.scala 69:18]
  assign FullAdder_406_io_b = io_pp_57[20]; // @[wallace.scala 70:18]
  assign FullAdder_406_io_ci = io_pp_58[19]; // @[wallace.scala 71:19]
  assign FullAdder_407_io_a = io_pp_59[18]; // @[wallace.scala 69:18]
  assign FullAdder_407_io_b = io_pp_60[17]; // @[wallace.scala 70:18]
  assign FullAdder_407_io_ci = io_pp_61[16]; // @[wallace.scala 71:19]
  assign HalfAdder_13_io_a = io_pp_62[15]; // @[wallace.scala 59:18]
  assign HalfAdder_13_io_b = io_pp_63[14]; // @[wallace.scala 60:18]
  assign FullAdder_408_io_a = io_pp_13[63]; // @[wallace.scala 69:18]
  assign FullAdder_408_io_b = io_pp_14[62]; // @[wallace.scala 70:18]
  assign FullAdder_408_io_ci = io_pp_15[61]; // @[wallace.scala 71:19]
  assign FullAdder_409_io_a = io_pp_16[60]; // @[wallace.scala 69:18]
  assign FullAdder_409_io_b = io_pp_17[59]; // @[wallace.scala 70:18]
  assign FullAdder_409_io_ci = io_pp_18[58]; // @[wallace.scala 71:19]
  assign FullAdder_410_io_a = io_pp_19[57]; // @[wallace.scala 69:18]
  assign FullAdder_410_io_b = io_pp_20[56]; // @[wallace.scala 70:18]
  assign FullAdder_410_io_ci = io_pp_21[55]; // @[wallace.scala 71:19]
  assign FullAdder_411_io_a = io_pp_22[54]; // @[wallace.scala 69:18]
  assign FullAdder_411_io_b = io_pp_23[53]; // @[wallace.scala 70:18]
  assign FullAdder_411_io_ci = io_pp_24[52]; // @[wallace.scala 71:19]
  assign FullAdder_412_io_a = io_pp_25[51]; // @[wallace.scala 69:18]
  assign FullAdder_412_io_b = io_pp_26[50]; // @[wallace.scala 70:18]
  assign FullAdder_412_io_ci = io_pp_27[49]; // @[wallace.scala 71:19]
  assign FullAdder_413_io_a = io_pp_28[48]; // @[wallace.scala 69:18]
  assign FullAdder_413_io_b = io_pp_29[47]; // @[wallace.scala 70:18]
  assign FullAdder_413_io_ci = io_pp_30[46]; // @[wallace.scala 71:19]
  assign FullAdder_414_io_a = io_pp_31[45]; // @[wallace.scala 69:18]
  assign FullAdder_414_io_b = io_pp_32[44]; // @[wallace.scala 70:18]
  assign FullAdder_414_io_ci = io_pp_33[43]; // @[wallace.scala 71:19]
  assign FullAdder_415_io_a = io_pp_34[42]; // @[wallace.scala 69:18]
  assign FullAdder_415_io_b = io_pp_35[41]; // @[wallace.scala 70:18]
  assign FullAdder_415_io_ci = io_pp_36[40]; // @[wallace.scala 71:19]
  assign FullAdder_416_io_a = io_pp_37[39]; // @[wallace.scala 69:18]
  assign FullAdder_416_io_b = io_pp_38[38]; // @[wallace.scala 70:18]
  assign FullAdder_416_io_ci = io_pp_39[37]; // @[wallace.scala 71:19]
  assign FullAdder_417_io_a = io_pp_40[36]; // @[wallace.scala 69:18]
  assign FullAdder_417_io_b = io_pp_41[35]; // @[wallace.scala 70:18]
  assign FullAdder_417_io_ci = io_pp_42[34]; // @[wallace.scala 71:19]
  assign FullAdder_418_io_a = io_pp_43[33]; // @[wallace.scala 69:18]
  assign FullAdder_418_io_b = io_pp_44[32]; // @[wallace.scala 70:18]
  assign FullAdder_418_io_ci = io_pp_45[31]; // @[wallace.scala 71:19]
  assign FullAdder_419_io_a = io_pp_46[30]; // @[wallace.scala 69:18]
  assign FullAdder_419_io_b = io_pp_47[29]; // @[wallace.scala 70:18]
  assign FullAdder_419_io_ci = io_pp_48[28]; // @[wallace.scala 71:19]
  assign FullAdder_420_io_a = io_pp_49[27]; // @[wallace.scala 69:18]
  assign FullAdder_420_io_b = io_pp_50[26]; // @[wallace.scala 70:18]
  assign FullAdder_420_io_ci = io_pp_51[25]; // @[wallace.scala 71:19]
  assign FullAdder_421_io_a = io_pp_52[24]; // @[wallace.scala 69:18]
  assign FullAdder_421_io_b = io_pp_53[23]; // @[wallace.scala 70:18]
  assign FullAdder_421_io_ci = io_pp_54[22]; // @[wallace.scala 71:19]
  assign FullAdder_422_io_a = io_pp_55[21]; // @[wallace.scala 69:18]
  assign FullAdder_422_io_b = io_pp_56[20]; // @[wallace.scala 70:18]
  assign FullAdder_422_io_ci = io_pp_57[19]; // @[wallace.scala 71:19]
  assign FullAdder_423_io_a = io_pp_58[18]; // @[wallace.scala 69:18]
  assign FullAdder_423_io_b = io_pp_59[17]; // @[wallace.scala 70:18]
  assign FullAdder_423_io_ci = io_pp_60[16]; // @[wallace.scala 71:19]
  assign FullAdder_424_io_a = io_pp_61[15]; // @[wallace.scala 69:18]
  assign FullAdder_424_io_b = io_pp_62[14]; // @[wallace.scala 70:18]
  assign FullAdder_424_io_ci = io_pp_63[13]; // @[wallace.scala 71:19]
  assign FullAdder_425_io_a = io_pp_12[63]; // @[wallace.scala 69:18]
  assign FullAdder_425_io_b = io_pp_13[62]; // @[wallace.scala 70:18]
  assign FullAdder_425_io_ci = io_pp_14[61]; // @[wallace.scala 71:19]
  assign FullAdder_426_io_a = io_pp_15[60]; // @[wallace.scala 69:18]
  assign FullAdder_426_io_b = io_pp_16[59]; // @[wallace.scala 70:18]
  assign FullAdder_426_io_ci = io_pp_17[58]; // @[wallace.scala 71:19]
  assign FullAdder_427_io_a = io_pp_18[57]; // @[wallace.scala 69:18]
  assign FullAdder_427_io_b = io_pp_19[56]; // @[wallace.scala 70:18]
  assign FullAdder_427_io_ci = io_pp_20[55]; // @[wallace.scala 71:19]
  assign FullAdder_428_io_a = io_pp_21[54]; // @[wallace.scala 69:18]
  assign FullAdder_428_io_b = io_pp_22[53]; // @[wallace.scala 70:18]
  assign FullAdder_428_io_ci = io_pp_23[52]; // @[wallace.scala 71:19]
  assign FullAdder_429_io_a = io_pp_24[51]; // @[wallace.scala 69:18]
  assign FullAdder_429_io_b = io_pp_25[50]; // @[wallace.scala 70:18]
  assign FullAdder_429_io_ci = io_pp_26[49]; // @[wallace.scala 71:19]
  assign FullAdder_430_io_a = io_pp_27[48]; // @[wallace.scala 69:18]
  assign FullAdder_430_io_b = io_pp_28[47]; // @[wallace.scala 70:18]
  assign FullAdder_430_io_ci = io_pp_29[46]; // @[wallace.scala 71:19]
  assign FullAdder_431_io_a = io_pp_30[45]; // @[wallace.scala 69:18]
  assign FullAdder_431_io_b = io_pp_31[44]; // @[wallace.scala 70:18]
  assign FullAdder_431_io_ci = io_pp_32[43]; // @[wallace.scala 71:19]
  assign FullAdder_432_io_a = io_pp_33[42]; // @[wallace.scala 69:18]
  assign FullAdder_432_io_b = io_pp_34[41]; // @[wallace.scala 70:18]
  assign FullAdder_432_io_ci = io_pp_35[40]; // @[wallace.scala 71:19]
  assign FullAdder_433_io_a = io_pp_36[39]; // @[wallace.scala 69:18]
  assign FullAdder_433_io_b = io_pp_37[38]; // @[wallace.scala 70:18]
  assign FullAdder_433_io_ci = io_pp_38[37]; // @[wallace.scala 71:19]
  assign FullAdder_434_io_a = io_pp_39[36]; // @[wallace.scala 69:18]
  assign FullAdder_434_io_b = io_pp_40[35]; // @[wallace.scala 70:18]
  assign FullAdder_434_io_ci = io_pp_41[34]; // @[wallace.scala 71:19]
  assign FullAdder_435_io_a = io_pp_42[33]; // @[wallace.scala 69:18]
  assign FullAdder_435_io_b = io_pp_43[32]; // @[wallace.scala 70:18]
  assign FullAdder_435_io_ci = io_pp_44[31]; // @[wallace.scala 71:19]
  assign FullAdder_436_io_a = io_pp_45[30]; // @[wallace.scala 69:18]
  assign FullAdder_436_io_b = io_pp_46[29]; // @[wallace.scala 70:18]
  assign FullAdder_436_io_ci = io_pp_47[28]; // @[wallace.scala 71:19]
  assign FullAdder_437_io_a = io_pp_48[27]; // @[wallace.scala 69:18]
  assign FullAdder_437_io_b = io_pp_49[26]; // @[wallace.scala 70:18]
  assign FullAdder_437_io_ci = io_pp_50[25]; // @[wallace.scala 71:19]
  assign FullAdder_438_io_a = io_pp_51[24]; // @[wallace.scala 69:18]
  assign FullAdder_438_io_b = io_pp_52[23]; // @[wallace.scala 70:18]
  assign FullAdder_438_io_ci = io_pp_53[22]; // @[wallace.scala 71:19]
  assign FullAdder_439_io_a = io_pp_54[21]; // @[wallace.scala 69:18]
  assign FullAdder_439_io_b = io_pp_55[20]; // @[wallace.scala 70:18]
  assign FullAdder_439_io_ci = io_pp_56[19]; // @[wallace.scala 71:19]
  assign FullAdder_440_io_a = io_pp_57[18]; // @[wallace.scala 69:18]
  assign FullAdder_440_io_b = io_pp_58[17]; // @[wallace.scala 70:18]
  assign FullAdder_440_io_ci = io_pp_59[16]; // @[wallace.scala 71:19]
  assign FullAdder_441_io_a = io_pp_60[15]; // @[wallace.scala 69:18]
  assign FullAdder_441_io_b = io_pp_61[14]; // @[wallace.scala 70:18]
  assign FullAdder_441_io_ci = io_pp_62[13]; // @[wallace.scala 71:19]
  assign FullAdder_442_io_a = io_pp_11[63]; // @[wallace.scala 69:18]
  assign FullAdder_442_io_b = io_pp_12[62]; // @[wallace.scala 70:18]
  assign FullAdder_442_io_ci = io_pp_13[61]; // @[wallace.scala 71:19]
  assign FullAdder_443_io_a = io_pp_14[60]; // @[wallace.scala 69:18]
  assign FullAdder_443_io_b = io_pp_15[59]; // @[wallace.scala 70:18]
  assign FullAdder_443_io_ci = io_pp_16[58]; // @[wallace.scala 71:19]
  assign FullAdder_444_io_a = io_pp_17[57]; // @[wallace.scala 69:18]
  assign FullAdder_444_io_b = io_pp_18[56]; // @[wallace.scala 70:18]
  assign FullAdder_444_io_ci = io_pp_19[55]; // @[wallace.scala 71:19]
  assign FullAdder_445_io_a = io_pp_20[54]; // @[wallace.scala 69:18]
  assign FullAdder_445_io_b = io_pp_21[53]; // @[wallace.scala 70:18]
  assign FullAdder_445_io_ci = io_pp_22[52]; // @[wallace.scala 71:19]
  assign FullAdder_446_io_a = io_pp_23[51]; // @[wallace.scala 69:18]
  assign FullAdder_446_io_b = io_pp_24[50]; // @[wallace.scala 70:18]
  assign FullAdder_446_io_ci = io_pp_25[49]; // @[wallace.scala 71:19]
  assign FullAdder_447_io_a = io_pp_26[48]; // @[wallace.scala 69:18]
  assign FullAdder_447_io_b = io_pp_27[47]; // @[wallace.scala 70:18]
  assign FullAdder_447_io_ci = io_pp_28[46]; // @[wallace.scala 71:19]
  assign FullAdder_448_io_a = io_pp_29[45]; // @[wallace.scala 69:18]
  assign FullAdder_448_io_b = io_pp_30[44]; // @[wallace.scala 70:18]
  assign FullAdder_448_io_ci = io_pp_31[43]; // @[wallace.scala 71:19]
  assign FullAdder_449_io_a = io_pp_32[42]; // @[wallace.scala 69:18]
  assign FullAdder_449_io_b = io_pp_33[41]; // @[wallace.scala 70:18]
  assign FullAdder_449_io_ci = io_pp_34[40]; // @[wallace.scala 71:19]
  assign FullAdder_450_io_a = io_pp_35[39]; // @[wallace.scala 69:18]
  assign FullAdder_450_io_b = io_pp_36[38]; // @[wallace.scala 70:18]
  assign FullAdder_450_io_ci = io_pp_37[37]; // @[wallace.scala 71:19]
  assign FullAdder_451_io_a = io_pp_38[36]; // @[wallace.scala 69:18]
  assign FullAdder_451_io_b = io_pp_39[35]; // @[wallace.scala 70:18]
  assign FullAdder_451_io_ci = io_pp_40[34]; // @[wallace.scala 71:19]
  assign FullAdder_452_io_a = io_pp_41[33]; // @[wallace.scala 69:18]
  assign FullAdder_452_io_b = io_pp_42[32]; // @[wallace.scala 70:18]
  assign FullAdder_452_io_ci = io_pp_43[31]; // @[wallace.scala 71:19]
  assign FullAdder_453_io_a = io_pp_44[30]; // @[wallace.scala 69:18]
  assign FullAdder_453_io_b = io_pp_45[29]; // @[wallace.scala 70:18]
  assign FullAdder_453_io_ci = io_pp_46[28]; // @[wallace.scala 71:19]
  assign FullAdder_454_io_a = io_pp_47[27]; // @[wallace.scala 69:18]
  assign FullAdder_454_io_b = io_pp_48[26]; // @[wallace.scala 70:18]
  assign FullAdder_454_io_ci = io_pp_49[25]; // @[wallace.scala 71:19]
  assign FullAdder_455_io_a = io_pp_50[24]; // @[wallace.scala 69:18]
  assign FullAdder_455_io_b = io_pp_51[23]; // @[wallace.scala 70:18]
  assign FullAdder_455_io_ci = io_pp_52[22]; // @[wallace.scala 71:19]
  assign FullAdder_456_io_a = io_pp_53[21]; // @[wallace.scala 69:18]
  assign FullAdder_456_io_b = io_pp_54[20]; // @[wallace.scala 70:18]
  assign FullAdder_456_io_ci = io_pp_55[19]; // @[wallace.scala 71:19]
  assign FullAdder_457_io_a = io_pp_56[18]; // @[wallace.scala 69:18]
  assign FullAdder_457_io_b = io_pp_57[17]; // @[wallace.scala 70:18]
  assign FullAdder_457_io_ci = io_pp_58[16]; // @[wallace.scala 71:19]
  assign FullAdder_458_io_a = io_pp_59[15]; // @[wallace.scala 69:18]
  assign FullAdder_458_io_b = io_pp_60[14]; // @[wallace.scala 70:18]
  assign FullAdder_458_io_ci = io_pp_61[13]; // @[wallace.scala 71:19]
  assign HalfAdder_14_io_a = io_pp_62[12]; // @[wallace.scala 59:18]
  assign HalfAdder_14_io_b = io_pp_63[11]; // @[wallace.scala 60:18]
  assign FullAdder_459_io_a = io_pp_10[63]; // @[wallace.scala 69:18]
  assign FullAdder_459_io_b = io_pp_11[62]; // @[wallace.scala 70:18]
  assign FullAdder_459_io_ci = io_pp_12[61]; // @[wallace.scala 71:19]
  assign FullAdder_460_io_a = io_pp_13[60]; // @[wallace.scala 69:18]
  assign FullAdder_460_io_b = io_pp_14[59]; // @[wallace.scala 70:18]
  assign FullAdder_460_io_ci = io_pp_15[58]; // @[wallace.scala 71:19]
  assign FullAdder_461_io_a = io_pp_16[57]; // @[wallace.scala 69:18]
  assign FullAdder_461_io_b = io_pp_17[56]; // @[wallace.scala 70:18]
  assign FullAdder_461_io_ci = io_pp_18[55]; // @[wallace.scala 71:19]
  assign FullAdder_462_io_a = io_pp_19[54]; // @[wallace.scala 69:18]
  assign FullAdder_462_io_b = io_pp_20[53]; // @[wallace.scala 70:18]
  assign FullAdder_462_io_ci = io_pp_21[52]; // @[wallace.scala 71:19]
  assign FullAdder_463_io_a = io_pp_22[51]; // @[wallace.scala 69:18]
  assign FullAdder_463_io_b = io_pp_23[50]; // @[wallace.scala 70:18]
  assign FullAdder_463_io_ci = io_pp_24[49]; // @[wallace.scala 71:19]
  assign FullAdder_464_io_a = io_pp_25[48]; // @[wallace.scala 69:18]
  assign FullAdder_464_io_b = io_pp_26[47]; // @[wallace.scala 70:18]
  assign FullAdder_464_io_ci = io_pp_27[46]; // @[wallace.scala 71:19]
  assign FullAdder_465_io_a = io_pp_28[45]; // @[wallace.scala 69:18]
  assign FullAdder_465_io_b = io_pp_29[44]; // @[wallace.scala 70:18]
  assign FullAdder_465_io_ci = io_pp_30[43]; // @[wallace.scala 71:19]
  assign FullAdder_466_io_a = io_pp_31[42]; // @[wallace.scala 69:18]
  assign FullAdder_466_io_b = io_pp_32[41]; // @[wallace.scala 70:18]
  assign FullAdder_466_io_ci = io_pp_33[40]; // @[wallace.scala 71:19]
  assign FullAdder_467_io_a = io_pp_34[39]; // @[wallace.scala 69:18]
  assign FullAdder_467_io_b = io_pp_35[38]; // @[wallace.scala 70:18]
  assign FullAdder_467_io_ci = io_pp_36[37]; // @[wallace.scala 71:19]
  assign FullAdder_468_io_a = io_pp_37[36]; // @[wallace.scala 69:18]
  assign FullAdder_468_io_b = io_pp_38[35]; // @[wallace.scala 70:18]
  assign FullAdder_468_io_ci = io_pp_39[34]; // @[wallace.scala 71:19]
  assign FullAdder_469_io_a = io_pp_40[33]; // @[wallace.scala 69:18]
  assign FullAdder_469_io_b = io_pp_41[32]; // @[wallace.scala 70:18]
  assign FullAdder_469_io_ci = io_pp_42[31]; // @[wallace.scala 71:19]
  assign FullAdder_470_io_a = io_pp_43[30]; // @[wallace.scala 69:18]
  assign FullAdder_470_io_b = io_pp_44[29]; // @[wallace.scala 70:18]
  assign FullAdder_470_io_ci = io_pp_45[28]; // @[wallace.scala 71:19]
  assign FullAdder_471_io_a = io_pp_46[27]; // @[wallace.scala 69:18]
  assign FullAdder_471_io_b = io_pp_47[26]; // @[wallace.scala 70:18]
  assign FullAdder_471_io_ci = io_pp_48[25]; // @[wallace.scala 71:19]
  assign FullAdder_472_io_a = io_pp_49[24]; // @[wallace.scala 69:18]
  assign FullAdder_472_io_b = io_pp_50[23]; // @[wallace.scala 70:18]
  assign FullAdder_472_io_ci = io_pp_51[22]; // @[wallace.scala 71:19]
  assign FullAdder_473_io_a = io_pp_52[21]; // @[wallace.scala 69:18]
  assign FullAdder_473_io_b = io_pp_53[20]; // @[wallace.scala 70:18]
  assign FullAdder_473_io_ci = io_pp_54[19]; // @[wallace.scala 71:19]
  assign FullAdder_474_io_a = io_pp_55[18]; // @[wallace.scala 69:18]
  assign FullAdder_474_io_b = io_pp_56[17]; // @[wallace.scala 70:18]
  assign FullAdder_474_io_ci = io_pp_57[16]; // @[wallace.scala 71:19]
  assign FullAdder_475_io_a = io_pp_58[15]; // @[wallace.scala 69:18]
  assign FullAdder_475_io_b = io_pp_59[14]; // @[wallace.scala 70:18]
  assign FullAdder_475_io_ci = io_pp_60[13]; // @[wallace.scala 71:19]
  assign FullAdder_476_io_a = io_pp_61[12]; // @[wallace.scala 69:18]
  assign FullAdder_476_io_b = io_pp_62[11]; // @[wallace.scala 70:18]
  assign FullAdder_476_io_ci = io_pp_63[10]; // @[wallace.scala 71:19]
  assign FullAdder_477_io_a = io_pp_9[63]; // @[wallace.scala 69:18]
  assign FullAdder_477_io_b = io_pp_10[62]; // @[wallace.scala 70:18]
  assign FullAdder_477_io_ci = io_pp_11[61]; // @[wallace.scala 71:19]
  assign FullAdder_478_io_a = io_pp_12[60]; // @[wallace.scala 69:18]
  assign FullAdder_478_io_b = io_pp_13[59]; // @[wallace.scala 70:18]
  assign FullAdder_478_io_ci = io_pp_14[58]; // @[wallace.scala 71:19]
  assign FullAdder_479_io_a = io_pp_15[57]; // @[wallace.scala 69:18]
  assign FullAdder_479_io_b = io_pp_16[56]; // @[wallace.scala 70:18]
  assign FullAdder_479_io_ci = io_pp_17[55]; // @[wallace.scala 71:19]
  assign FullAdder_480_io_a = io_pp_18[54]; // @[wallace.scala 69:18]
  assign FullAdder_480_io_b = io_pp_19[53]; // @[wallace.scala 70:18]
  assign FullAdder_480_io_ci = io_pp_20[52]; // @[wallace.scala 71:19]
  assign FullAdder_481_io_a = io_pp_21[51]; // @[wallace.scala 69:18]
  assign FullAdder_481_io_b = io_pp_22[50]; // @[wallace.scala 70:18]
  assign FullAdder_481_io_ci = io_pp_23[49]; // @[wallace.scala 71:19]
  assign FullAdder_482_io_a = io_pp_24[48]; // @[wallace.scala 69:18]
  assign FullAdder_482_io_b = io_pp_25[47]; // @[wallace.scala 70:18]
  assign FullAdder_482_io_ci = io_pp_26[46]; // @[wallace.scala 71:19]
  assign FullAdder_483_io_a = io_pp_27[45]; // @[wallace.scala 69:18]
  assign FullAdder_483_io_b = io_pp_28[44]; // @[wallace.scala 70:18]
  assign FullAdder_483_io_ci = io_pp_29[43]; // @[wallace.scala 71:19]
  assign FullAdder_484_io_a = io_pp_30[42]; // @[wallace.scala 69:18]
  assign FullAdder_484_io_b = io_pp_31[41]; // @[wallace.scala 70:18]
  assign FullAdder_484_io_ci = io_pp_32[40]; // @[wallace.scala 71:19]
  assign FullAdder_485_io_a = io_pp_33[39]; // @[wallace.scala 69:18]
  assign FullAdder_485_io_b = io_pp_34[38]; // @[wallace.scala 70:18]
  assign FullAdder_485_io_ci = io_pp_35[37]; // @[wallace.scala 71:19]
  assign FullAdder_486_io_a = io_pp_36[36]; // @[wallace.scala 69:18]
  assign FullAdder_486_io_b = io_pp_37[35]; // @[wallace.scala 70:18]
  assign FullAdder_486_io_ci = io_pp_38[34]; // @[wallace.scala 71:19]
  assign FullAdder_487_io_a = io_pp_39[33]; // @[wallace.scala 69:18]
  assign FullAdder_487_io_b = io_pp_40[32]; // @[wallace.scala 70:18]
  assign FullAdder_487_io_ci = io_pp_41[31]; // @[wallace.scala 71:19]
  assign FullAdder_488_io_a = io_pp_42[30]; // @[wallace.scala 69:18]
  assign FullAdder_488_io_b = io_pp_43[29]; // @[wallace.scala 70:18]
  assign FullAdder_488_io_ci = io_pp_44[28]; // @[wallace.scala 71:19]
  assign FullAdder_489_io_a = io_pp_45[27]; // @[wallace.scala 69:18]
  assign FullAdder_489_io_b = io_pp_46[26]; // @[wallace.scala 70:18]
  assign FullAdder_489_io_ci = io_pp_47[25]; // @[wallace.scala 71:19]
  assign FullAdder_490_io_a = io_pp_48[24]; // @[wallace.scala 69:18]
  assign FullAdder_490_io_b = io_pp_49[23]; // @[wallace.scala 70:18]
  assign FullAdder_490_io_ci = io_pp_50[22]; // @[wallace.scala 71:19]
  assign FullAdder_491_io_a = io_pp_51[21]; // @[wallace.scala 69:18]
  assign FullAdder_491_io_b = io_pp_52[20]; // @[wallace.scala 70:18]
  assign FullAdder_491_io_ci = io_pp_53[19]; // @[wallace.scala 71:19]
  assign FullAdder_492_io_a = io_pp_54[18]; // @[wallace.scala 69:18]
  assign FullAdder_492_io_b = io_pp_55[17]; // @[wallace.scala 70:18]
  assign FullAdder_492_io_ci = io_pp_56[16]; // @[wallace.scala 71:19]
  assign FullAdder_493_io_a = io_pp_57[15]; // @[wallace.scala 69:18]
  assign FullAdder_493_io_b = io_pp_58[14]; // @[wallace.scala 70:18]
  assign FullAdder_493_io_ci = io_pp_59[13]; // @[wallace.scala 71:19]
  assign FullAdder_494_io_a = io_pp_60[12]; // @[wallace.scala 69:18]
  assign FullAdder_494_io_b = io_pp_61[11]; // @[wallace.scala 70:18]
  assign FullAdder_494_io_ci = io_pp_62[10]; // @[wallace.scala 71:19]
  assign FullAdder_495_io_a = io_pp_8[63]; // @[wallace.scala 69:18]
  assign FullAdder_495_io_b = io_pp_9[62]; // @[wallace.scala 70:18]
  assign FullAdder_495_io_ci = io_pp_10[61]; // @[wallace.scala 71:19]
  assign FullAdder_496_io_a = io_pp_11[60]; // @[wallace.scala 69:18]
  assign FullAdder_496_io_b = io_pp_12[59]; // @[wallace.scala 70:18]
  assign FullAdder_496_io_ci = io_pp_13[58]; // @[wallace.scala 71:19]
  assign FullAdder_497_io_a = io_pp_14[57]; // @[wallace.scala 69:18]
  assign FullAdder_497_io_b = io_pp_15[56]; // @[wallace.scala 70:18]
  assign FullAdder_497_io_ci = io_pp_16[55]; // @[wallace.scala 71:19]
  assign FullAdder_498_io_a = io_pp_17[54]; // @[wallace.scala 69:18]
  assign FullAdder_498_io_b = io_pp_18[53]; // @[wallace.scala 70:18]
  assign FullAdder_498_io_ci = io_pp_19[52]; // @[wallace.scala 71:19]
  assign FullAdder_499_io_a = io_pp_20[51]; // @[wallace.scala 69:18]
  assign FullAdder_499_io_b = io_pp_21[50]; // @[wallace.scala 70:18]
  assign FullAdder_499_io_ci = io_pp_22[49]; // @[wallace.scala 71:19]
  assign FullAdder_500_io_a = io_pp_23[48]; // @[wallace.scala 69:18]
  assign FullAdder_500_io_b = io_pp_24[47]; // @[wallace.scala 70:18]
  assign FullAdder_500_io_ci = io_pp_25[46]; // @[wallace.scala 71:19]
  assign FullAdder_501_io_a = io_pp_26[45]; // @[wallace.scala 69:18]
  assign FullAdder_501_io_b = io_pp_27[44]; // @[wallace.scala 70:18]
  assign FullAdder_501_io_ci = io_pp_28[43]; // @[wallace.scala 71:19]
  assign FullAdder_502_io_a = io_pp_29[42]; // @[wallace.scala 69:18]
  assign FullAdder_502_io_b = io_pp_30[41]; // @[wallace.scala 70:18]
  assign FullAdder_502_io_ci = io_pp_31[40]; // @[wallace.scala 71:19]
  assign FullAdder_503_io_a = io_pp_32[39]; // @[wallace.scala 69:18]
  assign FullAdder_503_io_b = io_pp_33[38]; // @[wallace.scala 70:18]
  assign FullAdder_503_io_ci = io_pp_34[37]; // @[wallace.scala 71:19]
  assign FullAdder_504_io_a = io_pp_35[36]; // @[wallace.scala 69:18]
  assign FullAdder_504_io_b = io_pp_36[35]; // @[wallace.scala 70:18]
  assign FullAdder_504_io_ci = io_pp_37[34]; // @[wallace.scala 71:19]
  assign FullAdder_505_io_a = io_pp_38[33]; // @[wallace.scala 69:18]
  assign FullAdder_505_io_b = io_pp_39[32]; // @[wallace.scala 70:18]
  assign FullAdder_505_io_ci = io_pp_40[31]; // @[wallace.scala 71:19]
  assign FullAdder_506_io_a = io_pp_41[30]; // @[wallace.scala 69:18]
  assign FullAdder_506_io_b = io_pp_42[29]; // @[wallace.scala 70:18]
  assign FullAdder_506_io_ci = io_pp_43[28]; // @[wallace.scala 71:19]
  assign FullAdder_507_io_a = io_pp_44[27]; // @[wallace.scala 69:18]
  assign FullAdder_507_io_b = io_pp_45[26]; // @[wallace.scala 70:18]
  assign FullAdder_507_io_ci = io_pp_46[25]; // @[wallace.scala 71:19]
  assign FullAdder_508_io_a = io_pp_47[24]; // @[wallace.scala 69:18]
  assign FullAdder_508_io_b = io_pp_48[23]; // @[wallace.scala 70:18]
  assign FullAdder_508_io_ci = io_pp_49[22]; // @[wallace.scala 71:19]
  assign FullAdder_509_io_a = io_pp_50[21]; // @[wallace.scala 69:18]
  assign FullAdder_509_io_b = io_pp_51[20]; // @[wallace.scala 70:18]
  assign FullAdder_509_io_ci = io_pp_52[19]; // @[wallace.scala 71:19]
  assign FullAdder_510_io_a = io_pp_53[18]; // @[wallace.scala 69:18]
  assign FullAdder_510_io_b = io_pp_54[17]; // @[wallace.scala 70:18]
  assign FullAdder_510_io_ci = io_pp_55[16]; // @[wallace.scala 71:19]
  assign FullAdder_511_io_a = io_pp_56[15]; // @[wallace.scala 69:18]
  assign FullAdder_511_io_b = io_pp_57[14]; // @[wallace.scala 70:18]
  assign FullAdder_511_io_ci = io_pp_58[13]; // @[wallace.scala 71:19]
  assign FullAdder_512_io_a = io_pp_59[12]; // @[wallace.scala 69:18]
  assign FullAdder_512_io_b = io_pp_60[11]; // @[wallace.scala 70:18]
  assign FullAdder_512_io_ci = io_pp_61[10]; // @[wallace.scala 71:19]
  assign HalfAdder_15_io_a = io_pp_62[9]; // @[wallace.scala 59:18]
  assign HalfAdder_15_io_b = io_pp_63[8]; // @[wallace.scala 60:18]
  assign FullAdder_513_io_a = io_pp_7[63]; // @[wallace.scala 69:18]
  assign FullAdder_513_io_b = io_pp_8[62]; // @[wallace.scala 70:18]
  assign FullAdder_513_io_ci = io_pp_9[61]; // @[wallace.scala 71:19]
  assign FullAdder_514_io_a = io_pp_10[60]; // @[wallace.scala 69:18]
  assign FullAdder_514_io_b = io_pp_11[59]; // @[wallace.scala 70:18]
  assign FullAdder_514_io_ci = io_pp_12[58]; // @[wallace.scala 71:19]
  assign FullAdder_515_io_a = io_pp_13[57]; // @[wallace.scala 69:18]
  assign FullAdder_515_io_b = io_pp_14[56]; // @[wallace.scala 70:18]
  assign FullAdder_515_io_ci = io_pp_15[55]; // @[wallace.scala 71:19]
  assign FullAdder_516_io_a = io_pp_16[54]; // @[wallace.scala 69:18]
  assign FullAdder_516_io_b = io_pp_17[53]; // @[wallace.scala 70:18]
  assign FullAdder_516_io_ci = io_pp_18[52]; // @[wallace.scala 71:19]
  assign FullAdder_517_io_a = io_pp_19[51]; // @[wallace.scala 69:18]
  assign FullAdder_517_io_b = io_pp_20[50]; // @[wallace.scala 70:18]
  assign FullAdder_517_io_ci = io_pp_21[49]; // @[wallace.scala 71:19]
  assign FullAdder_518_io_a = io_pp_22[48]; // @[wallace.scala 69:18]
  assign FullAdder_518_io_b = io_pp_23[47]; // @[wallace.scala 70:18]
  assign FullAdder_518_io_ci = io_pp_24[46]; // @[wallace.scala 71:19]
  assign FullAdder_519_io_a = io_pp_25[45]; // @[wallace.scala 69:18]
  assign FullAdder_519_io_b = io_pp_26[44]; // @[wallace.scala 70:18]
  assign FullAdder_519_io_ci = io_pp_27[43]; // @[wallace.scala 71:19]
  assign FullAdder_520_io_a = io_pp_28[42]; // @[wallace.scala 69:18]
  assign FullAdder_520_io_b = io_pp_29[41]; // @[wallace.scala 70:18]
  assign FullAdder_520_io_ci = io_pp_30[40]; // @[wallace.scala 71:19]
  assign FullAdder_521_io_a = io_pp_31[39]; // @[wallace.scala 69:18]
  assign FullAdder_521_io_b = io_pp_32[38]; // @[wallace.scala 70:18]
  assign FullAdder_521_io_ci = io_pp_33[37]; // @[wallace.scala 71:19]
  assign FullAdder_522_io_a = io_pp_34[36]; // @[wallace.scala 69:18]
  assign FullAdder_522_io_b = io_pp_35[35]; // @[wallace.scala 70:18]
  assign FullAdder_522_io_ci = io_pp_36[34]; // @[wallace.scala 71:19]
  assign FullAdder_523_io_a = io_pp_37[33]; // @[wallace.scala 69:18]
  assign FullAdder_523_io_b = io_pp_38[32]; // @[wallace.scala 70:18]
  assign FullAdder_523_io_ci = io_pp_39[31]; // @[wallace.scala 71:19]
  assign FullAdder_524_io_a = io_pp_40[30]; // @[wallace.scala 69:18]
  assign FullAdder_524_io_b = io_pp_41[29]; // @[wallace.scala 70:18]
  assign FullAdder_524_io_ci = io_pp_42[28]; // @[wallace.scala 71:19]
  assign FullAdder_525_io_a = io_pp_43[27]; // @[wallace.scala 69:18]
  assign FullAdder_525_io_b = io_pp_44[26]; // @[wallace.scala 70:18]
  assign FullAdder_525_io_ci = io_pp_45[25]; // @[wallace.scala 71:19]
  assign FullAdder_526_io_a = io_pp_46[24]; // @[wallace.scala 69:18]
  assign FullAdder_526_io_b = io_pp_47[23]; // @[wallace.scala 70:18]
  assign FullAdder_526_io_ci = io_pp_48[22]; // @[wallace.scala 71:19]
  assign FullAdder_527_io_a = io_pp_49[21]; // @[wallace.scala 69:18]
  assign FullAdder_527_io_b = io_pp_50[20]; // @[wallace.scala 70:18]
  assign FullAdder_527_io_ci = io_pp_51[19]; // @[wallace.scala 71:19]
  assign FullAdder_528_io_a = io_pp_52[18]; // @[wallace.scala 69:18]
  assign FullAdder_528_io_b = io_pp_53[17]; // @[wallace.scala 70:18]
  assign FullAdder_528_io_ci = io_pp_54[16]; // @[wallace.scala 71:19]
  assign FullAdder_529_io_a = io_pp_55[15]; // @[wallace.scala 69:18]
  assign FullAdder_529_io_b = io_pp_56[14]; // @[wallace.scala 70:18]
  assign FullAdder_529_io_ci = io_pp_57[13]; // @[wallace.scala 71:19]
  assign FullAdder_530_io_a = io_pp_58[12]; // @[wallace.scala 69:18]
  assign FullAdder_530_io_b = io_pp_59[11]; // @[wallace.scala 70:18]
  assign FullAdder_530_io_ci = io_pp_60[10]; // @[wallace.scala 71:19]
  assign FullAdder_531_io_a = io_pp_61[9]; // @[wallace.scala 69:18]
  assign FullAdder_531_io_b = io_pp_62[8]; // @[wallace.scala 70:18]
  assign FullAdder_531_io_ci = io_pp_63[7]; // @[wallace.scala 71:19]
  assign FullAdder_532_io_a = io_pp_6[63]; // @[wallace.scala 69:18]
  assign FullAdder_532_io_b = io_pp_7[62]; // @[wallace.scala 70:18]
  assign FullAdder_532_io_ci = io_pp_8[61]; // @[wallace.scala 71:19]
  assign FullAdder_533_io_a = io_pp_9[60]; // @[wallace.scala 69:18]
  assign FullAdder_533_io_b = io_pp_10[59]; // @[wallace.scala 70:18]
  assign FullAdder_533_io_ci = io_pp_11[58]; // @[wallace.scala 71:19]
  assign FullAdder_534_io_a = io_pp_12[57]; // @[wallace.scala 69:18]
  assign FullAdder_534_io_b = io_pp_13[56]; // @[wallace.scala 70:18]
  assign FullAdder_534_io_ci = io_pp_14[55]; // @[wallace.scala 71:19]
  assign FullAdder_535_io_a = io_pp_15[54]; // @[wallace.scala 69:18]
  assign FullAdder_535_io_b = io_pp_16[53]; // @[wallace.scala 70:18]
  assign FullAdder_535_io_ci = io_pp_17[52]; // @[wallace.scala 71:19]
  assign FullAdder_536_io_a = io_pp_18[51]; // @[wallace.scala 69:18]
  assign FullAdder_536_io_b = io_pp_19[50]; // @[wallace.scala 70:18]
  assign FullAdder_536_io_ci = io_pp_20[49]; // @[wallace.scala 71:19]
  assign FullAdder_537_io_a = io_pp_21[48]; // @[wallace.scala 69:18]
  assign FullAdder_537_io_b = io_pp_22[47]; // @[wallace.scala 70:18]
  assign FullAdder_537_io_ci = io_pp_23[46]; // @[wallace.scala 71:19]
  assign FullAdder_538_io_a = io_pp_24[45]; // @[wallace.scala 69:18]
  assign FullAdder_538_io_b = io_pp_25[44]; // @[wallace.scala 70:18]
  assign FullAdder_538_io_ci = io_pp_26[43]; // @[wallace.scala 71:19]
  assign FullAdder_539_io_a = io_pp_27[42]; // @[wallace.scala 69:18]
  assign FullAdder_539_io_b = io_pp_28[41]; // @[wallace.scala 70:18]
  assign FullAdder_539_io_ci = io_pp_29[40]; // @[wallace.scala 71:19]
  assign FullAdder_540_io_a = io_pp_30[39]; // @[wallace.scala 69:18]
  assign FullAdder_540_io_b = io_pp_31[38]; // @[wallace.scala 70:18]
  assign FullAdder_540_io_ci = io_pp_32[37]; // @[wallace.scala 71:19]
  assign FullAdder_541_io_a = io_pp_33[36]; // @[wallace.scala 69:18]
  assign FullAdder_541_io_b = io_pp_34[35]; // @[wallace.scala 70:18]
  assign FullAdder_541_io_ci = io_pp_35[34]; // @[wallace.scala 71:19]
  assign FullAdder_542_io_a = io_pp_36[33]; // @[wallace.scala 69:18]
  assign FullAdder_542_io_b = io_pp_37[32]; // @[wallace.scala 70:18]
  assign FullAdder_542_io_ci = io_pp_38[31]; // @[wallace.scala 71:19]
  assign FullAdder_543_io_a = io_pp_39[30]; // @[wallace.scala 69:18]
  assign FullAdder_543_io_b = io_pp_40[29]; // @[wallace.scala 70:18]
  assign FullAdder_543_io_ci = io_pp_41[28]; // @[wallace.scala 71:19]
  assign FullAdder_544_io_a = io_pp_42[27]; // @[wallace.scala 69:18]
  assign FullAdder_544_io_b = io_pp_43[26]; // @[wallace.scala 70:18]
  assign FullAdder_544_io_ci = io_pp_44[25]; // @[wallace.scala 71:19]
  assign FullAdder_545_io_a = io_pp_45[24]; // @[wallace.scala 69:18]
  assign FullAdder_545_io_b = io_pp_46[23]; // @[wallace.scala 70:18]
  assign FullAdder_545_io_ci = io_pp_47[22]; // @[wallace.scala 71:19]
  assign FullAdder_546_io_a = io_pp_48[21]; // @[wallace.scala 69:18]
  assign FullAdder_546_io_b = io_pp_49[20]; // @[wallace.scala 70:18]
  assign FullAdder_546_io_ci = io_pp_50[19]; // @[wallace.scala 71:19]
  assign FullAdder_547_io_a = io_pp_51[18]; // @[wallace.scala 69:18]
  assign FullAdder_547_io_b = io_pp_52[17]; // @[wallace.scala 70:18]
  assign FullAdder_547_io_ci = io_pp_53[16]; // @[wallace.scala 71:19]
  assign FullAdder_548_io_a = io_pp_54[15]; // @[wallace.scala 69:18]
  assign FullAdder_548_io_b = io_pp_55[14]; // @[wallace.scala 70:18]
  assign FullAdder_548_io_ci = io_pp_56[13]; // @[wallace.scala 71:19]
  assign FullAdder_549_io_a = io_pp_57[12]; // @[wallace.scala 69:18]
  assign FullAdder_549_io_b = io_pp_58[11]; // @[wallace.scala 70:18]
  assign FullAdder_549_io_ci = io_pp_59[10]; // @[wallace.scala 71:19]
  assign FullAdder_550_io_a = io_pp_60[9]; // @[wallace.scala 69:18]
  assign FullAdder_550_io_b = io_pp_61[8]; // @[wallace.scala 70:18]
  assign FullAdder_550_io_ci = io_pp_62[7]; // @[wallace.scala 71:19]
  assign FullAdder_551_io_a = io_pp_5[63]; // @[wallace.scala 69:18]
  assign FullAdder_551_io_b = io_pp_6[62]; // @[wallace.scala 70:18]
  assign FullAdder_551_io_ci = io_pp_7[61]; // @[wallace.scala 71:19]
  assign FullAdder_552_io_a = io_pp_8[60]; // @[wallace.scala 69:18]
  assign FullAdder_552_io_b = io_pp_9[59]; // @[wallace.scala 70:18]
  assign FullAdder_552_io_ci = io_pp_10[58]; // @[wallace.scala 71:19]
  assign FullAdder_553_io_a = io_pp_11[57]; // @[wallace.scala 69:18]
  assign FullAdder_553_io_b = io_pp_12[56]; // @[wallace.scala 70:18]
  assign FullAdder_553_io_ci = io_pp_13[55]; // @[wallace.scala 71:19]
  assign FullAdder_554_io_a = io_pp_14[54]; // @[wallace.scala 69:18]
  assign FullAdder_554_io_b = io_pp_15[53]; // @[wallace.scala 70:18]
  assign FullAdder_554_io_ci = io_pp_16[52]; // @[wallace.scala 71:19]
  assign FullAdder_555_io_a = io_pp_17[51]; // @[wallace.scala 69:18]
  assign FullAdder_555_io_b = io_pp_18[50]; // @[wallace.scala 70:18]
  assign FullAdder_555_io_ci = io_pp_19[49]; // @[wallace.scala 71:19]
  assign FullAdder_556_io_a = io_pp_20[48]; // @[wallace.scala 69:18]
  assign FullAdder_556_io_b = io_pp_21[47]; // @[wallace.scala 70:18]
  assign FullAdder_556_io_ci = io_pp_22[46]; // @[wallace.scala 71:19]
  assign FullAdder_557_io_a = io_pp_23[45]; // @[wallace.scala 69:18]
  assign FullAdder_557_io_b = io_pp_24[44]; // @[wallace.scala 70:18]
  assign FullAdder_557_io_ci = io_pp_25[43]; // @[wallace.scala 71:19]
  assign FullAdder_558_io_a = io_pp_26[42]; // @[wallace.scala 69:18]
  assign FullAdder_558_io_b = io_pp_27[41]; // @[wallace.scala 70:18]
  assign FullAdder_558_io_ci = io_pp_28[40]; // @[wallace.scala 71:19]
  assign FullAdder_559_io_a = io_pp_29[39]; // @[wallace.scala 69:18]
  assign FullAdder_559_io_b = io_pp_30[38]; // @[wallace.scala 70:18]
  assign FullAdder_559_io_ci = io_pp_31[37]; // @[wallace.scala 71:19]
  assign FullAdder_560_io_a = io_pp_32[36]; // @[wallace.scala 69:18]
  assign FullAdder_560_io_b = io_pp_33[35]; // @[wallace.scala 70:18]
  assign FullAdder_560_io_ci = io_pp_34[34]; // @[wallace.scala 71:19]
  assign FullAdder_561_io_a = io_pp_35[33]; // @[wallace.scala 69:18]
  assign FullAdder_561_io_b = io_pp_36[32]; // @[wallace.scala 70:18]
  assign FullAdder_561_io_ci = io_pp_37[31]; // @[wallace.scala 71:19]
  assign FullAdder_562_io_a = io_pp_38[30]; // @[wallace.scala 69:18]
  assign FullAdder_562_io_b = io_pp_39[29]; // @[wallace.scala 70:18]
  assign FullAdder_562_io_ci = io_pp_40[28]; // @[wallace.scala 71:19]
  assign FullAdder_563_io_a = io_pp_41[27]; // @[wallace.scala 69:18]
  assign FullAdder_563_io_b = io_pp_42[26]; // @[wallace.scala 70:18]
  assign FullAdder_563_io_ci = io_pp_43[25]; // @[wallace.scala 71:19]
  assign FullAdder_564_io_a = io_pp_44[24]; // @[wallace.scala 69:18]
  assign FullAdder_564_io_b = io_pp_45[23]; // @[wallace.scala 70:18]
  assign FullAdder_564_io_ci = io_pp_46[22]; // @[wallace.scala 71:19]
  assign FullAdder_565_io_a = io_pp_47[21]; // @[wallace.scala 69:18]
  assign FullAdder_565_io_b = io_pp_48[20]; // @[wallace.scala 70:18]
  assign FullAdder_565_io_ci = io_pp_49[19]; // @[wallace.scala 71:19]
  assign FullAdder_566_io_a = io_pp_50[18]; // @[wallace.scala 69:18]
  assign FullAdder_566_io_b = io_pp_51[17]; // @[wallace.scala 70:18]
  assign FullAdder_566_io_ci = io_pp_52[16]; // @[wallace.scala 71:19]
  assign FullAdder_567_io_a = io_pp_53[15]; // @[wallace.scala 69:18]
  assign FullAdder_567_io_b = io_pp_54[14]; // @[wallace.scala 70:18]
  assign FullAdder_567_io_ci = io_pp_55[13]; // @[wallace.scala 71:19]
  assign FullAdder_568_io_a = io_pp_56[12]; // @[wallace.scala 69:18]
  assign FullAdder_568_io_b = io_pp_57[11]; // @[wallace.scala 70:18]
  assign FullAdder_568_io_ci = io_pp_58[10]; // @[wallace.scala 71:19]
  assign FullAdder_569_io_a = io_pp_59[9]; // @[wallace.scala 69:18]
  assign FullAdder_569_io_b = io_pp_60[8]; // @[wallace.scala 70:18]
  assign FullAdder_569_io_ci = io_pp_61[7]; // @[wallace.scala 71:19]
  assign HalfAdder_16_io_a = io_pp_62[6]; // @[wallace.scala 59:18]
  assign HalfAdder_16_io_b = io_pp_63[5]; // @[wallace.scala 60:18]
  assign FullAdder_570_io_a = io_pp_4[63]; // @[wallace.scala 69:18]
  assign FullAdder_570_io_b = io_pp_5[62]; // @[wallace.scala 70:18]
  assign FullAdder_570_io_ci = io_pp_6[61]; // @[wallace.scala 71:19]
  assign FullAdder_571_io_a = io_pp_7[60]; // @[wallace.scala 69:18]
  assign FullAdder_571_io_b = io_pp_8[59]; // @[wallace.scala 70:18]
  assign FullAdder_571_io_ci = io_pp_9[58]; // @[wallace.scala 71:19]
  assign FullAdder_572_io_a = io_pp_10[57]; // @[wallace.scala 69:18]
  assign FullAdder_572_io_b = io_pp_11[56]; // @[wallace.scala 70:18]
  assign FullAdder_572_io_ci = io_pp_12[55]; // @[wallace.scala 71:19]
  assign FullAdder_573_io_a = io_pp_13[54]; // @[wallace.scala 69:18]
  assign FullAdder_573_io_b = io_pp_14[53]; // @[wallace.scala 70:18]
  assign FullAdder_573_io_ci = io_pp_15[52]; // @[wallace.scala 71:19]
  assign FullAdder_574_io_a = io_pp_16[51]; // @[wallace.scala 69:18]
  assign FullAdder_574_io_b = io_pp_17[50]; // @[wallace.scala 70:18]
  assign FullAdder_574_io_ci = io_pp_18[49]; // @[wallace.scala 71:19]
  assign FullAdder_575_io_a = io_pp_19[48]; // @[wallace.scala 69:18]
  assign FullAdder_575_io_b = io_pp_20[47]; // @[wallace.scala 70:18]
  assign FullAdder_575_io_ci = io_pp_21[46]; // @[wallace.scala 71:19]
  assign FullAdder_576_io_a = io_pp_22[45]; // @[wallace.scala 69:18]
  assign FullAdder_576_io_b = io_pp_23[44]; // @[wallace.scala 70:18]
  assign FullAdder_576_io_ci = io_pp_24[43]; // @[wallace.scala 71:19]
  assign FullAdder_577_io_a = io_pp_25[42]; // @[wallace.scala 69:18]
  assign FullAdder_577_io_b = io_pp_26[41]; // @[wallace.scala 70:18]
  assign FullAdder_577_io_ci = io_pp_27[40]; // @[wallace.scala 71:19]
  assign FullAdder_578_io_a = io_pp_28[39]; // @[wallace.scala 69:18]
  assign FullAdder_578_io_b = io_pp_29[38]; // @[wallace.scala 70:18]
  assign FullAdder_578_io_ci = io_pp_30[37]; // @[wallace.scala 71:19]
  assign FullAdder_579_io_a = io_pp_31[36]; // @[wallace.scala 69:18]
  assign FullAdder_579_io_b = io_pp_32[35]; // @[wallace.scala 70:18]
  assign FullAdder_579_io_ci = io_pp_33[34]; // @[wallace.scala 71:19]
  assign FullAdder_580_io_a = io_pp_34[33]; // @[wallace.scala 69:18]
  assign FullAdder_580_io_b = io_pp_35[32]; // @[wallace.scala 70:18]
  assign FullAdder_580_io_ci = io_pp_36[31]; // @[wallace.scala 71:19]
  assign FullAdder_581_io_a = io_pp_37[30]; // @[wallace.scala 69:18]
  assign FullAdder_581_io_b = io_pp_38[29]; // @[wallace.scala 70:18]
  assign FullAdder_581_io_ci = io_pp_39[28]; // @[wallace.scala 71:19]
  assign FullAdder_582_io_a = io_pp_40[27]; // @[wallace.scala 69:18]
  assign FullAdder_582_io_b = io_pp_41[26]; // @[wallace.scala 70:18]
  assign FullAdder_582_io_ci = io_pp_42[25]; // @[wallace.scala 71:19]
  assign FullAdder_583_io_a = io_pp_43[24]; // @[wallace.scala 69:18]
  assign FullAdder_583_io_b = io_pp_44[23]; // @[wallace.scala 70:18]
  assign FullAdder_583_io_ci = io_pp_45[22]; // @[wallace.scala 71:19]
  assign FullAdder_584_io_a = io_pp_46[21]; // @[wallace.scala 69:18]
  assign FullAdder_584_io_b = io_pp_47[20]; // @[wallace.scala 70:18]
  assign FullAdder_584_io_ci = io_pp_48[19]; // @[wallace.scala 71:19]
  assign FullAdder_585_io_a = io_pp_49[18]; // @[wallace.scala 69:18]
  assign FullAdder_585_io_b = io_pp_50[17]; // @[wallace.scala 70:18]
  assign FullAdder_585_io_ci = io_pp_51[16]; // @[wallace.scala 71:19]
  assign FullAdder_586_io_a = io_pp_52[15]; // @[wallace.scala 69:18]
  assign FullAdder_586_io_b = io_pp_53[14]; // @[wallace.scala 70:18]
  assign FullAdder_586_io_ci = io_pp_54[13]; // @[wallace.scala 71:19]
  assign FullAdder_587_io_a = io_pp_55[12]; // @[wallace.scala 69:18]
  assign FullAdder_587_io_b = io_pp_56[11]; // @[wallace.scala 70:18]
  assign FullAdder_587_io_ci = io_pp_57[10]; // @[wallace.scala 71:19]
  assign FullAdder_588_io_a = io_pp_58[9]; // @[wallace.scala 69:18]
  assign FullAdder_588_io_b = io_pp_59[8]; // @[wallace.scala 70:18]
  assign FullAdder_588_io_ci = io_pp_60[7]; // @[wallace.scala 71:19]
  assign FullAdder_589_io_a = io_pp_61[6]; // @[wallace.scala 69:18]
  assign FullAdder_589_io_b = io_pp_62[5]; // @[wallace.scala 70:18]
  assign FullAdder_589_io_ci = io_pp_63[4]; // @[wallace.scala 71:19]
  assign FullAdder_590_io_a = io_pp_3[63]; // @[wallace.scala 69:18]
  assign FullAdder_590_io_b = io_pp_4[62]; // @[wallace.scala 70:18]
  assign FullAdder_590_io_ci = io_pp_5[61]; // @[wallace.scala 71:19]
  assign FullAdder_591_io_a = io_pp_6[60]; // @[wallace.scala 69:18]
  assign FullAdder_591_io_b = io_pp_7[59]; // @[wallace.scala 70:18]
  assign FullAdder_591_io_ci = io_pp_8[58]; // @[wallace.scala 71:19]
  assign FullAdder_592_io_a = io_pp_9[57]; // @[wallace.scala 69:18]
  assign FullAdder_592_io_b = io_pp_10[56]; // @[wallace.scala 70:18]
  assign FullAdder_592_io_ci = io_pp_11[55]; // @[wallace.scala 71:19]
  assign FullAdder_593_io_a = io_pp_12[54]; // @[wallace.scala 69:18]
  assign FullAdder_593_io_b = io_pp_13[53]; // @[wallace.scala 70:18]
  assign FullAdder_593_io_ci = io_pp_14[52]; // @[wallace.scala 71:19]
  assign FullAdder_594_io_a = io_pp_15[51]; // @[wallace.scala 69:18]
  assign FullAdder_594_io_b = io_pp_16[50]; // @[wallace.scala 70:18]
  assign FullAdder_594_io_ci = io_pp_17[49]; // @[wallace.scala 71:19]
  assign FullAdder_595_io_a = io_pp_18[48]; // @[wallace.scala 69:18]
  assign FullAdder_595_io_b = io_pp_19[47]; // @[wallace.scala 70:18]
  assign FullAdder_595_io_ci = io_pp_20[46]; // @[wallace.scala 71:19]
  assign FullAdder_596_io_a = io_pp_21[45]; // @[wallace.scala 69:18]
  assign FullAdder_596_io_b = io_pp_22[44]; // @[wallace.scala 70:18]
  assign FullAdder_596_io_ci = io_pp_23[43]; // @[wallace.scala 71:19]
  assign FullAdder_597_io_a = io_pp_24[42]; // @[wallace.scala 69:18]
  assign FullAdder_597_io_b = io_pp_25[41]; // @[wallace.scala 70:18]
  assign FullAdder_597_io_ci = io_pp_26[40]; // @[wallace.scala 71:19]
  assign FullAdder_598_io_a = io_pp_27[39]; // @[wallace.scala 69:18]
  assign FullAdder_598_io_b = io_pp_28[38]; // @[wallace.scala 70:18]
  assign FullAdder_598_io_ci = io_pp_29[37]; // @[wallace.scala 71:19]
  assign FullAdder_599_io_a = io_pp_30[36]; // @[wallace.scala 69:18]
  assign FullAdder_599_io_b = io_pp_31[35]; // @[wallace.scala 70:18]
  assign FullAdder_599_io_ci = io_pp_32[34]; // @[wallace.scala 71:19]
  assign FullAdder_600_io_a = io_pp_33[33]; // @[wallace.scala 69:18]
  assign FullAdder_600_io_b = io_pp_34[32]; // @[wallace.scala 70:18]
  assign FullAdder_600_io_ci = io_pp_35[31]; // @[wallace.scala 71:19]
  assign FullAdder_601_io_a = io_pp_36[30]; // @[wallace.scala 69:18]
  assign FullAdder_601_io_b = io_pp_37[29]; // @[wallace.scala 70:18]
  assign FullAdder_601_io_ci = io_pp_38[28]; // @[wallace.scala 71:19]
  assign FullAdder_602_io_a = io_pp_39[27]; // @[wallace.scala 69:18]
  assign FullAdder_602_io_b = io_pp_40[26]; // @[wallace.scala 70:18]
  assign FullAdder_602_io_ci = io_pp_41[25]; // @[wallace.scala 71:19]
  assign FullAdder_603_io_a = io_pp_42[24]; // @[wallace.scala 69:18]
  assign FullAdder_603_io_b = io_pp_43[23]; // @[wallace.scala 70:18]
  assign FullAdder_603_io_ci = io_pp_44[22]; // @[wallace.scala 71:19]
  assign FullAdder_604_io_a = io_pp_45[21]; // @[wallace.scala 69:18]
  assign FullAdder_604_io_b = io_pp_46[20]; // @[wallace.scala 70:18]
  assign FullAdder_604_io_ci = io_pp_47[19]; // @[wallace.scala 71:19]
  assign FullAdder_605_io_a = io_pp_48[18]; // @[wallace.scala 69:18]
  assign FullAdder_605_io_b = io_pp_49[17]; // @[wallace.scala 70:18]
  assign FullAdder_605_io_ci = io_pp_50[16]; // @[wallace.scala 71:19]
  assign FullAdder_606_io_a = io_pp_51[15]; // @[wallace.scala 69:18]
  assign FullAdder_606_io_b = io_pp_52[14]; // @[wallace.scala 70:18]
  assign FullAdder_606_io_ci = io_pp_53[13]; // @[wallace.scala 71:19]
  assign FullAdder_607_io_a = io_pp_54[12]; // @[wallace.scala 69:18]
  assign FullAdder_607_io_b = io_pp_55[11]; // @[wallace.scala 70:18]
  assign FullAdder_607_io_ci = io_pp_56[10]; // @[wallace.scala 71:19]
  assign FullAdder_608_io_a = io_pp_57[9]; // @[wallace.scala 69:18]
  assign FullAdder_608_io_b = io_pp_58[8]; // @[wallace.scala 70:18]
  assign FullAdder_608_io_ci = io_pp_59[7]; // @[wallace.scala 71:19]
  assign FullAdder_609_io_a = io_pp_60[6]; // @[wallace.scala 69:18]
  assign FullAdder_609_io_b = io_pp_61[5]; // @[wallace.scala 70:18]
  assign FullAdder_609_io_ci = io_pp_62[4]; // @[wallace.scala 71:19]
  assign FullAdder_610_io_a = io_pp_2[63]; // @[wallace.scala 69:18]
  assign FullAdder_610_io_b = io_pp_3[62]; // @[wallace.scala 70:18]
  assign FullAdder_610_io_ci = io_pp_4[61]; // @[wallace.scala 71:19]
  assign FullAdder_611_io_a = io_pp_5[60]; // @[wallace.scala 69:18]
  assign FullAdder_611_io_b = io_pp_6[59]; // @[wallace.scala 70:18]
  assign FullAdder_611_io_ci = io_pp_7[58]; // @[wallace.scala 71:19]
  assign FullAdder_612_io_a = io_pp_8[57]; // @[wallace.scala 69:18]
  assign FullAdder_612_io_b = io_pp_9[56]; // @[wallace.scala 70:18]
  assign FullAdder_612_io_ci = io_pp_10[55]; // @[wallace.scala 71:19]
  assign FullAdder_613_io_a = io_pp_11[54]; // @[wallace.scala 69:18]
  assign FullAdder_613_io_b = io_pp_12[53]; // @[wallace.scala 70:18]
  assign FullAdder_613_io_ci = io_pp_13[52]; // @[wallace.scala 71:19]
  assign FullAdder_614_io_a = io_pp_14[51]; // @[wallace.scala 69:18]
  assign FullAdder_614_io_b = io_pp_15[50]; // @[wallace.scala 70:18]
  assign FullAdder_614_io_ci = io_pp_16[49]; // @[wallace.scala 71:19]
  assign FullAdder_615_io_a = io_pp_17[48]; // @[wallace.scala 69:18]
  assign FullAdder_615_io_b = io_pp_18[47]; // @[wallace.scala 70:18]
  assign FullAdder_615_io_ci = io_pp_19[46]; // @[wallace.scala 71:19]
  assign FullAdder_616_io_a = io_pp_20[45]; // @[wallace.scala 69:18]
  assign FullAdder_616_io_b = io_pp_21[44]; // @[wallace.scala 70:18]
  assign FullAdder_616_io_ci = io_pp_22[43]; // @[wallace.scala 71:19]
  assign FullAdder_617_io_a = io_pp_23[42]; // @[wallace.scala 69:18]
  assign FullAdder_617_io_b = io_pp_24[41]; // @[wallace.scala 70:18]
  assign FullAdder_617_io_ci = io_pp_25[40]; // @[wallace.scala 71:19]
  assign FullAdder_618_io_a = io_pp_26[39]; // @[wallace.scala 69:18]
  assign FullAdder_618_io_b = io_pp_27[38]; // @[wallace.scala 70:18]
  assign FullAdder_618_io_ci = io_pp_28[37]; // @[wallace.scala 71:19]
  assign FullAdder_619_io_a = io_pp_29[36]; // @[wallace.scala 69:18]
  assign FullAdder_619_io_b = io_pp_30[35]; // @[wallace.scala 70:18]
  assign FullAdder_619_io_ci = io_pp_31[34]; // @[wallace.scala 71:19]
  assign FullAdder_620_io_a = io_pp_32[33]; // @[wallace.scala 69:18]
  assign FullAdder_620_io_b = io_pp_33[32]; // @[wallace.scala 70:18]
  assign FullAdder_620_io_ci = io_pp_34[31]; // @[wallace.scala 71:19]
  assign FullAdder_621_io_a = io_pp_35[30]; // @[wallace.scala 69:18]
  assign FullAdder_621_io_b = io_pp_36[29]; // @[wallace.scala 70:18]
  assign FullAdder_621_io_ci = io_pp_37[28]; // @[wallace.scala 71:19]
  assign FullAdder_622_io_a = io_pp_38[27]; // @[wallace.scala 69:18]
  assign FullAdder_622_io_b = io_pp_39[26]; // @[wallace.scala 70:18]
  assign FullAdder_622_io_ci = io_pp_40[25]; // @[wallace.scala 71:19]
  assign FullAdder_623_io_a = io_pp_41[24]; // @[wallace.scala 69:18]
  assign FullAdder_623_io_b = io_pp_42[23]; // @[wallace.scala 70:18]
  assign FullAdder_623_io_ci = io_pp_43[22]; // @[wallace.scala 71:19]
  assign FullAdder_624_io_a = io_pp_44[21]; // @[wallace.scala 69:18]
  assign FullAdder_624_io_b = io_pp_45[20]; // @[wallace.scala 70:18]
  assign FullAdder_624_io_ci = io_pp_46[19]; // @[wallace.scala 71:19]
  assign FullAdder_625_io_a = io_pp_47[18]; // @[wallace.scala 69:18]
  assign FullAdder_625_io_b = io_pp_48[17]; // @[wallace.scala 70:18]
  assign FullAdder_625_io_ci = io_pp_49[16]; // @[wallace.scala 71:19]
  assign FullAdder_626_io_a = io_pp_50[15]; // @[wallace.scala 69:18]
  assign FullAdder_626_io_b = io_pp_51[14]; // @[wallace.scala 70:18]
  assign FullAdder_626_io_ci = io_pp_52[13]; // @[wallace.scala 71:19]
  assign FullAdder_627_io_a = io_pp_53[12]; // @[wallace.scala 69:18]
  assign FullAdder_627_io_b = io_pp_54[11]; // @[wallace.scala 70:18]
  assign FullAdder_627_io_ci = io_pp_55[10]; // @[wallace.scala 71:19]
  assign FullAdder_628_io_a = io_pp_56[9]; // @[wallace.scala 69:18]
  assign FullAdder_628_io_b = io_pp_57[8]; // @[wallace.scala 70:18]
  assign FullAdder_628_io_ci = io_pp_58[7]; // @[wallace.scala 71:19]
  assign FullAdder_629_io_a = io_pp_59[6]; // @[wallace.scala 69:18]
  assign FullAdder_629_io_b = io_pp_60[5]; // @[wallace.scala 70:18]
  assign FullAdder_629_io_ci = io_pp_61[4]; // @[wallace.scala 71:19]
  assign HalfAdder_17_io_a = io_pp_62[3]; // @[wallace.scala 59:18]
  assign HalfAdder_17_io_b = io_pp_63[2]; // @[wallace.scala 60:18]
  assign FullAdder_630_io_a = io_pp_1[63]; // @[wallace.scala 69:18]
  assign FullAdder_630_io_b = io_pp_2[62]; // @[wallace.scala 70:18]
  assign FullAdder_630_io_ci = io_pp_3[61]; // @[wallace.scala 71:19]
  assign FullAdder_631_io_a = io_pp_4[60]; // @[wallace.scala 69:18]
  assign FullAdder_631_io_b = io_pp_5[59]; // @[wallace.scala 70:18]
  assign FullAdder_631_io_ci = io_pp_6[58]; // @[wallace.scala 71:19]
  assign FullAdder_632_io_a = io_pp_7[57]; // @[wallace.scala 69:18]
  assign FullAdder_632_io_b = io_pp_8[56]; // @[wallace.scala 70:18]
  assign FullAdder_632_io_ci = io_pp_9[55]; // @[wallace.scala 71:19]
  assign FullAdder_633_io_a = io_pp_10[54]; // @[wallace.scala 69:18]
  assign FullAdder_633_io_b = io_pp_11[53]; // @[wallace.scala 70:18]
  assign FullAdder_633_io_ci = io_pp_12[52]; // @[wallace.scala 71:19]
  assign FullAdder_634_io_a = io_pp_13[51]; // @[wallace.scala 69:18]
  assign FullAdder_634_io_b = io_pp_14[50]; // @[wallace.scala 70:18]
  assign FullAdder_634_io_ci = io_pp_15[49]; // @[wallace.scala 71:19]
  assign FullAdder_635_io_a = io_pp_16[48]; // @[wallace.scala 69:18]
  assign FullAdder_635_io_b = io_pp_17[47]; // @[wallace.scala 70:18]
  assign FullAdder_635_io_ci = io_pp_18[46]; // @[wallace.scala 71:19]
  assign FullAdder_636_io_a = io_pp_19[45]; // @[wallace.scala 69:18]
  assign FullAdder_636_io_b = io_pp_20[44]; // @[wallace.scala 70:18]
  assign FullAdder_636_io_ci = io_pp_21[43]; // @[wallace.scala 71:19]
  assign FullAdder_637_io_a = io_pp_22[42]; // @[wallace.scala 69:18]
  assign FullAdder_637_io_b = io_pp_23[41]; // @[wallace.scala 70:18]
  assign FullAdder_637_io_ci = io_pp_24[40]; // @[wallace.scala 71:19]
  assign FullAdder_638_io_a = io_pp_25[39]; // @[wallace.scala 69:18]
  assign FullAdder_638_io_b = io_pp_26[38]; // @[wallace.scala 70:18]
  assign FullAdder_638_io_ci = io_pp_27[37]; // @[wallace.scala 71:19]
  assign FullAdder_639_io_a = io_pp_28[36]; // @[wallace.scala 69:18]
  assign FullAdder_639_io_b = io_pp_29[35]; // @[wallace.scala 70:18]
  assign FullAdder_639_io_ci = io_pp_30[34]; // @[wallace.scala 71:19]
  assign FullAdder_640_io_a = io_pp_31[33]; // @[wallace.scala 69:18]
  assign FullAdder_640_io_b = io_pp_32[32]; // @[wallace.scala 70:18]
  assign FullAdder_640_io_ci = io_pp_33[31]; // @[wallace.scala 71:19]
  assign FullAdder_641_io_a = io_pp_34[30]; // @[wallace.scala 69:18]
  assign FullAdder_641_io_b = io_pp_35[29]; // @[wallace.scala 70:18]
  assign FullAdder_641_io_ci = io_pp_36[28]; // @[wallace.scala 71:19]
  assign FullAdder_642_io_a = io_pp_37[27]; // @[wallace.scala 69:18]
  assign FullAdder_642_io_b = io_pp_38[26]; // @[wallace.scala 70:18]
  assign FullAdder_642_io_ci = io_pp_39[25]; // @[wallace.scala 71:19]
  assign FullAdder_643_io_a = io_pp_40[24]; // @[wallace.scala 69:18]
  assign FullAdder_643_io_b = io_pp_41[23]; // @[wallace.scala 70:18]
  assign FullAdder_643_io_ci = io_pp_42[22]; // @[wallace.scala 71:19]
  assign FullAdder_644_io_a = io_pp_43[21]; // @[wallace.scala 69:18]
  assign FullAdder_644_io_b = io_pp_44[20]; // @[wallace.scala 70:18]
  assign FullAdder_644_io_ci = io_pp_45[19]; // @[wallace.scala 71:19]
  assign FullAdder_645_io_a = io_pp_46[18]; // @[wallace.scala 69:18]
  assign FullAdder_645_io_b = io_pp_47[17]; // @[wallace.scala 70:18]
  assign FullAdder_645_io_ci = io_pp_48[16]; // @[wallace.scala 71:19]
  assign FullAdder_646_io_a = io_pp_49[15]; // @[wallace.scala 69:18]
  assign FullAdder_646_io_b = io_pp_50[14]; // @[wallace.scala 70:18]
  assign FullAdder_646_io_ci = io_pp_51[13]; // @[wallace.scala 71:19]
  assign FullAdder_647_io_a = io_pp_52[12]; // @[wallace.scala 69:18]
  assign FullAdder_647_io_b = io_pp_53[11]; // @[wallace.scala 70:18]
  assign FullAdder_647_io_ci = io_pp_54[10]; // @[wallace.scala 71:19]
  assign FullAdder_648_io_a = io_pp_55[9]; // @[wallace.scala 69:18]
  assign FullAdder_648_io_b = io_pp_56[8]; // @[wallace.scala 70:18]
  assign FullAdder_648_io_ci = io_pp_57[7]; // @[wallace.scala 71:19]
  assign FullAdder_649_io_a = io_pp_58[6]; // @[wallace.scala 69:18]
  assign FullAdder_649_io_b = io_pp_59[5]; // @[wallace.scala 70:18]
  assign FullAdder_649_io_ci = io_pp_60[4]; // @[wallace.scala 71:19]
  assign FullAdder_650_io_a = io_pp_61[3]; // @[wallace.scala 69:18]
  assign FullAdder_650_io_b = io_pp_62[2]; // @[wallace.scala 70:18]
  assign FullAdder_650_io_ci = io_pp_63[1]; // @[wallace.scala 71:19]
  assign FullAdder_651_io_a = io_pp_0[63]; // @[wallace.scala 69:18]
  assign FullAdder_651_io_b = io_pp_1[62]; // @[wallace.scala 70:18]
  assign FullAdder_651_io_ci = io_pp_2[61]; // @[wallace.scala 71:19]
  assign FullAdder_652_io_a = io_pp_3[60]; // @[wallace.scala 69:18]
  assign FullAdder_652_io_b = io_pp_4[59]; // @[wallace.scala 70:18]
  assign FullAdder_652_io_ci = io_pp_5[58]; // @[wallace.scala 71:19]
  assign FullAdder_653_io_a = io_pp_6[57]; // @[wallace.scala 69:18]
  assign FullAdder_653_io_b = io_pp_7[56]; // @[wallace.scala 70:18]
  assign FullAdder_653_io_ci = io_pp_8[55]; // @[wallace.scala 71:19]
  assign FullAdder_654_io_a = io_pp_9[54]; // @[wallace.scala 69:18]
  assign FullAdder_654_io_b = io_pp_10[53]; // @[wallace.scala 70:18]
  assign FullAdder_654_io_ci = io_pp_11[52]; // @[wallace.scala 71:19]
  assign FullAdder_655_io_a = io_pp_12[51]; // @[wallace.scala 69:18]
  assign FullAdder_655_io_b = io_pp_13[50]; // @[wallace.scala 70:18]
  assign FullAdder_655_io_ci = io_pp_14[49]; // @[wallace.scala 71:19]
  assign FullAdder_656_io_a = io_pp_15[48]; // @[wallace.scala 69:18]
  assign FullAdder_656_io_b = io_pp_16[47]; // @[wallace.scala 70:18]
  assign FullAdder_656_io_ci = io_pp_17[46]; // @[wallace.scala 71:19]
  assign FullAdder_657_io_a = io_pp_18[45]; // @[wallace.scala 69:18]
  assign FullAdder_657_io_b = io_pp_19[44]; // @[wallace.scala 70:18]
  assign FullAdder_657_io_ci = io_pp_20[43]; // @[wallace.scala 71:19]
  assign FullAdder_658_io_a = io_pp_21[42]; // @[wallace.scala 69:18]
  assign FullAdder_658_io_b = io_pp_22[41]; // @[wallace.scala 70:18]
  assign FullAdder_658_io_ci = io_pp_23[40]; // @[wallace.scala 71:19]
  assign FullAdder_659_io_a = io_pp_24[39]; // @[wallace.scala 69:18]
  assign FullAdder_659_io_b = io_pp_25[38]; // @[wallace.scala 70:18]
  assign FullAdder_659_io_ci = io_pp_26[37]; // @[wallace.scala 71:19]
  assign FullAdder_660_io_a = io_pp_27[36]; // @[wallace.scala 69:18]
  assign FullAdder_660_io_b = io_pp_28[35]; // @[wallace.scala 70:18]
  assign FullAdder_660_io_ci = io_pp_29[34]; // @[wallace.scala 71:19]
  assign FullAdder_661_io_a = io_pp_30[33]; // @[wallace.scala 69:18]
  assign FullAdder_661_io_b = io_pp_31[32]; // @[wallace.scala 70:18]
  assign FullAdder_661_io_ci = io_pp_32[31]; // @[wallace.scala 71:19]
  assign FullAdder_662_io_a = io_pp_33[30]; // @[wallace.scala 69:18]
  assign FullAdder_662_io_b = io_pp_34[29]; // @[wallace.scala 70:18]
  assign FullAdder_662_io_ci = io_pp_35[28]; // @[wallace.scala 71:19]
  assign FullAdder_663_io_a = io_pp_36[27]; // @[wallace.scala 69:18]
  assign FullAdder_663_io_b = io_pp_37[26]; // @[wallace.scala 70:18]
  assign FullAdder_663_io_ci = io_pp_38[25]; // @[wallace.scala 71:19]
  assign FullAdder_664_io_a = io_pp_39[24]; // @[wallace.scala 69:18]
  assign FullAdder_664_io_b = io_pp_40[23]; // @[wallace.scala 70:18]
  assign FullAdder_664_io_ci = io_pp_41[22]; // @[wallace.scala 71:19]
  assign FullAdder_665_io_a = io_pp_42[21]; // @[wallace.scala 69:18]
  assign FullAdder_665_io_b = io_pp_43[20]; // @[wallace.scala 70:18]
  assign FullAdder_665_io_ci = io_pp_44[19]; // @[wallace.scala 71:19]
  assign FullAdder_666_io_a = io_pp_45[18]; // @[wallace.scala 69:18]
  assign FullAdder_666_io_b = io_pp_46[17]; // @[wallace.scala 70:18]
  assign FullAdder_666_io_ci = io_pp_47[16]; // @[wallace.scala 71:19]
  assign FullAdder_667_io_a = io_pp_48[15]; // @[wallace.scala 69:18]
  assign FullAdder_667_io_b = io_pp_49[14]; // @[wallace.scala 70:18]
  assign FullAdder_667_io_ci = io_pp_50[13]; // @[wallace.scala 71:19]
  assign FullAdder_668_io_a = io_pp_51[12]; // @[wallace.scala 69:18]
  assign FullAdder_668_io_b = io_pp_52[11]; // @[wallace.scala 70:18]
  assign FullAdder_668_io_ci = io_pp_53[10]; // @[wallace.scala 71:19]
  assign FullAdder_669_io_a = io_pp_54[9]; // @[wallace.scala 69:18]
  assign FullAdder_669_io_b = io_pp_55[8]; // @[wallace.scala 70:18]
  assign FullAdder_669_io_ci = io_pp_56[7]; // @[wallace.scala 71:19]
  assign FullAdder_670_io_a = io_pp_57[6]; // @[wallace.scala 69:18]
  assign FullAdder_670_io_b = io_pp_58[5]; // @[wallace.scala 70:18]
  assign FullAdder_670_io_ci = io_pp_59[4]; // @[wallace.scala 71:19]
  assign FullAdder_671_io_a = io_pp_60[3]; // @[wallace.scala 69:18]
  assign FullAdder_671_io_b = io_pp_61[2]; // @[wallace.scala 70:18]
  assign FullAdder_671_io_ci = io_pp_62[1]; // @[wallace.scala 71:19]
  assign FullAdder_672_io_a = io_pp_0[62]; // @[wallace.scala 69:18]
  assign FullAdder_672_io_b = io_pp_1[61]; // @[wallace.scala 70:18]
  assign FullAdder_672_io_ci = io_pp_2[60]; // @[wallace.scala 71:19]
  assign FullAdder_673_io_a = io_pp_3[59]; // @[wallace.scala 69:18]
  assign FullAdder_673_io_b = io_pp_4[58]; // @[wallace.scala 70:18]
  assign FullAdder_673_io_ci = io_pp_5[57]; // @[wallace.scala 71:19]
  assign FullAdder_674_io_a = io_pp_6[56]; // @[wallace.scala 69:18]
  assign FullAdder_674_io_b = io_pp_7[55]; // @[wallace.scala 70:18]
  assign FullAdder_674_io_ci = io_pp_8[54]; // @[wallace.scala 71:19]
  assign FullAdder_675_io_a = io_pp_9[53]; // @[wallace.scala 69:18]
  assign FullAdder_675_io_b = io_pp_10[52]; // @[wallace.scala 70:18]
  assign FullAdder_675_io_ci = io_pp_11[51]; // @[wallace.scala 71:19]
  assign FullAdder_676_io_a = io_pp_12[50]; // @[wallace.scala 69:18]
  assign FullAdder_676_io_b = io_pp_13[49]; // @[wallace.scala 70:18]
  assign FullAdder_676_io_ci = io_pp_14[48]; // @[wallace.scala 71:19]
  assign FullAdder_677_io_a = io_pp_15[47]; // @[wallace.scala 69:18]
  assign FullAdder_677_io_b = io_pp_16[46]; // @[wallace.scala 70:18]
  assign FullAdder_677_io_ci = io_pp_17[45]; // @[wallace.scala 71:19]
  assign FullAdder_678_io_a = io_pp_18[44]; // @[wallace.scala 69:18]
  assign FullAdder_678_io_b = io_pp_19[43]; // @[wallace.scala 70:18]
  assign FullAdder_678_io_ci = io_pp_20[42]; // @[wallace.scala 71:19]
  assign FullAdder_679_io_a = io_pp_21[41]; // @[wallace.scala 69:18]
  assign FullAdder_679_io_b = io_pp_22[40]; // @[wallace.scala 70:18]
  assign FullAdder_679_io_ci = io_pp_23[39]; // @[wallace.scala 71:19]
  assign FullAdder_680_io_a = io_pp_24[38]; // @[wallace.scala 69:18]
  assign FullAdder_680_io_b = io_pp_25[37]; // @[wallace.scala 70:18]
  assign FullAdder_680_io_ci = io_pp_26[36]; // @[wallace.scala 71:19]
  assign FullAdder_681_io_a = io_pp_27[35]; // @[wallace.scala 69:18]
  assign FullAdder_681_io_b = io_pp_28[34]; // @[wallace.scala 70:18]
  assign FullAdder_681_io_ci = io_pp_29[33]; // @[wallace.scala 71:19]
  assign FullAdder_682_io_a = io_pp_30[32]; // @[wallace.scala 69:18]
  assign FullAdder_682_io_b = io_pp_31[31]; // @[wallace.scala 70:18]
  assign FullAdder_682_io_ci = io_pp_32[30]; // @[wallace.scala 71:19]
  assign FullAdder_683_io_a = io_pp_33[29]; // @[wallace.scala 69:18]
  assign FullAdder_683_io_b = io_pp_34[28]; // @[wallace.scala 70:18]
  assign FullAdder_683_io_ci = io_pp_35[27]; // @[wallace.scala 71:19]
  assign FullAdder_684_io_a = io_pp_36[26]; // @[wallace.scala 69:18]
  assign FullAdder_684_io_b = io_pp_37[25]; // @[wallace.scala 70:18]
  assign FullAdder_684_io_ci = io_pp_38[24]; // @[wallace.scala 71:19]
  assign FullAdder_685_io_a = io_pp_39[23]; // @[wallace.scala 69:18]
  assign FullAdder_685_io_b = io_pp_40[22]; // @[wallace.scala 70:18]
  assign FullAdder_685_io_ci = io_pp_41[21]; // @[wallace.scala 71:19]
  assign FullAdder_686_io_a = io_pp_42[20]; // @[wallace.scala 69:18]
  assign FullAdder_686_io_b = io_pp_43[19]; // @[wallace.scala 70:18]
  assign FullAdder_686_io_ci = io_pp_44[18]; // @[wallace.scala 71:19]
  assign FullAdder_687_io_a = io_pp_45[17]; // @[wallace.scala 69:18]
  assign FullAdder_687_io_b = io_pp_46[16]; // @[wallace.scala 70:18]
  assign FullAdder_687_io_ci = io_pp_47[15]; // @[wallace.scala 71:19]
  assign FullAdder_688_io_a = io_pp_48[14]; // @[wallace.scala 69:18]
  assign FullAdder_688_io_b = io_pp_49[13]; // @[wallace.scala 70:18]
  assign FullAdder_688_io_ci = io_pp_50[12]; // @[wallace.scala 71:19]
  assign FullAdder_689_io_a = io_pp_51[11]; // @[wallace.scala 69:18]
  assign FullAdder_689_io_b = io_pp_52[10]; // @[wallace.scala 70:18]
  assign FullAdder_689_io_ci = io_pp_53[9]; // @[wallace.scala 71:19]
  assign FullAdder_690_io_a = io_pp_54[8]; // @[wallace.scala 69:18]
  assign FullAdder_690_io_b = io_pp_55[7]; // @[wallace.scala 70:18]
  assign FullAdder_690_io_ci = io_pp_56[6]; // @[wallace.scala 71:19]
  assign FullAdder_691_io_a = io_pp_57[5]; // @[wallace.scala 69:18]
  assign FullAdder_691_io_b = io_pp_58[4]; // @[wallace.scala 70:18]
  assign FullAdder_691_io_ci = io_pp_59[3]; // @[wallace.scala 71:19]
  assign FullAdder_692_io_a = io_pp_60[2]; // @[wallace.scala 69:18]
  assign FullAdder_692_io_b = io_pp_61[1]; // @[wallace.scala 70:18]
  assign FullAdder_692_io_ci = io_pp_62[0]; // @[wallace.scala 71:19]
  assign FullAdder_693_io_a = io_pp_0[61]; // @[wallace.scala 69:18]
  assign FullAdder_693_io_b = io_pp_1[60]; // @[wallace.scala 70:18]
  assign FullAdder_693_io_ci = io_pp_2[59]; // @[wallace.scala 71:19]
  assign FullAdder_694_io_a = io_pp_3[58]; // @[wallace.scala 69:18]
  assign FullAdder_694_io_b = io_pp_4[57]; // @[wallace.scala 70:18]
  assign FullAdder_694_io_ci = io_pp_5[56]; // @[wallace.scala 71:19]
  assign FullAdder_695_io_a = io_pp_6[55]; // @[wallace.scala 69:18]
  assign FullAdder_695_io_b = io_pp_7[54]; // @[wallace.scala 70:18]
  assign FullAdder_695_io_ci = io_pp_8[53]; // @[wallace.scala 71:19]
  assign FullAdder_696_io_a = io_pp_9[52]; // @[wallace.scala 69:18]
  assign FullAdder_696_io_b = io_pp_10[51]; // @[wallace.scala 70:18]
  assign FullAdder_696_io_ci = io_pp_11[50]; // @[wallace.scala 71:19]
  assign FullAdder_697_io_a = io_pp_12[49]; // @[wallace.scala 69:18]
  assign FullAdder_697_io_b = io_pp_13[48]; // @[wallace.scala 70:18]
  assign FullAdder_697_io_ci = io_pp_14[47]; // @[wallace.scala 71:19]
  assign FullAdder_698_io_a = io_pp_15[46]; // @[wallace.scala 69:18]
  assign FullAdder_698_io_b = io_pp_16[45]; // @[wallace.scala 70:18]
  assign FullAdder_698_io_ci = io_pp_17[44]; // @[wallace.scala 71:19]
  assign FullAdder_699_io_a = io_pp_18[43]; // @[wallace.scala 69:18]
  assign FullAdder_699_io_b = io_pp_19[42]; // @[wallace.scala 70:18]
  assign FullAdder_699_io_ci = io_pp_20[41]; // @[wallace.scala 71:19]
  assign FullAdder_700_io_a = io_pp_21[40]; // @[wallace.scala 69:18]
  assign FullAdder_700_io_b = io_pp_22[39]; // @[wallace.scala 70:18]
  assign FullAdder_700_io_ci = io_pp_23[38]; // @[wallace.scala 71:19]
  assign FullAdder_701_io_a = io_pp_24[37]; // @[wallace.scala 69:18]
  assign FullAdder_701_io_b = io_pp_25[36]; // @[wallace.scala 70:18]
  assign FullAdder_701_io_ci = io_pp_26[35]; // @[wallace.scala 71:19]
  assign FullAdder_702_io_a = io_pp_27[34]; // @[wallace.scala 69:18]
  assign FullAdder_702_io_b = io_pp_28[33]; // @[wallace.scala 70:18]
  assign FullAdder_702_io_ci = io_pp_29[32]; // @[wallace.scala 71:19]
  assign FullAdder_703_io_a = io_pp_30[31]; // @[wallace.scala 69:18]
  assign FullAdder_703_io_b = io_pp_31[30]; // @[wallace.scala 70:18]
  assign FullAdder_703_io_ci = io_pp_32[29]; // @[wallace.scala 71:19]
  assign FullAdder_704_io_a = io_pp_33[28]; // @[wallace.scala 69:18]
  assign FullAdder_704_io_b = io_pp_34[27]; // @[wallace.scala 70:18]
  assign FullAdder_704_io_ci = io_pp_35[26]; // @[wallace.scala 71:19]
  assign FullAdder_705_io_a = io_pp_36[25]; // @[wallace.scala 69:18]
  assign FullAdder_705_io_b = io_pp_37[24]; // @[wallace.scala 70:18]
  assign FullAdder_705_io_ci = io_pp_38[23]; // @[wallace.scala 71:19]
  assign FullAdder_706_io_a = io_pp_39[22]; // @[wallace.scala 69:18]
  assign FullAdder_706_io_b = io_pp_40[21]; // @[wallace.scala 70:18]
  assign FullAdder_706_io_ci = io_pp_41[20]; // @[wallace.scala 71:19]
  assign FullAdder_707_io_a = io_pp_42[19]; // @[wallace.scala 69:18]
  assign FullAdder_707_io_b = io_pp_43[18]; // @[wallace.scala 70:18]
  assign FullAdder_707_io_ci = io_pp_44[17]; // @[wallace.scala 71:19]
  assign FullAdder_708_io_a = io_pp_45[16]; // @[wallace.scala 69:18]
  assign FullAdder_708_io_b = io_pp_46[15]; // @[wallace.scala 70:18]
  assign FullAdder_708_io_ci = io_pp_47[14]; // @[wallace.scala 71:19]
  assign FullAdder_709_io_a = io_pp_48[13]; // @[wallace.scala 69:18]
  assign FullAdder_709_io_b = io_pp_49[12]; // @[wallace.scala 70:18]
  assign FullAdder_709_io_ci = io_pp_50[11]; // @[wallace.scala 71:19]
  assign FullAdder_710_io_a = io_pp_51[10]; // @[wallace.scala 69:18]
  assign FullAdder_710_io_b = io_pp_52[9]; // @[wallace.scala 70:18]
  assign FullAdder_710_io_ci = io_pp_53[8]; // @[wallace.scala 71:19]
  assign FullAdder_711_io_a = io_pp_54[7]; // @[wallace.scala 69:18]
  assign FullAdder_711_io_b = io_pp_55[6]; // @[wallace.scala 70:18]
  assign FullAdder_711_io_ci = io_pp_56[5]; // @[wallace.scala 71:19]
  assign FullAdder_712_io_a = io_pp_57[4]; // @[wallace.scala 69:18]
  assign FullAdder_712_io_b = io_pp_58[3]; // @[wallace.scala 70:18]
  assign FullAdder_712_io_ci = io_pp_59[2]; // @[wallace.scala 71:19]
  assign HalfAdder_18_io_a = io_pp_60[1]; // @[wallace.scala 59:18]
  assign HalfAdder_18_io_b = io_pp_61[0]; // @[wallace.scala 60:18]
  assign FullAdder_713_io_a = io_pp_0[60]; // @[wallace.scala 69:18]
  assign FullAdder_713_io_b = io_pp_1[59]; // @[wallace.scala 70:18]
  assign FullAdder_713_io_ci = io_pp_2[58]; // @[wallace.scala 71:19]
  assign FullAdder_714_io_a = io_pp_3[57]; // @[wallace.scala 69:18]
  assign FullAdder_714_io_b = io_pp_4[56]; // @[wallace.scala 70:18]
  assign FullAdder_714_io_ci = io_pp_5[55]; // @[wallace.scala 71:19]
  assign FullAdder_715_io_a = io_pp_6[54]; // @[wallace.scala 69:18]
  assign FullAdder_715_io_b = io_pp_7[53]; // @[wallace.scala 70:18]
  assign FullAdder_715_io_ci = io_pp_8[52]; // @[wallace.scala 71:19]
  assign FullAdder_716_io_a = io_pp_9[51]; // @[wallace.scala 69:18]
  assign FullAdder_716_io_b = io_pp_10[50]; // @[wallace.scala 70:18]
  assign FullAdder_716_io_ci = io_pp_11[49]; // @[wallace.scala 71:19]
  assign FullAdder_717_io_a = io_pp_12[48]; // @[wallace.scala 69:18]
  assign FullAdder_717_io_b = io_pp_13[47]; // @[wallace.scala 70:18]
  assign FullAdder_717_io_ci = io_pp_14[46]; // @[wallace.scala 71:19]
  assign FullAdder_718_io_a = io_pp_15[45]; // @[wallace.scala 69:18]
  assign FullAdder_718_io_b = io_pp_16[44]; // @[wallace.scala 70:18]
  assign FullAdder_718_io_ci = io_pp_17[43]; // @[wallace.scala 71:19]
  assign FullAdder_719_io_a = io_pp_18[42]; // @[wallace.scala 69:18]
  assign FullAdder_719_io_b = io_pp_19[41]; // @[wallace.scala 70:18]
  assign FullAdder_719_io_ci = io_pp_20[40]; // @[wallace.scala 71:19]
  assign FullAdder_720_io_a = io_pp_21[39]; // @[wallace.scala 69:18]
  assign FullAdder_720_io_b = io_pp_22[38]; // @[wallace.scala 70:18]
  assign FullAdder_720_io_ci = io_pp_23[37]; // @[wallace.scala 71:19]
  assign FullAdder_721_io_a = io_pp_24[36]; // @[wallace.scala 69:18]
  assign FullAdder_721_io_b = io_pp_25[35]; // @[wallace.scala 70:18]
  assign FullAdder_721_io_ci = io_pp_26[34]; // @[wallace.scala 71:19]
  assign FullAdder_722_io_a = io_pp_27[33]; // @[wallace.scala 69:18]
  assign FullAdder_722_io_b = io_pp_28[32]; // @[wallace.scala 70:18]
  assign FullAdder_722_io_ci = io_pp_29[31]; // @[wallace.scala 71:19]
  assign FullAdder_723_io_a = io_pp_30[30]; // @[wallace.scala 69:18]
  assign FullAdder_723_io_b = io_pp_31[29]; // @[wallace.scala 70:18]
  assign FullAdder_723_io_ci = io_pp_32[28]; // @[wallace.scala 71:19]
  assign FullAdder_724_io_a = io_pp_33[27]; // @[wallace.scala 69:18]
  assign FullAdder_724_io_b = io_pp_34[26]; // @[wallace.scala 70:18]
  assign FullAdder_724_io_ci = io_pp_35[25]; // @[wallace.scala 71:19]
  assign FullAdder_725_io_a = io_pp_36[24]; // @[wallace.scala 69:18]
  assign FullAdder_725_io_b = io_pp_37[23]; // @[wallace.scala 70:18]
  assign FullAdder_725_io_ci = io_pp_38[22]; // @[wallace.scala 71:19]
  assign FullAdder_726_io_a = io_pp_39[21]; // @[wallace.scala 69:18]
  assign FullAdder_726_io_b = io_pp_40[20]; // @[wallace.scala 70:18]
  assign FullAdder_726_io_ci = io_pp_41[19]; // @[wallace.scala 71:19]
  assign FullAdder_727_io_a = io_pp_42[18]; // @[wallace.scala 69:18]
  assign FullAdder_727_io_b = io_pp_43[17]; // @[wallace.scala 70:18]
  assign FullAdder_727_io_ci = io_pp_44[16]; // @[wallace.scala 71:19]
  assign FullAdder_728_io_a = io_pp_45[15]; // @[wallace.scala 69:18]
  assign FullAdder_728_io_b = io_pp_46[14]; // @[wallace.scala 70:18]
  assign FullAdder_728_io_ci = io_pp_47[13]; // @[wallace.scala 71:19]
  assign FullAdder_729_io_a = io_pp_48[12]; // @[wallace.scala 69:18]
  assign FullAdder_729_io_b = io_pp_49[11]; // @[wallace.scala 70:18]
  assign FullAdder_729_io_ci = io_pp_50[10]; // @[wallace.scala 71:19]
  assign FullAdder_730_io_a = io_pp_51[9]; // @[wallace.scala 69:18]
  assign FullAdder_730_io_b = io_pp_52[8]; // @[wallace.scala 70:18]
  assign FullAdder_730_io_ci = io_pp_53[7]; // @[wallace.scala 71:19]
  assign FullAdder_731_io_a = io_pp_54[6]; // @[wallace.scala 69:18]
  assign FullAdder_731_io_b = io_pp_55[5]; // @[wallace.scala 70:18]
  assign FullAdder_731_io_ci = io_pp_56[4]; // @[wallace.scala 71:19]
  assign FullAdder_732_io_a = io_pp_57[3]; // @[wallace.scala 69:18]
  assign FullAdder_732_io_b = io_pp_58[2]; // @[wallace.scala 70:18]
  assign FullAdder_732_io_ci = io_pp_59[1]; // @[wallace.scala 71:19]
  assign FullAdder_733_io_a = io_pp_0[59]; // @[wallace.scala 69:18]
  assign FullAdder_733_io_b = io_pp_1[58]; // @[wallace.scala 70:18]
  assign FullAdder_733_io_ci = io_pp_2[57]; // @[wallace.scala 71:19]
  assign FullAdder_734_io_a = io_pp_3[56]; // @[wallace.scala 69:18]
  assign FullAdder_734_io_b = io_pp_4[55]; // @[wallace.scala 70:18]
  assign FullAdder_734_io_ci = io_pp_5[54]; // @[wallace.scala 71:19]
  assign FullAdder_735_io_a = io_pp_6[53]; // @[wallace.scala 69:18]
  assign FullAdder_735_io_b = io_pp_7[52]; // @[wallace.scala 70:18]
  assign FullAdder_735_io_ci = io_pp_8[51]; // @[wallace.scala 71:19]
  assign FullAdder_736_io_a = io_pp_9[50]; // @[wallace.scala 69:18]
  assign FullAdder_736_io_b = io_pp_10[49]; // @[wallace.scala 70:18]
  assign FullAdder_736_io_ci = io_pp_11[48]; // @[wallace.scala 71:19]
  assign FullAdder_737_io_a = io_pp_12[47]; // @[wallace.scala 69:18]
  assign FullAdder_737_io_b = io_pp_13[46]; // @[wallace.scala 70:18]
  assign FullAdder_737_io_ci = io_pp_14[45]; // @[wallace.scala 71:19]
  assign FullAdder_738_io_a = io_pp_15[44]; // @[wallace.scala 69:18]
  assign FullAdder_738_io_b = io_pp_16[43]; // @[wallace.scala 70:18]
  assign FullAdder_738_io_ci = io_pp_17[42]; // @[wallace.scala 71:19]
  assign FullAdder_739_io_a = io_pp_18[41]; // @[wallace.scala 69:18]
  assign FullAdder_739_io_b = io_pp_19[40]; // @[wallace.scala 70:18]
  assign FullAdder_739_io_ci = io_pp_20[39]; // @[wallace.scala 71:19]
  assign FullAdder_740_io_a = io_pp_21[38]; // @[wallace.scala 69:18]
  assign FullAdder_740_io_b = io_pp_22[37]; // @[wallace.scala 70:18]
  assign FullAdder_740_io_ci = io_pp_23[36]; // @[wallace.scala 71:19]
  assign FullAdder_741_io_a = io_pp_24[35]; // @[wallace.scala 69:18]
  assign FullAdder_741_io_b = io_pp_25[34]; // @[wallace.scala 70:18]
  assign FullAdder_741_io_ci = io_pp_26[33]; // @[wallace.scala 71:19]
  assign FullAdder_742_io_a = io_pp_27[32]; // @[wallace.scala 69:18]
  assign FullAdder_742_io_b = io_pp_28[31]; // @[wallace.scala 70:18]
  assign FullAdder_742_io_ci = io_pp_29[30]; // @[wallace.scala 71:19]
  assign FullAdder_743_io_a = io_pp_30[29]; // @[wallace.scala 69:18]
  assign FullAdder_743_io_b = io_pp_31[28]; // @[wallace.scala 70:18]
  assign FullAdder_743_io_ci = io_pp_32[27]; // @[wallace.scala 71:19]
  assign FullAdder_744_io_a = io_pp_33[26]; // @[wallace.scala 69:18]
  assign FullAdder_744_io_b = io_pp_34[25]; // @[wallace.scala 70:18]
  assign FullAdder_744_io_ci = io_pp_35[24]; // @[wallace.scala 71:19]
  assign FullAdder_745_io_a = io_pp_36[23]; // @[wallace.scala 69:18]
  assign FullAdder_745_io_b = io_pp_37[22]; // @[wallace.scala 70:18]
  assign FullAdder_745_io_ci = io_pp_38[21]; // @[wallace.scala 71:19]
  assign FullAdder_746_io_a = io_pp_39[20]; // @[wallace.scala 69:18]
  assign FullAdder_746_io_b = io_pp_40[19]; // @[wallace.scala 70:18]
  assign FullAdder_746_io_ci = io_pp_41[18]; // @[wallace.scala 71:19]
  assign FullAdder_747_io_a = io_pp_42[17]; // @[wallace.scala 69:18]
  assign FullAdder_747_io_b = io_pp_43[16]; // @[wallace.scala 70:18]
  assign FullAdder_747_io_ci = io_pp_44[15]; // @[wallace.scala 71:19]
  assign FullAdder_748_io_a = io_pp_45[14]; // @[wallace.scala 69:18]
  assign FullAdder_748_io_b = io_pp_46[13]; // @[wallace.scala 70:18]
  assign FullAdder_748_io_ci = io_pp_47[12]; // @[wallace.scala 71:19]
  assign FullAdder_749_io_a = io_pp_48[11]; // @[wallace.scala 69:18]
  assign FullAdder_749_io_b = io_pp_49[10]; // @[wallace.scala 70:18]
  assign FullAdder_749_io_ci = io_pp_50[9]; // @[wallace.scala 71:19]
  assign FullAdder_750_io_a = io_pp_51[8]; // @[wallace.scala 69:18]
  assign FullAdder_750_io_b = io_pp_52[7]; // @[wallace.scala 70:18]
  assign FullAdder_750_io_ci = io_pp_53[6]; // @[wallace.scala 71:19]
  assign FullAdder_751_io_a = io_pp_54[5]; // @[wallace.scala 69:18]
  assign FullAdder_751_io_b = io_pp_55[4]; // @[wallace.scala 70:18]
  assign FullAdder_751_io_ci = io_pp_56[3]; // @[wallace.scala 71:19]
  assign FullAdder_752_io_a = io_pp_57[2]; // @[wallace.scala 69:18]
  assign FullAdder_752_io_b = io_pp_58[1]; // @[wallace.scala 70:18]
  assign FullAdder_752_io_ci = io_pp_59[0]; // @[wallace.scala 71:19]
  assign FullAdder_753_io_a = io_pp_0[58]; // @[wallace.scala 69:18]
  assign FullAdder_753_io_b = io_pp_1[57]; // @[wallace.scala 70:18]
  assign FullAdder_753_io_ci = io_pp_2[56]; // @[wallace.scala 71:19]
  assign FullAdder_754_io_a = io_pp_3[55]; // @[wallace.scala 69:18]
  assign FullAdder_754_io_b = io_pp_4[54]; // @[wallace.scala 70:18]
  assign FullAdder_754_io_ci = io_pp_5[53]; // @[wallace.scala 71:19]
  assign FullAdder_755_io_a = io_pp_6[52]; // @[wallace.scala 69:18]
  assign FullAdder_755_io_b = io_pp_7[51]; // @[wallace.scala 70:18]
  assign FullAdder_755_io_ci = io_pp_8[50]; // @[wallace.scala 71:19]
  assign FullAdder_756_io_a = io_pp_9[49]; // @[wallace.scala 69:18]
  assign FullAdder_756_io_b = io_pp_10[48]; // @[wallace.scala 70:18]
  assign FullAdder_756_io_ci = io_pp_11[47]; // @[wallace.scala 71:19]
  assign FullAdder_757_io_a = io_pp_12[46]; // @[wallace.scala 69:18]
  assign FullAdder_757_io_b = io_pp_13[45]; // @[wallace.scala 70:18]
  assign FullAdder_757_io_ci = io_pp_14[44]; // @[wallace.scala 71:19]
  assign FullAdder_758_io_a = io_pp_15[43]; // @[wallace.scala 69:18]
  assign FullAdder_758_io_b = io_pp_16[42]; // @[wallace.scala 70:18]
  assign FullAdder_758_io_ci = io_pp_17[41]; // @[wallace.scala 71:19]
  assign FullAdder_759_io_a = io_pp_18[40]; // @[wallace.scala 69:18]
  assign FullAdder_759_io_b = io_pp_19[39]; // @[wallace.scala 70:18]
  assign FullAdder_759_io_ci = io_pp_20[38]; // @[wallace.scala 71:19]
  assign FullAdder_760_io_a = io_pp_21[37]; // @[wallace.scala 69:18]
  assign FullAdder_760_io_b = io_pp_22[36]; // @[wallace.scala 70:18]
  assign FullAdder_760_io_ci = io_pp_23[35]; // @[wallace.scala 71:19]
  assign FullAdder_761_io_a = io_pp_24[34]; // @[wallace.scala 69:18]
  assign FullAdder_761_io_b = io_pp_25[33]; // @[wallace.scala 70:18]
  assign FullAdder_761_io_ci = io_pp_26[32]; // @[wallace.scala 71:19]
  assign FullAdder_762_io_a = io_pp_27[31]; // @[wallace.scala 69:18]
  assign FullAdder_762_io_b = io_pp_28[30]; // @[wallace.scala 70:18]
  assign FullAdder_762_io_ci = io_pp_29[29]; // @[wallace.scala 71:19]
  assign FullAdder_763_io_a = io_pp_30[28]; // @[wallace.scala 69:18]
  assign FullAdder_763_io_b = io_pp_31[27]; // @[wallace.scala 70:18]
  assign FullAdder_763_io_ci = io_pp_32[26]; // @[wallace.scala 71:19]
  assign FullAdder_764_io_a = io_pp_33[25]; // @[wallace.scala 69:18]
  assign FullAdder_764_io_b = io_pp_34[24]; // @[wallace.scala 70:18]
  assign FullAdder_764_io_ci = io_pp_35[23]; // @[wallace.scala 71:19]
  assign FullAdder_765_io_a = io_pp_36[22]; // @[wallace.scala 69:18]
  assign FullAdder_765_io_b = io_pp_37[21]; // @[wallace.scala 70:18]
  assign FullAdder_765_io_ci = io_pp_38[20]; // @[wallace.scala 71:19]
  assign FullAdder_766_io_a = io_pp_39[19]; // @[wallace.scala 69:18]
  assign FullAdder_766_io_b = io_pp_40[18]; // @[wallace.scala 70:18]
  assign FullAdder_766_io_ci = io_pp_41[17]; // @[wallace.scala 71:19]
  assign FullAdder_767_io_a = io_pp_42[16]; // @[wallace.scala 69:18]
  assign FullAdder_767_io_b = io_pp_43[15]; // @[wallace.scala 70:18]
  assign FullAdder_767_io_ci = io_pp_44[14]; // @[wallace.scala 71:19]
  assign FullAdder_768_io_a = io_pp_45[13]; // @[wallace.scala 69:18]
  assign FullAdder_768_io_b = io_pp_46[12]; // @[wallace.scala 70:18]
  assign FullAdder_768_io_ci = io_pp_47[11]; // @[wallace.scala 71:19]
  assign FullAdder_769_io_a = io_pp_48[10]; // @[wallace.scala 69:18]
  assign FullAdder_769_io_b = io_pp_49[9]; // @[wallace.scala 70:18]
  assign FullAdder_769_io_ci = io_pp_50[8]; // @[wallace.scala 71:19]
  assign FullAdder_770_io_a = io_pp_51[7]; // @[wallace.scala 69:18]
  assign FullAdder_770_io_b = io_pp_52[6]; // @[wallace.scala 70:18]
  assign FullAdder_770_io_ci = io_pp_53[5]; // @[wallace.scala 71:19]
  assign FullAdder_771_io_a = io_pp_54[4]; // @[wallace.scala 69:18]
  assign FullAdder_771_io_b = io_pp_55[3]; // @[wallace.scala 70:18]
  assign FullAdder_771_io_ci = io_pp_56[2]; // @[wallace.scala 71:19]
  assign HalfAdder_19_io_a = io_pp_57[1]; // @[wallace.scala 59:18]
  assign HalfAdder_19_io_b = io_pp_58[0]; // @[wallace.scala 60:18]
  assign FullAdder_772_io_a = io_pp_0[57]; // @[wallace.scala 69:18]
  assign FullAdder_772_io_b = io_pp_1[56]; // @[wallace.scala 70:18]
  assign FullAdder_772_io_ci = io_pp_2[55]; // @[wallace.scala 71:19]
  assign FullAdder_773_io_a = io_pp_3[54]; // @[wallace.scala 69:18]
  assign FullAdder_773_io_b = io_pp_4[53]; // @[wallace.scala 70:18]
  assign FullAdder_773_io_ci = io_pp_5[52]; // @[wallace.scala 71:19]
  assign FullAdder_774_io_a = io_pp_6[51]; // @[wallace.scala 69:18]
  assign FullAdder_774_io_b = io_pp_7[50]; // @[wallace.scala 70:18]
  assign FullAdder_774_io_ci = io_pp_8[49]; // @[wallace.scala 71:19]
  assign FullAdder_775_io_a = io_pp_9[48]; // @[wallace.scala 69:18]
  assign FullAdder_775_io_b = io_pp_10[47]; // @[wallace.scala 70:18]
  assign FullAdder_775_io_ci = io_pp_11[46]; // @[wallace.scala 71:19]
  assign FullAdder_776_io_a = io_pp_12[45]; // @[wallace.scala 69:18]
  assign FullAdder_776_io_b = io_pp_13[44]; // @[wallace.scala 70:18]
  assign FullAdder_776_io_ci = io_pp_14[43]; // @[wallace.scala 71:19]
  assign FullAdder_777_io_a = io_pp_15[42]; // @[wallace.scala 69:18]
  assign FullAdder_777_io_b = io_pp_16[41]; // @[wallace.scala 70:18]
  assign FullAdder_777_io_ci = io_pp_17[40]; // @[wallace.scala 71:19]
  assign FullAdder_778_io_a = io_pp_18[39]; // @[wallace.scala 69:18]
  assign FullAdder_778_io_b = io_pp_19[38]; // @[wallace.scala 70:18]
  assign FullAdder_778_io_ci = io_pp_20[37]; // @[wallace.scala 71:19]
  assign FullAdder_779_io_a = io_pp_21[36]; // @[wallace.scala 69:18]
  assign FullAdder_779_io_b = io_pp_22[35]; // @[wallace.scala 70:18]
  assign FullAdder_779_io_ci = io_pp_23[34]; // @[wallace.scala 71:19]
  assign FullAdder_780_io_a = io_pp_24[33]; // @[wallace.scala 69:18]
  assign FullAdder_780_io_b = io_pp_25[32]; // @[wallace.scala 70:18]
  assign FullAdder_780_io_ci = io_pp_26[31]; // @[wallace.scala 71:19]
  assign FullAdder_781_io_a = io_pp_27[30]; // @[wallace.scala 69:18]
  assign FullAdder_781_io_b = io_pp_28[29]; // @[wallace.scala 70:18]
  assign FullAdder_781_io_ci = io_pp_29[28]; // @[wallace.scala 71:19]
  assign FullAdder_782_io_a = io_pp_30[27]; // @[wallace.scala 69:18]
  assign FullAdder_782_io_b = io_pp_31[26]; // @[wallace.scala 70:18]
  assign FullAdder_782_io_ci = io_pp_32[25]; // @[wallace.scala 71:19]
  assign FullAdder_783_io_a = io_pp_33[24]; // @[wallace.scala 69:18]
  assign FullAdder_783_io_b = io_pp_34[23]; // @[wallace.scala 70:18]
  assign FullAdder_783_io_ci = io_pp_35[22]; // @[wallace.scala 71:19]
  assign FullAdder_784_io_a = io_pp_36[21]; // @[wallace.scala 69:18]
  assign FullAdder_784_io_b = io_pp_37[20]; // @[wallace.scala 70:18]
  assign FullAdder_784_io_ci = io_pp_38[19]; // @[wallace.scala 71:19]
  assign FullAdder_785_io_a = io_pp_39[18]; // @[wallace.scala 69:18]
  assign FullAdder_785_io_b = io_pp_40[17]; // @[wallace.scala 70:18]
  assign FullAdder_785_io_ci = io_pp_41[16]; // @[wallace.scala 71:19]
  assign FullAdder_786_io_a = io_pp_42[15]; // @[wallace.scala 69:18]
  assign FullAdder_786_io_b = io_pp_43[14]; // @[wallace.scala 70:18]
  assign FullAdder_786_io_ci = io_pp_44[13]; // @[wallace.scala 71:19]
  assign FullAdder_787_io_a = io_pp_45[12]; // @[wallace.scala 69:18]
  assign FullAdder_787_io_b = io_pp_46[11]; // @[wallace.scala 70:18]
  assign FullAdder_787_io_ci = io_pp_47[10]; // @[wallace.scala 71:19]
  assign FullAdder_788_io_a = io_pp_48[9]; // @[wallace.scala 69:18]
  assign FullAdder_788_io_b = io_pp_49[8]; // @[wallace.scala 70:18]
  assign FullAdder_788_io_ci = io_pp_50[7]; // @[wallace.scala 71:19]
  assign FullAdder_789_io_a = io_pp_51[6]; // @[wallace.scala 69:18]
  assign FullAdder_789_io_b = io_pp_52[5]; // @[wallace.scala 70:18]
  assign FullAdder_789_io_ci = io_pp_53[4]; // @[wallace.scala 71:19]
  assign FullAdder_790_io_a = io_pp_54[3]; // @[wallace.scala 69:18]
  assign FullAdder_790_io_b = io_pp_55[2]; // @[wallace.scala 70:18]
  assign FullAdder_790_io_ci = io_pp_56[1]; // @[wallace.scala 71:19]
  assign FullAdder_791_io_a = io_pp_0[56]; // @[wallace.scala 69:18]
  assign FullAdder_791_io_b = io_pp_1[55]; // @[wallace.scala 70:18]
  assign FullAdder_791_io_ci = io_pp_2[54]; // @[wallace.scala 71:19]
  assign FullAdder_792_io_a = io_pp_3[53]; // @[wallace.scala 69:18]
  assign FullAdder_792_io_b = io_pp_4[52]; // @[wallace.scala 70:18]
  assign FullAdder_792_io_ci = io_pp_5[51]; // @[wallace.scala 71:19]
  assign FullAdder_793_io_a = io_pp_6[50]; // @[wallace.scala 69:18]
  assign FullAdder_793_io_b = io_pp_7[49]; // @[wallace.scala 70:18]
  assign FullAdder_793_io_ci = io_pp_8[48]; // @[wallace.scala 71:19]
  assign FullAdder_794_io_a = io_pp_9[47]; // @[wallace.scala 69:18]
  assign FullAdder_794_io_b = io_pp_10[46]; // @[wallace.scala 70:18]
  assign FullAdder_794_io_ci = io_pp_11[45]; // @[wallace.scala 71:19]
  assign FullAdder_795_io_a = io_pp_12[44]; // @[wallace.scala 69:18]
  assign FullAdder_795_io_b = io_pp_13[43]; // @[wallace.scala 70:18]
  assign FullAdder_795_io_ci = io_pp_14[42]; // @[wallace.scala 71:19]
  assign FullAdder_796_io_a = io_pp_15[41]; // @[wallace.scala 69:18]
  assign FullAdder_796_io_b = io_pp_16[40]; // @[wallace.scala 70:18]
  assign FullAdder_796_io_ci = io_pp_17[39]; // @[wallace.scala 71:19]
  assign FullAdder_797_io_a = io_pp_18[38]; // @[wallace.scala 69:18]
  assign FullAdder_797_io_b = io_pp_19[37]; // @[wallace.scala 70:18]
  assign FullAdder_797_io_ci = io_pp_20[36]; // @[wallace.scala 71:19]
  assign FullAdder_798_io_a = io_pp_21[35]; // @[wallace.scala 69:18]
  assign FullAdder_798_io_b = io_pp_22[34]; // @[wallace.scala 70:18]
  assign FullAdder_798_io_ci = io_pp_23[33]; // @[wallace.scala 71:19]
  assign FullAdder_799_io_a = io_pp_24[32]; // @[wallace.scala 69:18]
  assign FullAdder_799_io_b = io_pp_25[31]; // @[wallace.scala 70:18]
  assign FullAdder_799_io_ci = io_pp_26[30]; // @[wallace.scala 71:19]
  assign FullAdder_800_io_a = io_pp_27[29]; // @[wallace.scala 69:18]
  assign FullAdder_800_io_b = io_pp_28[28]; // @[wallace.scala 70:18]
  assign FullAdder_800_io_ci = io_pp_29[27]; // @[wallace.scala 71:19]
  assign FullAdder_801_io_a = io_pp_30[26]; // @[wallace.scala 69:18]
  assign FullAdder_801_io_b = io_pp_31[25]; // @[wallace.scala 70:18]
  assign FullAdder_801_io_ci = io_pp_32[24]; // @[wallace.scala 71:19]
  assign FullAdder_802_io_a = io_pp_33[23]; // @[wallace.scala 69:18]
  assign FullAdder_802_io_b = io_pp_34[22]; // @[wallace.scala 70:18]
  assign FullAdder_802_io_ci = io_pp_35[21]; // @[wallace.scala 71:19]
  assign FullAdder_803_io_a = io_pp_36[20]; // @[wallace.scala 69:18]
  assign FullAdder_803_io_b = io_pp_37[19]; // @[wallace.scala 70:18]
  assign FullAdder_803_io_ci = io_pp_38[18]; // @[wallace.scala 71:19]
  assign FullAdder_804_io_a = io_pp_39[17]; // @[wallace.scala 69:18]
  assign FullAdder_804_io_b = io_pp_40[16]; // @[wallace.scala 70:18]
  assign FullAdder_804_io_ci = io_pp_41[15]; // @[wallace.scala 71:19]
  assign FullAdder_805_io_a = io_pp_42[14]; // @[wallace.scala 69:18]
  assign FullAdder_805_io_b = io_pp_43[13]; // @[wallace.scala 70:18]
  assign FullAdder_805_io_ci = io_pp_44[12]; // @[wallace.scala 71:19]
  assign FullAdder_806_io_a = io_pp_45[11]; // @[wallace.scala 69:18]
  assign FullAdder_806_io_b = io_pp_46[10]; // @[wallace.scala 70:18]
  assign FullAdder_806_io_ci = io_pp_47[9]; // @[wallace.scala 71:19]
  assign FullAdder_807_io_a = io_pp_48[8]; // @[wallace.scala 69:18]
  assign FullAdder_807_io_b = io_pp_49[7]; // @[wallace.scala 70:18]
  assign FullAdder_807_io_ci = io_pp_50[6]; // @[wallace.scala 71:19]
  assign FullAdder_808_io_a = io_pp_51[5]; // @[wallace.scala 69:18]
  assign FullAdder_808_io_b = io_pp_52[4]; // @[wallace.scala 70:18]
  assign FullAdder_808_io_ci = io_pp_53[3]; // @[wallace.scala 71:19]
  assign FullAdder_809_io_a = io_pp_54[2]; // @[wallace.scala 69:18]
  assign FullAdder_809_io_b = io_pp_55[1]; // @[wallace.scala 70:18]
  assign FullAdder_809_io_ci = io_pp_56[0]; // @[wallace.scala 71:19]
  assign FullAdder_810_io_a = io_pp_0[55]; // @[wallace.scala 69:18]
  assign FullAdder_810_io_b = io_pp_1[54]; // @[wallace.scala 70:18]
  assign FullAdder_810_io_ci = io_pp_2[53]; // @[wallace.scala 71:19]
  assign FullAdder_811_io_a = io_pp_3[52]; // @[wallace.scala 69:18]
  assign FullAdder_811_io_b = io_pp_4[51]; // @[wallace.scala 70:18]
  assign FullAdder_811_io_ci = io_pp_5[50]; // @[wallace.scala 71:19]
  assign FullAdder_812_io_a = io_pp_6[49]; // @[wallace.scala 69:18]
  assign FullAdder_812_io_b = io_pp_7[48]; // @[wallace.scala 70:18]
  assign FullAdder_812_io_ci = io_pp_8[47]; // @[wallace.scala 71:19]
  assign FullAdder_813_io_a = io_pp_9[46]; // @[wallace.scala 69:18]
  assign FullAdder_813_io_b = io_pp_10[45]; // @[wallace.scala 70:18]
  assign FullAdder_813_io_ci = io_pp_11[44]; // @[wallace.scala 71:19]
  assign FullAdder_814_io_a = io_pp_12[43]; // @[wallace.scala 69:18]
  assign FullAdder_814_io_b = io_pp_13[42]; // @[wallace.scala 70:18]
  assign FullAdder_814_io_ci = io_pp_14[41]; // @[wallace.scala 71:19]
  assign FullAdder_815_io_a = io_pp_15[40]; // @[wallace.scala 69:18]
  assign FullAdder_815_io_b = io_pp_16[39]; // @[wallace.scala 70:18]
  assign FullAdder_815_io_ci = io_pp_17[38]; // @[wallace.scala 71:19]
  assign FullAdder_816_io_a = io_pp_18[37]; // @[wallace.scala 69:18]
  assign FullAdder_816_io_b = io_pp_19[36]; // @[wallace.scala 70:18]
  assign FullAdder_816_io_ci = io_pp_20[35]; // @[wallace.scala 71:19]
  assign FullAdder_817_io_a = io_pp_21[34]; // @[wallace.scala 69:18]
  assign FullAdder_817_io_b = io_pp_22[33]; // @[wallace.scala 70:18]
  assign FullAdder_817_io_ci = io_pp_23[32]; // @[wallace.scala 71:19]
  assign FullAdder_818_io_a = io_pp_24[31]; // @[wallace.scala 69:18]
  assign FullAdder_818_io_b = io_pp_25[30]; // @[wallace.scala 70:18]
  assign FullAdder_818_io_ci = io_pp_26[29]; // @[wallace.scala 71:19]
  assign FullAdder_819_io_a = io_pp_27[28]; // @[wallace.scala 69:18]
  assign FullAdder_819_io_b = io_pp_28[27]; // @[wallace.scala 70:18]
  assign FullAdder_819_io_ci = io_pp_29[26]; // @[wallace.scala 71:19]
  assign FullAdder_820_io_a = io_pp_30[25]; // @[wallace.scala 69:18]
  assign FullAdder_820_io_b = io_pp_31[24]; // @[wallace.scala 70:18]
  assign FullAdder_820_io_ci = io_pp_32[23]; // @[wallace.scala 71:19]
  assign FullAdder_821_io_a = io_pp_33[22]; // @[wallace.scala 69:18]
  assign FullAdder_821_io_b = io_pp_34[21]; // @[wallace.scala 70:18]
  assign FullAdder_821_io_ci = io_pp_35[20]; // @[wallace.scala 71:19]
  assign FullAdder_822_io_a = io_pp_36[19]; // @[wallace.scala 69:18]
  assign FullAdder_822_io_b = io_pp_37[18]; // @[wallace.scala 70:18]
  assign FullAdder_822_io_ci = io_pp_38[17]; // @[wallace.scala 71:19]
  assign FullAdder_823_io_a = io_pp_39[16]; // @[wallace.scala 69:18]
  assign FullAdder_823_io_b = io_pp_40[15]; // @[wallace.scala 70:18]
  assign FullAdder_823_io_ci = io_pp_41[14]; // @[wallace.scala 71:19]
  assign FullAdder_824_io_a = io_pp_42[13]; // @[wallace.scala 69:18]
  assign FullAdder_824_io_b = io_pp_43[12]; // @[wallace.scala 70:18]
  assign FullAdder_824_io_ci = io_pp_44[11]; // @[wallace.scala 71:19]
  assign FullAdder_825_io_a = io_pp_45[10]; // @[wallace.scala 69:18]
  assign FullAdder_825_io_b = io_pp_46[9]; // @[wallace.scala 70:18]
  assign FullAdder_825_io_ci = io_pp_47[8]; // @[wallace.scala 71:19]
  assign FullAdder_826_io_a = io_pp_48[7]; // @[wallace.scala 69:18]
  assign FullAdder_826_io_b = io_pp_49[6]; // @[wallace.scala 70:18]
  assign FullAdder_826_io_ci = io_pp_50[5]; // @[wallace.scala 71:19]
  assign FullAdder_827_io_a = io_pp_51[4]; // @[wallace.scala 69:18]
  assign FullAdder_827_io_b = io_pp_52[3]; // @[wallace.scala 70:18]
  assign FullAdder_827_io_ci = io_pp_53[2]; // @[wallace.scala 71:19]
  assign FullAdder_828_io_a = io_pp_0[54]; // @[wallace.scala 69:18]
  assign FullAdder_828_io_b = io_pp_1[53]; // @[wallace.scala 70:18]
  assign FullAdder_828_io_ci = io_pp_2[52]; // @[wallace.scala 71:19]
  assign FullAdder_829_io_a = io_pp_3[51]; // @[wallace.scala 69:18]
  assign FullAdder_829_io_b = io_pp_4[50]; // @[wallace.scala 70:18]
  assign FullAdder_829_io_ci = io_pp_5[49]; // @[wallace.scala 71:19]
  assign FullAdder_830_io_a = io_pp_6[48]; // @[wallace.scala 69:18]
  assign FullAdder_830_io_b = io_pp_7[47]; // @[wallace.scala 70:18]
  assign FullAdder_830_io_ci = io_pp_8[46]; // @[wallace.scala 71:19]
  assign FullAdder_831_io_a = io_pp_9[45]; // @[wallace.scala 69:18]
  assign FullAdder_831_io_b = io_pp_10[44]; // @[wallace.scala 70:18]
  assign FullAdder_831_io_ci = io_pp_11[43]; // @[wallace.scala 71:19]
  assign FullAdder_832_io_a = io_pp_12[42]; // @[wallace.scala 69:18]
  assign FullAdder_832_io_b = io_pp_13[41]; // @[wallace.scala 70:18]
  assign FullAdder_832_io_ci = io_pp_14[40]; // @[wallace.scala 71:19]
  assign FullAdder_833_io_a = io_pp_15[39]; // @[wallace.scala 69:18]
  assign FullAdder_833_io_b = io_pp_16[38]; // @[wallace.scala 70:18]
  assign FullAdder_833_io_ci = io_pp_17[37]; // @[wallace.scala 71:19]
  assign FullAdder_834_io_a = io_pp_18[36]; // @[wallace.scala 69:18]
  assign FullAdder_834_io_b = io_pp_19[35]; // @[wallace.scala 70:18]
  assign FullAdder_834_io_ci = io_pp_20[34]; // @[wallace.scala 71:19]
  assign FullAdder_835_io_a = io_pp_21[33]; // @[wallace.scala 69:18]
  assign FullAdder_835_io_b = io_pp_22[32]; // @[wallace.scala 70:18]
  assign FullAdder_835_io_ci = io_pp_23[31]; // @[wallace.scala 71:19]
  assign FullAdder_836_io_a = io_pp_24[30]; // @[wallace.scala 69:18]
  assign FullAdder_836_io_b = io_pp_25[29]; // @[wallace.scala 70:18]
  assign FullAdder_836_io_ci = io_pp_26[28]; // @[wallace.scala 71:19]
  assign FullAdder_837_io_a = io_pp_27[27]; // @[wallace.scala 69:18]
  assign FullAdder_837_io_b = io_pp_28[26]; // @[wallace.scala 70:18]
  assign FullAdder_837_io_ci = io_pp_29[25]; // @[wallace.scala 71:19]
  assign FullAdder_838_io_a = io_pp_30[24]; // @[wallace.scala 69:18]
  assign FullAdder_838_io_b = io_pp_31[23]; // @[wallace.scala 70:18]
  assign FullAdder_838_io_ci = io_pp_32[22]; // @[wallace.scala 71:19]
  assign FullAdder_839_io_a = io_pp_33[21]; // @[wallace.scala 69:18]
  assign FullAdder_839_io_b = io_pp_34[20]; // @[wallace.scala 70:18]
  assign FullAdder_839_io_ci = io_pp_35[19]; // @[wallace.scala 71:19]
  assign FullAdder_840_io_a = io_pp_36[18]; // @[wallace.scala 69:18]
  assign FullAdder_840_io_b = io_pp_37[17]; // @[wallace.scala 70:18]
  assign FullAdder_840_io_ci = io_pp_38[16]; // @[wallace.scala 71:19]
  assign FullAdder_841_io_a = io_pp_39[15]; // @[wallace.scala 69:18]
  assign FullAdder_841_io_b = io_pp_40[14]; // @[wallace.scala 70:18]
  assign FullAdder_841_io_ci = io_pp_41[13]; // @[wallace.scala 71:19]
  assign FullAdder_842_io_a = io_pp_42[12]; // @[wallace.scala 69:18]
  assign FullAdder_842_io_b = io_pp_43[11]; // @[wallace.scala 70:18]
  assign FullAdder_842_io_ci = io_pp_44[10]; // @[wallace.scala 71:19]
  assign FullAdder_843_io_a = io_pp_45[9]; // @[wallace.scala 69:18]
  assign FullAdder_843_io_b = io_pp_46[8]; // @[wallace.scala 70:18]
  assign FullAdder_843_io_ci = io_pp_47[7]; // @[wallace.scala 71:19]
  assign FullAdder_844_io_a = io_pp_48[6]; // @[wallace.scala 69:18]
  assign FullAdder_844_io_b = io_pp_49[5]; // @[wallace.scala 70:18]
  assign FullAdder_844_io_ci = io_pp_50[4]; // @[wallace.scala 71:19]
  assign FullAdder_845_io_a = io_pp_51[3]; // @[wallace.scala 69:18]
  assign FullAdder_845_io_b = io_pp_52[2]; // @[wallace.scala 70:18]
  assign FullAdder_845_io_ci = io_pp_53[1]; // @[wallace.scala 71:19]
  assign FullAdder_846_io_a = io_pp_0[53]; // @[wallace.scala 69:18]
  assign FullAdder_846_io_b = io_pp_1[52]; // @[wallace.scala 70:18]
  assign FullAdder_846_io_ci = io_pp_2[51]; // @[wallace.scala 71:19]
  assign FullAdder_847_io_a = io_pp_3[50]; // @[wallace.scala 69:18]
  assign FullAdder_847_io_b = io_pp_4[49]; // @[wallace.scala 70:18]
  assign FullAdder_847_io_ci = io_pp_5[48]; // @[wallace.scala 71:19]
  assign FullAdder_848_io_a = io_pp_6[47]; // @[wallace.scala 69:18]
  assign FullAdder_848_io_b = io_pp_7[46]; // @[wallace.scala 70:18]
  assign FullAdder_848_io_ci = io_pp_8[45]; // @[wallace.scala 71:19]
  assign FullAdder_849_io_a = io_pp_9[44]; // @[wallace.scala 69:18]
  assign FullAdder_849_io_b = io_pp_10[43]; // @[wallace.scala 70:18]
  assign FullAdder_849_io_ci = io_pp_11[42]; // @[wallace.scala 71:19]
  assign FullAdder_850_io_a = io_pp_12[41]; // @[wallace.scala 69:18]
  assign FullAdder_850_io_b = io_pp_13[40]; // @[wallace.scala 70:18]
  assign FullAdder_850_io_ci = io_pp_14[39]; // @[wallace.scala 71:19]
  assign FullAdder_851_io_a = io_pp_15[38]; // @[wallace.scala 69:18]
  assign FullAdder_851_io_b = io_pp_16[37]; // @[wallace.scala 70:18]
  assign FullAdder_851_io_ci = io_pp_17[36]; // @[wallace.scala 71:19]
  assign FullAdder_852_io_a = io_pp_18[35]; // @[wallace.scala 69:18]
  assign FullAdder_852_io_b = io_pp_19[34]; // @[wallace.scala 70:18]
  assign FullAdder_852_io_ci = io_pp_20[33]; // @[wallace.scala 71:19]
  assign FullAdder_853_io_a = io_pp_21[32]; // @[wallace.scala 69:18]
  assign FullAdder_853_io_b = io_pp_22[31]; // @[wallace.scala 70:18]
  assign FullAdder_853_io_ci = io_pp_23[30]; // @[wallace.scala 71:19]
  assign FullAdder_854_io_a = io_pp_24[29]; // @[wallace.scala 69:18]
  assign FullAdder_854_io_b = io_pp_25[28]; // @[wallace.scala 70:18]
  assign FullAdder_854_io_ci = io_pp_26[27]; // @[wallace.scala 71:19]
  assign FullAdder_855_io_a = io_pp_27[26]; // @[wallace.scala 69:18]
  assign FullAdder_855_io_b = io_pp_28[25]; // @[wallace.scala 70:18]
  assign FullAdder_855_io_ci = io_pp_29[24]; // @[wallace.scala 71:19]
  assign FullAdder_856_io_a = io_pp_30[23]; // @[wallace.scala 69:18]
  assign FullAdder_856_io_b = io_pp_31[22]; // @[wallace.scala 70:18]
  assign FullAdder_856_io_ci = io_pp_32[21]; // @[wallace.scala 71:19]
  assign FullAdder_857_io_a = io_pp_33[20]; // @[wallace.scala 69:18]
  assign FullAdder_857_io_b = io_pp_34[19]; // @[wallace.scala 70:18]
  assign FullAdder_857_io_ci = io_pp_35[18]; // @[wallace.scala 71:19]
  assign FullAdder_858_io_a = io_pp_36[17]; // @[wallace.scala 69:18]
  assign FullAdder_858_io_b = io_pp_37[16]; // @[wallace.scala 70:18]
  assign FullAdder_858_io_ci = io_pp_38[15]; // @[wallace.scala 71:19]
  assign FullAdder_859_io_a = io_pp_39[14]; // @[wallace.scala 69:18]
  assign FullAdder_859_io_b = io_pp_40[13]; // @[wallace.scala 70:18]
  assign FullAdder_859_io_ci = io_pp_41[12]; // @[wallace.scala 71:19]
  assign FullAdder_860_io_a = io_pp_42[11]; // @[wallace.scala 69:18]
  assign FullAdder_860_io_b = io_pp_43[10]; // @[wallace.scala 70:18]
  assign FullAdder_860_io_ci = io_pp_44[9]; // @[wallace.scala 71:19]
  assign FullAdder_861_io_a = io_pp_45[8]; // @[wallace.scala 69:18]
  assign FullAdder_861_io_b = io_pp_46[7]; // @[wallace.scala 70:18]
  assign FullAdder_861_io_ci = io_pp_47[6]; // @[wallace.scala 71:19]
  assign FullAdder_862_io_a = io_pp_48[5]; // @[wallace.scala 69:18]
  assign FullAdder_862_io_b = io_pp_49[4]; // @[wallace.scala 70:18]
  assign FullAdder_862_io_ci = io_pp_50[3]; // @[wallace.scala 71:19]
  assign FullAdder_863_io_a = io_pp_51[2]; // @[wallace.scala 69:18]
  assign FullAdder_863_io_b = io_pp_52[1]; // @[wallace.scala 70:18]
  assign FullAdder_863_io_ci = io_pp_53[0]; // @[wallace.scala 71:19]
  assign FullAdder_864_io_a = io_pp_0[52]; // @[wallace.scala 69:18]
  assign FullAdder_864_io_b = io_pp_1[51]; // @[wallace.scala 70:18]
  assign FullAdder_864_io_ci = io_pp_2[50]; // @[wallace.scala 71:19]
  assign FullAdder_865_io_a = io_pp_3[49]; // @[wallace.scala 69:18]
  assign FullAdder_865_io_b = io_pp_4[48]; // @[wallace.scala 70:18]
  assign FullAdder_865_io_ci = io_pp_5[47]; // @[wallace.scala 71:19]
  assign FullAdder_866_io_a = io_pp_6[46]; // @[wallace.scala 69:18]
  assign FullAdder_866_io_b = io_pp_7[45]; // @[wallace.scala 70:18]
  assign FullAdder_866_io_ci = io_pp_8[44]; // @[wallace.scala 71:19]
  assign FullAdder_867_io_a = io_pp_9[43]; // @[wallace.scala 69:18]
  assign FullAdder_867_io_b = io_pp_10[42]; // @[wallace.scala 70:18]
  assign FullAdder_867_io_ci = io_pp_11[41]; // @[wallace.scala 71:19]
  assign FullAdder_868_io_a = io_pp_12[40]; // @[wallace.scala 69:18]
  assign FullAdder_868_io_b = io_pp_13[39]; // @[wallace.scala 70:18]
  assign FullAdder_868_io_ci = io_pp_14[38]; // @[wallace.scala 71:19]
  assign FullAdder_869_io_a = io_pp_15[37]; // @[wallace.scala 69:18]
  assign FullAdder_869_io_b = io_pp_16[36]; // @[wallace.scala 70:18]
  assign FullAdder_869_io_ci = io_pp_17[35]; // @[wallace.scala 71:19]
  assign FullAdder_870_io_a = io_pp_18[34]; // @[wallace.scala 69:18]
  assign FullAdder_870_io_b = io_pp_19[33]; // @[wallace.scala 70:18]
  assign FullAdder_870_io_ci = io_pp_20[32]; // @[wallace.scala 71:19]
  assign FullAdder_871_io_a = io_pp_21[31]; // @[wallace.scala 69:18]
  assign FullAdder_871_io_b = io_pp_22[30]; // @[wallace.scala 70:18]
  assign FullAdder_871_io_ci = io_pp_23[29]; // @[wallace.scala 71:19]
  assign FullAdder_872_io_a = io_pp_24[28]; // @[wallace.scala 69:18]
  assign FullAdder_872_io_b = io_pp_25[27]; // @[wallace.scala 70:18]
  assign FullAdder_872_io_ci = io_pp_26[26]; // @[wallace.scala 71:19]
  assign FullAdder_873_io_a = io_pp_27[25]; // @[wallace.scala 69:18]
  assign FullAdder_873_io_b = io_pp_28[24]; // @[wallace.scala 70:18]
  assign FullAdder_873_io_ci = io_pp_29[23]; // @[wallace.scala 71:19]
  assign FullAdder_874_io_a = io_pp_30[22]; // @[wallace.scala 69:18]
  assign FullAdder_874_io_b = io_pp_31[21]; // @[wallace.scala 70:18]
  assign FullAdder_874_io_ci = io_pp_32[20]; // @[wallace.scala 71:19]
  assign FullAdder_875_io_a = io_pp_33[19]; // @[wallace.scala 69:18]
  assign FullAdder_875_io_b = io_pp_34[18]; // @[wallace.scala 70:18]
  assign FullAdder_875_io_ci = io_pp_35[17]; // @[wallace.scala 71:19]
  assign FullAdder_876_io_a = io_pp_36[16]; // @[wallace.scala 69:18]
  assign FullAdder_876_io_b = io_pp_37[15]; // @[wallace.scala 70:18]
  assign FullAdder_876_io_ci = io_pp_38[14]; // @[wallace.scala 71:19]
  assign FullAdder_877_io_a = io_pp_39[13]; // @[wallace.scala 69:18]
  assign FullAdder_877_io_b = io_pp_40[12]; // @[wallace.scala 70:18]
  assign FullAdder_877_io_ci = io_pp_41[11]; // @[wallace.scala 71:19]
  assign FullAdder_878_io_a = io_pp_42[10]; // @[wallace.scala 69:18]
  assign FullAdder_878_io_b = io_pp_43[9]; // @[wallace.scala 70:18]
  assign FullAdder_878_io_ci = io_pp_44[8]; // @[wallace.scala 71:19]
  assign FullAdder_879_io_a = io_pp_45[7]; // @[wallace.scala 69:18]
  assign FullAdder_879_io_b = io_pp_46[6]; // @[wallace.scala 70:18]
  assign FullAdder_879_io_ci = io_pp_47[5]; // @[wallace.scala 71:19]
  assign FullAdder_880_io_a = io_pp_48[4]; // @[wallace.scala 69:18]
  assign FullAdder_880_io_b = io_pp_49[3]; // @[wallace.scala 70:18]
  assign FullAdder_880_io_ci = io_pp_50[2]; // @[wallace.scala 71:19]
  assign HalfAdder_20_io_a = io_pp_51[1]; // @[wallace.scala 59:18]
  assign HalfAdder_20_io_b = io_pp_52[0]; // @[wallace.scala 60:18]
  assign FullAdder_881_io_a = io_pp_0[51]; // @[wallace.scala 69:18]
  assign FullAdder_881_io_b = io_pp_1[50]; // @[wallace.scala 70:18]
  assign FullAdder_881_io_ci = io_pp_2[49]; // @[wallace.scala 71:19]
  assign FullAdder_882_io_a = io_pp_3[48]; // @[wallace.scala 69:18]
  assign FullAdder_882_io_b = io_pp_4[47]; // @[wallace.scala 70:18]
  assign FullAdder_882_io_ci = io_pp_5[46]; // @[wallace.scala 71:19]
  assign FullAdder_883_io_a = io_pp_6[45]; // @[wallace.scala 69:18]
  assign FullAdder_883_io_b = io_pp_7[44]; // @[wallace.scala 70:18]
  assign FullAdder_883_io_ci = io_pp_8[43]; // @[wallace.scala 71:19]
  assign FullAdder_884_io_a = io_pp_9[42]; // @[wallace.scala 69:18]
  assign FullAdder_884_io_b = io_pp_10[41]; // @[wallace.scala 70:18]
  assign FullAdder_884_io_ci = io_pp_11[40]; // @[wallace.scala 71:19]
  assign FullAdder_885_io_a = io_pp_12[39]; // @[wallace.scala 69:18]
  assign FullAdder_885_io_b = io_pp_13[38]; // @[wallace.scala 70:18]
  assign FullAdder_885_io_ci = io_pp_14[37]; // @[wallace.scala 71:19]
  assign FullAdder_886_io_a = io_pp_15[36]; // @[wallace.scala 69:18]
  assign FullAdder_886_io_b = io_pp_16[35]; // @[wallace.scala 70:18]
  assign FullAdder_886_io_ci = io_pp_17[34]; // @[wallace.scala 71:19]
  assign FullAdder_887_io_a = io_pp_18[33]; // @[wallace.scala 69:18]
  assign FullAdder_887_io_b = io_pp_19[32]; // @[wallace.scala 70:18]
  assign FullAdder_887_io_ci = io_pp_20[31]; // @[wallace.scala 71:19]
  assign FullAdder_888_io_a = io_pp_21[30]; // @[wallace.scala 69:18]
  assign FullAdder_888_io_b = io_pp_22[29]; // @[wallace.scala 70:18]
  assign FullAdder_888_io_ci = io_pp_23[28]; // @[wallace.scala 71:19]
  assign FullAdder_889_io_a = io_pp_24[27]; // @[wallace.scala 69:18]
  assign FullAdder_889_io_b = io_pp_25[26]; // @[wallace.scala 70:18]
  assign FullAdder_889_io_ci = io_pp_26[25]; // @[wallace.scala 71:19]
  assign FullAdder_890_io_a = io_pp_27[24]; // @[wallace.scala 69:18]
  assign FullAdder_890_io_b = io_pp_28[23]; // @[wallace.scala 70:18]
  assign FullAdder_890_io_ci = io_pp_29[22]; // @[wallace.scala 71:19]
  assign FullAdder_891_io_a = io_pp_30[21]; // @[wallace.scala 69:18]
  assign FullAdder_891_io_b = io_pp_31[20]; // @[wallace.scala 70:18]
  assign FullAdder_891_io_ci = io_pp_32[19]; // @[wallace.scala 71:19]
  assign FullAdder_892_io_a = io_pp_33[18]; // @[wallace.scala 69:18]
  assign FullAdder_892_io_b = io_pp_34[17]; // @[wallace.scala 70:18]
  assign FullAdder_892_io_ci = io_pp_35[16]; // @[wallace.scala 71:19]
  assign FullAdder_893_io_a = io_pp_36[15]; // @[wallace.scala 69:18]
  assign FullAdder_893_io_b = io_pp_37[14]; // @[wallace.scala 70:18]
  assign FullAdder_893_io_ci = io_pp_38[13]; // @[wallace.scala 71:19]
  assign FullAdder_894_io_a = io_pp_39[12]; // @[wallace.scala 69:18]
  assign FullAdder_894_io_b = io_pp_40[11]; // @[wallace.scala 70:18]
  assign FullAdder_894_io_ci = io_pp_41[10]; // @[wallace.scala 71:19]
  assign FullAdder_895_io_a = io_pp_42[9]; // @[wallace.scala 69:18]
  assign FullAdder_895_io_b = io_pp_43[8]; // @[wallace.scala 70:18]
  assign FullAdder_895_io_ci = io_pp_44[7]; // @[wallace.scala 71:19]
  assign FullAdder_896_io_a = io_pp_45[6]; // @[wallace.scala 69:18]
  assign FullAdder_896_io_b = io_pp_46[5]; // @[wallace.scala 70:18]
  assign FullAdder_896_io_ci = io_pp_47[4]; // @[wallace.scala 71:19]
  assign FullAdder_897_io_a = io_pp_48[3]; // @[wallace.scala 69:18]
  assign FullAdder_897_io_b = io_pp_49[2]; // @[wallace.scala 70:18]
  assign FullAdder_897_io_ci = io_pp_50[1]; // @[wallace.scala 71:19]
  assign FullAdder_898_io_a = io_pp_0[50]; // @[wallace.scala 69:18]
  assign FullAdder_898_io_b = io_pp_1[49]; // @[wallace.scala 70:18]
  assign FullAdder_898_io_ci = io_pp_2[48]; // @[wallace.scala 71:19]
  assign FullAdder_899_io_a = io_pp_3[47]; // @[wallace.scala 69:18]
  assign FullAdder_899_io_b = io_pp_4[46]; // @[wallace.scala 70:18]
  assign FullAdder_899_io_ci = io_pp_5[45]; // @[wallace.scala 71:19]
  assign FullAdder_900_io_a = io_pp_6[44]; // @[wallace.scala 69:18]
  assign FullAdder_900_io_b = io_pp_7[43]; // @[wallace.scala 70:18]
  assign FullAdder_900_io_ci = io_pp_8[42]; // @[wallace.scala 71:19]
  assign FullAdder_901_io_a = io_pp_9[41]; // @[wallace.scala 69:18]
  assign FullAdder_901_io_b = io_pp_10[40]; // @[wallace.scala 70:18]
  assign FullAdder_901_io_ci = io_pp_11[39]; // @[wallace.scala 71:19]
  assign FullAdder_902_io_a = io_pp_12[38]; // @[wallace.scala 69:18]
  assign FullAdder_902_io_b = io_pp_13[37]; // @[wallace.scala 70:18]
  assign FullAdder_902_io_ci = io_pp_14[36]; // @[wallace.scala 71:19]
  assign FullAdder_903_io_a = io_pp_15[35]; // @[wallace.scala 69:18]
  assign FullAdder_903_io_b = io_pp_16[34]; // @[wallace.scala 70:18]
  assign FullAdder_903_io_ci = io_pp_17[33]; // @[wallace.scala 71:19]
  assign FullAdder_904_io_a = io_pp_18[32]; // @[wallace.scala 69:18]
  assign FullAdder_904_io_b = io_pp_19[31]; // @[wallace.scala 70:18]
  assign FullAdder_904_io_ci = io_pp_20[30]; // @[wallace.scala 71:19]
  assign FullAdder_905_io_a = io_pp_21[29]; // @[wallace.scala 69:18]
  assign FullAdder_905_io_b = io_pp_22[28]; // @[wallace.scala 70:18]
  assign FullAdder_905_io_ci = io_pp_23[27]; // @[wallace.scala 71:19]
  assign FullAdder_906_io_a = io_pp_24[26]; // @[wallace.scala 69:18]
  assign FullAdder_906_io_b = io_pp_25[25]; // @[wallace.scala 70:18]
  assign FullAdder_906_io_ci = io_pp_26[24]; // @[wallace.scala 71:19]
  assign FullAdder_907_io_a = io_pp_27[23]; // @[wallace.scala 69:18]
  assign FullAdder_907_io_b = io_pp_28[22]; // @[wallace.scala 70:18]
  assign FullAdder_907_io_ci = io_pp_29[21]; // @[wallace.scala 71:19]
  assign FullAdder_908_io_a = io_pp_30[20]; // @[wallace.scala 69:18]
  assign FullAdder_908_io_b = io_pp_31[19]; // @[wallace.scala 70:18]
  assign FullAdder_908_io_ci = io_pp_32[18]; // @[wallace.scala 71:19]
  assign FullAdder_909_io_a = io_pp_33[17]; // @[wallace.scala 69:18]
  assign FullAdder_909_io_b = io_pp_34[16]; // @[wallace.scala 70:18]
  assign FullAdder_909_io_ci = io_pp_35[15]; // @[wallace.scala 71:19]
  assign FullAdder_910_io_a = io_pp_36[14]; // @[wallace.scala 69:18]
  assign FullAdder_910_io_b = io_pp_37[13]; // @[wallace.scala 70:18]
  assign FullAdder_910_io_ci = io_pp_38[12]; // @[wallace.scala 71:19]
  assign FullAdder_911_io_a = io_pp_39[11]; // @[wallace.scala 69:18]
  assign FullAdder_911_io_b = io_pp_40[10]; // @[wallace.scala 70:18]
  assign FullAdder_911_io_ci = io_pp_41[9]; // @[wallace.scala 71:19]
  assign FullAdder_912_io_a = io_pp_42[8]; // @[wallace.scala 69:18]
  assign FullAdder_912_io_b = io_pp_43[7]; // @[wallace.scala 70:18]
  assign FullAdder_912_io_ci = io_pp_44[6]; // @[wallace.scala 71:19]
  assign FullAdder_913_io_a = io_pp_45[5]; // @[wallace.scala 69:18]
  assign FullAdder_913_io_b = io_pp_46[4]; // @[wallace.scala 70:18]
  assign FullAdder_913_io_ci = io_pp_47[3]; // @[wallace.scala 71:19]
  assign FullAdder_914_io_a = io_pp_48[2]; // @[wallace.scala 69:18]
  assign FullAdder_914_io_b = io_pp_49[1]; // @[wallace.scala 70:18]
  assign FullAdder_914_io_ci = io_pp_50[0]; // @[wallace.scala 71:19]
  assign FullAdder_915_io_a = io_pp_0[49]; // @[wallace.scala 69:18]
  assign FullAdder_915_io_b = io_pp_1[48]; // @[wallace.scala 70:18]
  assign FullAdder_915_io_ci = io_pp_2[47]; // @[wallace.scala 71:19]
  assign FullAdder_916_io_a = io_pp_3[46]; // @[wallace.scala 69:18]
  assign FullAdder_916_io_b = io_pp_4[45]; // @[wallace.scala 70:18]
  assign FullAdder_916_io_ci = io_pp_5[44]; // @[wallace.scala 71:19]
  assign FullAdder_917_io_a = io_pp_6[43]; // @[wallace.scala 69:18]
  assign FullAdder_917_io_b = io_pp_7[42]; // @[wallace.scala 70:18]
  assign FullAdder_917_io_ci = io_pp_8[41]; // @[wallace.scala 71:19]
  assign FullAdder_918_io_a = io_pp_9[40]; // @[wallace.scala 69:18]
  assign FullAdder_918_io_b = io_pp_10[39]; // @[wallace.scala 70:18]
  assign FullAdder_918_io_ci = io_pp_11[38]; // @[wallace.scala 71:19]
  assign FullAdder_919_io_a = io_pp_12[37]; // @[wallace.scala 69:18]
  assign FullAdder_919_io_b = io_pp_13[36]; // @[wallace.scala 70:18]
  assign FullAdder_919_io_ci = io_pp_14[35]; // @[wallace.scala 71:19]
  assign FullAdder_920_io_a = io_pp_15[34]; // @[wallace.scala 69:18]
  assign FullAdder_920_io_b = io_pp_16[33]; // @[wallace.scala 70:18]
  assign FullAdder_920_io_ci = io_pp_17[32]; // @[wallace.scala 71:19]
  assign FullAdder_921_io_a = io_pp_18[31]; // @[wallace.scala 69:18]
  assign FullAdder_921_io_b = io_pp_19[30]; // @[wallace.scala 70:18]
  assign FullAdder_921_io_ci = io_pp_20[29]; // @[wallace.scala 71:19]
  assign FullAdder_922_io_a = io_pp_21[28]; // @[wallace.scala 69:18]
  assign FullAdder_922_io_b = io_pp_22[27]; // @[wallace.scala 70:18]
  assign FullAdder_922_io_ci = io_pp_23[26]; // @[wallace.scala 71:19]
  assign FullAdder_923_io_a = io_pp_24[25]; // @[wallace.scala 69:18]
  assign FullAdder_923_io_b = io_pp_25[24]; // @[wallace.scala 70:18]
  assign FullAdder_923_io_ci = io_pp_26[23]; // @[wallace.scala 71:19]
  assign FullAdder_924_io_a = io_pp_27[22]; // @[wallace.scala 69:18]
  assign FullAdder_924_io_b = io_pp_28[21]; // @[wallace.scala 70:18]
  assign FullAdder_924_io_ci = io_pp_29[20]; // @[wallace.scala 71:19]
  assign FullAdder_925_io_a = io_pp_30[19]; // @[wallace.scala 69:18]
  assign FullAdder_925_io_b = io_pp_31[18]; // @[wallace.scala 70:18]
  assign FullAdder_925_io_ci = io_pp_32[17]; // @[wallace.scala 71:19]
  assign FullAdder_926_io_a = io_pp_33[16]; // @[wallace.scala 69:18]
  assign FullAdder_926_io_b = io_pp_34[15]; // @[wallace.scala 70:18]
  assign FullAdder_926_io_ci = io_pp_35[14]; // @[wallace.scala 71:19]
  assign FullAdder_927_io_a = io_pp_36[13]; // @[wallace.scala 69:18]
  assign FullAdder_927_io_b = io_pp_37[12]; // @[wallace.scala 70:18]
  assign FullAdder_927_io_ci = io_pp_38[11]; // @[wallace.scala 71:19]
  assign FullAdder_928_io_a = io_pp_39[10]; // @[wallace.scala 69:18]
  assign FullAdder_928_io_b = io_pp_40[9]; // @[wallace.scala 70:18]
  assign FullAdder_928_io_ci = io_pp_41[8]; // @[wallace.scala 71:19]
  assign FullAdder_929_io_a = io_pp_42[7]; // @[wallace.scala 69:18]
  assign FullAdder_929_io_b = io_pp_43[6]; // @[wallace.scala 70:18]
  assign FullAdder_929_io_ci = io_pp_44[5]; // @[wallace.scala 71:19]
  assign FullAdder_930_io_a = io_pp_45[4]; // @[wallace.scala 69:18]
  assign FullAdder_930_io_b = io_pp_46[3]; // @[wallace.scala 70:18]
  assign FullAdder_930_io_ci = io_pp_47[2]; // @[wallace.scala 71:19]
  assign FullAdder_931_io_a = io_pp_0[48]; // @[wallace.scala 69:18]
  assign FullAdder_931_io_b = io_pp_1[47]; // @[wallace.scala 70:18]
  assign FullAdder_931_io_ci = io_pp_2[46]; // @[wallace.scala 71:19]
  assign FullAdder_932_io_a = io_pp_3[45]; // @[wallace.scala 69:18]
  assign FullAdder_932_io_b = io_pp_4[44]; // @[wallace.scala 70:18]
  assign FullAdder_932_io_ci = io_pp_5[43]; // @[wallace.scala 71:19]
  assign FullAdder_933_io_a = io_pp_6[42]; // @[wallace.scala 69:18]
  assign FullAdder_933_io_b = io_pp_7[41]; // @[wallace.scala 70:18]
  assign FullAdder_933_io_ci = io_pp_8[40]; // @[wallace.scala 71:19]
  assign FullAdder_934_io_a = io_pp_9[39]; // @[wallace.scala 69:18]
  assign FullAdder_934_io_b = io_pp_10[38]; // @[wallace.scala 70:18]
  assign FullAdder_934_io_ci = io_pp_11[37]; // @[wallace.scala 71:19]
  assign FullAdder_935_io_a = io_pp_12[36]; // @[wallace.scala 69:18]
  assign FullAdder_935_io_b = io_pp_13[35]; // @[wallace.scala 70:18]
  assign FullAdder_935_io_ci = io_pp_14[34]; // @[wallace.scala 71:19]
  assign FullAdder_936_io_a = io_pp_15[33]; // @[wallace.scala 69:18]
  assign FullAdder_936_io_b = io_pp_16[32]; // @[wallace.scala 70:18]
  assign FullAdder_936_io_ci = io_pp_17[31]; // @[wallace.scala 71:19]
  assign FullAdder_937_io_a = io_pp_18[30]; // @[wallace.scala 69:18]
  assign FullAdder_937_io_b = io_pp_19[29]; // @[wallace.scala 70:18]
  assign FullAdder_937_io_ci = io_pp_20[28]; // @[wallace.scala 71:19]
  assign FullAdder_938_io_a = io_pp_21[27]; // @[wallace.scala 69:18]
  assign FullAdder_938_io_b = io_pp_22[26]; // @[wallace.scala 70:18]
  assign FullAdder_938_io_ci = io_pp_23[25]; // @[wallace.scala 71:19]
  assign FullAdder_939_io_a = io_pp_24[24]; // @[wallace.scala 69:18]
  assign FullAdder_939_io_b = io_pp_25[23]; // @[wallace.scala 70:18]
  assign FullAdder_939_io_ci = io_pp_26[22]; // @[wallace.scala 71:19]
  assign FullAdder_940_io_a = io_pp_27[21]; // @[wallace.scala 69:18]
  assign FullAdder_940_io_b = io_pp_28[20]; // @[wallace.scala 70:18]
  assign FullAdder_940_io_ci = io_pp_29[19]; // @[wallace.scala 71:19]
  assign FullAdder_941_io_a = io_pp_30[18]; // @[wallace.scala 69:18]
  assign FullAdder_941_io_b = io_pp_31[17]; // @[wallace.scala 70:18]
  assign FullAdder_941_io_ci = io_pp_32[16]; // @[wallace.scala 71:19]
  assign FullAdder_942_io_a = io_pp_33[15]; // @[wallace.scala 69:18]
  assign FullAdder_942_io_b = io_pp_34[14]; // @[wallace.scala 70:18]
  assign FullAdder_942_io_ci = io_pp_35[13]; // @[wallace.scala 71:19]
  assign FullAdder_943_io_a = io_pp_36[12]; // @[wallace.scala 69:18]
  assign FullAdder_943_io_b = io_pp_37[11]; // @[wallace.scala 70:18]
  assign FullAdder_943_io_ci = io_pp_38[10]; // @[wallace.scala 71:19]
  assign FullAdder_944_io_a = io_pp_39[9]; // @[wallace.scala 69:18]
  assign FullAdder_944_io_b = io_pp_40[8]; // @[wallace.scala 70:18]
  assign FullAdder_944_io_ci = io_pp_41[7]; // @[wallace.scala 71:19]
  assign FullAdder_945_io_a = io_pp_42[6]; // @[wallace.scala 69:18]
  assign FullAdder_945_io_b = io_pp_43[5]; // @[wallace.scala 70:18]
  assign FullAdder_945_io_ci = io_pp_44[4]; // @[wallace.scala 71:19]
  assign FullAdder_946_io_a = io_pp_45[3]; // @[wallace.scala 69:18]
  assign FullAdder_946_io_b = io_pp_46[2]; // @[wallace.scala 70:18]
  assign FullAdder_946_io_ci = io_pp_47[1]; // @[wallace.scala 71:19]
  assign FullAdder_947_io_a = io_pp_0[47]; // @[wallace.scala 69:18]
  assign FullAdder_947_io_b = io_pp_1[46]; // @[wallace.scala 70:18]
  assign FullAdder_947_io_ci = io_pp_2[45]; // @[wallace.scala 71:19]
  assign FullAdder_948_io_a = io_pp_3[44]; // @[wallace.scala 69:18]
  assign FullAdder_948_io_b = io_pp_4[43]; // @[wallace.scala 70:18]
  assign FullAdder_948_io_ci = io_pp_5[42]; // @[wallace.scala 71:19]
  assign FullAdder_949_io_a = io_pp_6[41]; // @[wallace.scala 69:18]
  assign FullAdder_949_io_b = io_pp_7[40]; // @[wallace.scala 70:18]
  assign FullAdder_949_io_ci = io_pp_8[39]; // @[wallace.scala 71:19]
  assign FullAdder_950_io_a = io_pp_9[38]; // @[wallace.scala 69:18]
  assign FullAdder_950_io_b = io_pp_10[37]; // @[wallace.scala 70:18]
  assign FullAdder_950_io_ci = io_pp_11[36]; // @[wallace.scala 71:19]
  assign FullAdder_951_io_a = io_pp_12[35]; // @[wallace.scala 69:18]
  assign FullAdder_951_io_b = io_pp_13[34]; // @[wallace.scala 70:18]
  assign FullAdder_951_io_ci = io_pp_14[33]; // @[wallace.scala 71:19]
  assign FullAdder_952_io_a = io_pp_15[32]; // @[wallace.scala 69:18]
  assign FullAdder_952_io_b = io_pp_16[31]; // @[wallace.scala 70:18]
  assign FullAdder_952_io_ci = io_pp_17[30]; // @[wallace.scala 71:19]
  assign FullAdder_953_io_a = io_pp_18[29]; // @[wallace.scala 69:18]
  assign FullAdder_953_io_b = io_pp_19[28]; // @[wallace.scala 70:18]
  assign FullAdder_953_io_ci = io_pp_20[27]; // @[wallace.scala 71:19]
  assign FullAdder_954_io_a = io_pp_21[26]; // @[wallace.scala 69:18]
  assign FullAdder_954_io_b = io_pp_22[25]; // @[wallace.scala 70:18]
  assign FullAdder_954_io_ci = io_pp_23[24]; // @[wallace.scala 71:19]
  assign FullAdder_955_io_a = io_pp_24[23]; // @[wallace.scala 69:18]
  assign FullAdder_955_io_b = io_pp_25[22]; // @[wallace.scala 70:18]
  assign FullAdder_955_io_ci = io_pp_26[21]; // @[wallace.scala 71:19]
  assign FullAdder_956_io_a = io_pp_27[20]; // @[wallace.scala 69:18]
  assign FullAdder_956_io_b = io_pp_28[19]; // @[wallace.scala 70:18]
  assign FullAdder_956_io_ci = io_pp_29[18]; // @[wallace.scala 71:19]
  assign FullAdder_957_io_a = io_pp_30[17]; // @[wallace.scala 69:18]
  assign FullAdder_957_io_b = io_pp_31[16]; // @[wallace.scala 70:18]
  assign FullAdder_957_io_ci = io_pp_32[15]; // @[wallace.scala 71:19]
  assign FullAdder_958_io_a = io_pp_33[14]; // @[wallace.scala 69:18]
  assign FullAdder_958_io_b = io_pp_34[13]; // @[wallace.scala 70:18]
  assign FullAdder_958_io_ci = io_pp_35[12]; // @[wallace.scala 71:19]
  assign FullAdder_959_io_a = io_pp_36[11]; // @[wallace.scala 69:18]
  assign FullAdder_959_io_b = io_pp_37[10]; // @[wallace.scala 70:18]
  assign FullAdder_959_io_ci = io_pp_38[9]; // @[wallace.scala 71:19]
  assign FullAdder_960_io_a = io_pp_39[8]; // @[wallace.scala 69:18]
  assign FullAdder_960_io_b = io_pp_40[7]; // @[wallace.scala 70:18]
  assign FullAdder_960_io_ci = io_pp_41[6]; // @[wallace.scala 71:19]
  assign FullAdder_961_io_a = io_pp_42[5]; // @[wallace.scala 69:18]
  assign FullAdder_961_io_b = io_pp_43[4]; // @[wallace.scala 70:18]
  assign FullAdder_961_io_ci = io_pp_44[3]; // @[wallace.scala 71:19]
  assign FullAdder_962_io_a = io_pp_45[2]; // @[wallace.scala 69:18]
  assign FullAdder_962_io_b = io_pp_46[1]; // @[wallace.scala 70:18]
  assign FullAdder_962_io_ci = io_pp_47[0]; // @[wallace.scala 71:19]
  assign FullAdder_963_io_a = io_pp_0[46]; // @[wallace.scala 69:18]
  assign FullAdder_963_io_b = io_pp_1[45]; // @[wallace.scala 70:18]
  assign FullAdder_963_io_ci = io_pp_2[44]; // @[wallace.scala 71:19]
  assign FullAdder_964_io_a = io_pp_3[43]; // @[wallace.scala 69:18]
  assign FullAdder_964_io_b = io_pp_4[42]; // @[wallace.scala 70:18]
  assign FullAdder_964_io_ci = io_pp_5[41]; // @[wallace.scala 71:19]
  assign FullAdder_965_io_a = io_pp_6[40]; // @[wallace.scala 69:18]
  assign FullAdder_965_io_b = io_pp_7[39]; // @[wallace.scala 70:18]
  assign FullAdder_965_io_ci = io_pp_8[38]; // @[wallace.scala 71:19]
  assign FullAdder_966_io_a = io_pp_9[37]; // @[wallace.scala 69:18]
  assign FullAdder_966_io_b = io_pp_10[36]; // @[wallace.scala 70:18]
  assign FullAdder_966_io_ci = io_pp_11[35]; // @[wallace.scala 71:19]
  assign FullAdder_967_io_a = io_pp_12[34]; // @[wallace.scala 69:18]
  assign FullAdder_967_io_b = io_pp_13[33]; // @[wallace.scala 70:18]
  assign FullAdder_967_io_ci = io_pp_14[32]; // @[wallace.scala 71:19]
  assign FullAdder_968_io_a = io_pp_15[31]; // @[wallace.scala 69:18]
  assign FullAdder_968_io_b = io_pp_16[30]; // @[wallace.scala 70:18]
  assign FullAdder_968_io_ci = io_pp_17[29]; // @[wallace.scala 71:19]
  assign FullAdder_969_io_a = io_pp_18[28]; // @[wallace.scala 69:18]
  assign FullAdder_969_io_b = io_pp_19[27]; // @[wallace.scala 70:18]
  assign FullAdder_969_io_ci = io_pp_20[26]; // @[wallace.scala 71:19]
  assign FullAdder_970_io_a = io_pp_21[25]; // @[wallace.scala 69:18]
  assign FullAdder_970_io_b = io_pp_22[24]; // @[wallace.scala 70:18]
  assign FullAdder_970_io_ci = io_pp_23[23]; // @[wallace.scala 71:19]
  assign FullAdder_971_io_a = io_pp_24[22]; // @[wallace.scala 69:18]
  assign FullAdder_971_io_b = io_pp_25[21]; // @[wallace.scala 70:18]
  assign FullAdder_971_io_ci = io_pp_26[20]; // @[wallace.scala 71:19]
  assign FullAdder_972_io_a = io_pp_27[19]; // @[wallace.scala 69:18]
  assign FullAdder_972_io_b = io_pp_28[18]; // @[wallace.scala 70:18]
  assign FullAdder_972_io_ci = io_pp_29[17]; // @[wallace.scala 71:19]
  assign FullAdder_973_io_a = io_pp_30[16]; // @[wallace.scala 69:18]
  assign FullAdder_973_io_b = io_pp_31[15]; // @[wallace.scala 70:18]
  assign FullAdder_973_io_ci = io_pp_32[14]; // @[wallace.scala 71:19]
  assign FullAdder_974_io_a = io_pp_33[13]; // @[wallace.scala 69:18]
  assign FullAdder_974_io_b = io_pp_34[12]; // @[wallace.scala 70:18]
  assign FullAdder_974_io_ci = io_pp_35[11]; // @[wallace.scala 71:19]
  assign FullAdder_975_io_a = io_pp_36[10]; // @[wallace.scala 69:18]
  assign FullAdder_975_io_b = io_pp_37[9]; // @[wallace.scala 70:18]
  assign FullAdder_975_io_ci = io_pp_38[8]; // @[wallace.scala 71:19]
  assign FullAdder_976_io_a = io_pp_39[7]; // @[wallace.scala 69:18]
  assign FullAdder_976_io_b = io_pp_40[6]; // @[wallace.scala 70:18]
  assign FullAdder_976_io_ci = io_pp_41[5]; // @[wallace.scala 71:19]
  assign FullAdder_977_io_a = io_pp_42[4]; // @[wallace.scala 69:18]
  assign FullAdder_977_io_b = io_pp_43[3]; // @[wallace.scala 70:18]
  assign FullAdder_977_io_ci = io_pp_44[2]; // @[wallace.scala 71:19]
  assign HalfAdder_21_io_a = io_pp_45[1]; // @[wallace.scala 59:18]
  assign HalfAdder_21_io_b = io_pp_46[0]; // @[wallace.scala 60:18]
  assign FullAdder_978_io_a = io_pp_0[45]; // @[wallace.scala 69:18]
  assign FullAdder_978_io_b = io_pp_1[44]; // @[wallace.scala 70:18]
  assign FullAdder_978_io_ci = io_pp_2[43]; // @[wallace.scala 71:19]
  assign FullAdder_979_io_a = io_pp_3[42]; // @[wallace.scala 69:18]
  assign FullAdder_979_io_b = io_pp_4[41]; // @[wallace.scala 70:18]
  assign FullAdder_979_io_ci = io_pp_5[40]; // @[wallace.scala 71:19]
  assign FullAdder_980_io_a = io_pp_6[39]; // @[wallace.scala 69:18]
  assign FullAdder_980_io_b = io_pp_7[38]; // @[wallace.scala 70:18]
  assign FullAdder_980_io_ci = io_pp_8[37]; // @[wallace.scala 71:19]
  assign FullAdder_981_io_a = io_pp_9[36]; // @[wallace.scala 69:18]
  assign FullAdder_981_io_b = io_pp_10[35]; // @[wallace.scala 70:18]
  assign FullAdder_981_io_ci = io_pp_11[34]; // @[wallace.scala 71:19]
  assign FullAdder_982_io_a = io_pp_12[33]; // @[wallace.scala 69:18]
  assign FullAdder_982_io_b = io_pp_13[32]; // @[wallace.scala 70:18]
  assign FullAdder_982_io_ci = io_pp_14[31]; // @[wallace.scala 71:19]
  assign FullAdder_983_io_a = io_pp_15[30]; // @[wallace.scala 69:18]
  assign FullAdder_983_io_b = io_pp_16[29]; // @[wallace.scala 70:18]
  assign FullAdder_983_io_ci = io_pp_17[28]; // @[wallace.scala 71:19]
  assign FullAdder_984_io_a = io_pp_18[27]; // @[wallace.scala 69:18]
  assign FullAdder_984_io_b = io_pp_19[26]; // @[wallace.scala 70:18]
  assign FullAdder_984_io_ci = io_pp_20[25]; // @[wallace.scala 71:19]
  assign FullAdder_985_io_a = io_pp_21[24]; // @[wallace.scala 69:18]
  assign FullAdder_985_io_b = io_pp_22[23]; // @[wallace.scala 70:18]
  assign FullAdder_985_io_ci = io_pp_23[22]; // @[wallace.scala 71:19]
  assign FullAdder_986_io_a = io_pp_24[21]; // @[wallace.scala 69:18]
  assign FullAdder_986_io_b = io_pp_25[20]; // @[wallace.scala 70:18]
  assign FullAdder_986_io_ci = io_pp_26[19]; // @[wallace.scala 71:19]
  assign FullAdder_987_io_a = io_pp_27[18]; // @[wallace.scala 69:18]
  assign FullAdder_987_io_b = io_pp_28[17]; // @[wallace.scala 70:18]
  assign FullAdder_987_io_ci = io_pp_29[16]; // @[wallace.scala 71:19]
  assign FullAdder_988_io_a = io_pp_30[15]; // @[wallace.scala 69:18]
  assign FullAdder_988_io_b = io_pp_31[14]; // @[wallace.scala 70:18]
  assign FullAdder_988_io_ci = io_pp_32[13]; // @[wallace.scala 71:19]
  assign FullAdder_989_io_a = io_pp_33[12]; // @[wallace.scala 69:18]
  assign FullAdder_989_io_b = io_pp_34[11]; // @[wallace.scala 70:18]
  assign FullAdder_989_io_ci = io_pp_35[10]; // @[wallace.scala 71:19]
  assign FullAdder_990_io_a = io_pp_36[9]; // @[wallace.scala 69:18]
  assign FullAdder_990_io_b = io_pp_37[8]; // @[wallace.scala 70:18]
  assign FullAdder_990_io_ci = io_pp_38[7]; // @[wallace.scala 71:19]
  assign FullAdder_991_io_a = io_pp_39[6]; // @[wallace.scala 69:18]
  assign FullAdder_991_io_b = io_pp_40[5]; // @[wallace.scala 70:18]
  assign FullAdder_991_io_ci = io_pp_41[4]; // @[wallace.scala 71:19]
  assign FullAdder_992_io_a = io_pp_42[3]; // @[wallace.scala 69:18]
  assign FullAdder_992_io_b = io_pp_43[2]; // @[wallace.scala 70:18]
  assign FullAdder_992_io_ci = io_pp_44[1]; // @[wallace.scala 71:19]
  assign FullAdder_993_io_a = io_pp_0[44]; // @[wallace.scala 69:18]
  assign FullAdder_993_io_b = io_pp_1[43]; // @[wallace.scala 70:18]
  assign FullAdder_993_io_ci = io_pp_2[42]; // @[wallace.scala 71:19]
  assign FullAdder_994_io_a = io_pp_3[41]; // @[wallace.scala 69:18]
  assign FullAdder_994_io_b = io_pp_4[40]; // @[wallace.scala 70:18]
  assign FullAdder_994_io_ci = io_pp_5[39]; // @[wallace.scala 71:19]
  assign FullAdder_995_io_a = io_pp_6[38]; // @[wallace.scala 69:18]
  assign FullAdder_995_io_b = io_pp_7[37]; // @[wallace.scala 70:18]
  assign FullAdder_995_io_ci = io_pp_8[36]; // @[wallace.scala 71:19]
  assign FullAdder_996_io_a = io_pp_9[35]; // @[wallace.scala 69:18]
  assign FullAdder_996_io_b = io_pp_10[34]; // @[wallace.scala 70:18]
  assign FullAdder_996_io_ci = io_pp_11[33]; // @[wallace.scala 71:19]
  assign FullAdder_997_io_a = io_pp_12[32]; // @[wallace.scala 69:18]
  assign FullAdder_997_io_b = io_pp_13[31]; // @[wallace.scala 70:18]
  assign FullAdder_997_io_ci = io_pp_14[30]; // @[wallace.scala 71:19]
  assign FullAdder_998_io_a = io_pp_15[29]; // @[wallace.scala 69:18]
  assign FullAdder_998_io_b = io_pp_16[28]; // @[wallace.scala 70:18]
  assign FullAdder_998_io_ci = io_pp_17[27]; // @[wallace.scala 71:19]
  assign FullAdder_999_io_a = io_pp_18[26]; // @[wallace.scala 69:18]
  assign FullAdder_999_io_b = io_pp_19[25]; // @[wallace.scala 70:18]
  assign FullAdder_999_io_ci = io_pp_20[24]; // @[wallace.scala 71:19]
  assign FullAdder_1000_io_a = io_pp_21[23]; // @[wallace.scala 69:18]
  assign FullAdder_1000_io_b = io_pp_22[22]; // @[wallace.scala 70:18]
  assign FullAdder_1000_io_ci = io_pp_23[21]; // @[wallace.scala 71:19]
  assign FullAdder_1001_io_a = io_pp_24[20]; // @[wallace.scala 69:18]
  assign FullAdder_1001_io_b = io_pp_25[19]; // @[wallace.scala 70:18]
  assign FullAdder_1001_io_ci = io_pp_26[18]; // @[wallace.scala 71:19]
  assign FullAdder_1002_io_a = io_pp_27[17]; // @[wallace.scala 69:18]
  assign FullAdder_1002_io_b = io_pp_28[16]; // @[wallace.scala 70:18]
  assign FullAdder_1002_io_ci = io_pp_29[15]; // @[wallace.scala 71:19]
  assign FullAdder_1003_io_a = io_pp_30[14]; // @[wallace.scala 69:18]
  assign FullAdder_1003_io_b = io_pp_31[13]; // @[wallace.scala 70:18]
  assign FullAdder_1003_io_ci = io_pp_32[12]; // @[wallace.scala 71:19]
  assign FullAdder_1004_io_a = io_pp_33[11]; // @[wallace.scala 69:18]
  assign FullAdder_1004_io_b = io_pp_34[10]; // @[wallace.scala 70:18]
  assign FullAdder_1004_io_ci = io_pp_35[9]; // @[wallace.scala 71:19]
  assign FullAdder_1005_io_a = io_pp_36[8]; // @[wallace.scala 69:18]
  assign FullAdder_1005_io_b = io_pp_37[7]; // @[wallace.scala 70:18]
  assign FullAdder_1005_io_ci = io_pp_38[6]; // @[wallace.scala 71:19]
  assign FullAdder_1006_io_a = io_pp_39[5]; // @[wallace.scala 69:18]
  assign FullAdder_1006_io_b = io_pp_40[4]; // @[wallace.scala 70:18]
  assign FullAdder_1006_io_ci = io_pp_41[3]; // @[wallace.scala 71:19]
  assign FullAdder_1007_io_a = io_pp_42[2]; // @[wallace.scala 69:18]
  assign FullAdder_1007_io_b = io_pp_43[1]; // @[wallace.scala 70:18]
  assign FullAdder_1007_io_ci = io_pp_44[0]; // @[wallace.scala 71:19]
  assign FullAdder_1008_io_a = io_pp_0[43]; // @[wallace.scala 69:18]
  assign FullAdder_1008_io_b = io_pp_1[42]; // @[wallace.scala 70:18]
  assign FullAdder_1008_io_ci = io_pp_2[41]; // @[wallace.scala 71:19]
  assign FullAdder_1009_io_a = io_pp_3[40]; // @[wallace.scala 69:18]
  assign FullAdder_1009_io_b = io_pp_4[39]; // @[wallace.scala 70:18]
  assign FullAdder_1009_io_ci = io_pp_5[38]; // @[wallace.scala 71:19]
  assign FullAdder_1010_io_a = io_pp_6[37]; // @[wallace.scala 69:18]
  assign FullAdder_1010_io_b = io_pp_7[36]; // @[wallace.scala 70:18]
  assign FullAdder_1010_io_ci = io_pp_8[35]; // @[wallace.scala 71:19]
  assign FullAdder_1011_io_a = io_pp_9[34]; // @[wallace.scala 69:18]
  assign FullAdder_1011_io_b = io_pp_10[33]; // @[wallace.scala 70:18]
  assign FullAdder_1011_io_ci = io_pp_11[32]; // @[wallace.scala 71:19]
  assign FullAdder_1012_io_a = io_pp_12[31]; // @[wallace.scala 69:18]
  assign FullAdder_1012_io_b = io_pp_13[30]; // @[wallace.scala 70:18]
  assign FullAdder_1012_io_ci = io_pp_14[29]; // @[wallace.scala 71:19]
  assign FullAdder_1013_io_a = io_pp_15[28]; // @[wallace.scala 69:18]
  assign FullAdder_1013_io_b = io_pp_16[27]; // @[wallace.scala 70:18]
  assign FullAdder_1013_io_ci = io_pp_17[26]; // @[wallace.scala 71:19]
  assign FullAdder_1014_io_a = io_pp_18[25]; // @[wallace.scala 69:18]
  assign FullAdder_1014_io_b = io_pp_19[24]; // @[wallace.scala 70:18]
  assign FullAdder_1014_io_ci = io_pp_20[23]; // @[wallace.scala 71:19]
  assign FullAdder_1015_io_a = io_pp_21[22]; // @[wallace.scala 69:18]
  assign FullAdder_1015_io_b = io_pp_22[21]; // @[wallace.scala 70:18]
  assign FullAdder_1015_io_ci = io_pp_23[20]; // @[wallace.scala 71:19]
  assign FullAdder_1016_io_a = io_pp_24[19]; // @[wallace.scala 69:18]
  assign FullAdder_1016_io_b = io_pp_25[18]; // @[wallace.scala 70:18]
  assign FullAdder_1016_io_ci = io_pp_26[17]; // @[wallace.scala 71:19]
  assign FullAdder_1017_io_a = io_pp_27[16]; // @[wallace.scala 69:18]
  assign FullAdder_1017_io_b = io_pp_28[15]; // @[wallace.scala 70:18]
  assign FullAdder_1017_io_ci = io_pp_29[14]; // @[wallace.scala 71:19]
  assign FullAdder_1018_io_a = io_pp_30[13]; // @[wallace.scala 69:18]
  assign FullAdder_1018_io_b = io_pp_31[12]; // @[wallace.scala 70:18]
  assign FullAdder_1018_io_ci = io_pp_32[11]; // @[wallace.scala 71:19]
  assign FullAdder_1019_io_a = io_pp_33[10]; // @[wallace.scala 69:18]
  assign FullAdder_1019_io_b = io_pp_34[9]; // @[wallace.scala 70:18]
  assign FullAdder_1019_io_ci = io_pp_35[8]; // @[wallace.scala 71:19]
  assign FullAdder_1020_io_a = io_pp_36[7]; // @[wallace.scala 69:18]
  assign FullAdder_1020_io_b = io_pp_37[6]; // @[wallace.scala 70:18]
  assign FullAdder_1020_io_ci = io_pp_38[5]; // @[wallace.scala 71:19]
  assign FullAdder_1021_io_a = io_pp_39[4]; // @[wallace.scala 69:18]
  assign FullAdder_1021_io_b = io_pp_40[3]; // @[wallace.scala 70:18]
  assign FullAdder_1021_io_ci = io_pp_41[2]; // @[wallace.scala 71:19]
  assign FullAdder_1022_io_a = io_pp_0[42]; // @[wallace.scala 69:18]
  assign FullAdder_1022_io_b = io_pp_1[41]; // @[wallace.scala 70:18]
  assign FullAdder_1022_io_ci = io_pp_2[40]; // @[wallace.scala 71:19]
  assign FullAdder_1023_io_a = io_pp_3[39]; // @[wallace.scala 69:18]
  assign FullAdder_1023_io_b = io_pp_4[38]; // @[wallace.scala 70:18]
  assign FullAdder_1023_io_ci = io_pp_5[37]; // @[wallace.scala 71:19]
  assign FullAdder_1024_io_a = io_pp_6[36]; // @[wallace.scala 69:18]
  assign FullAdder_1024_io_b = io_pp_7[35]; // @[wallace.scala 70:18]
  assign FullAdder_1024_io_ci = io_pp_8[34]; // @[wallace.scala 71:19]
  assign FullAdder_1025_io_a = io_pp_9[33]; // @[wallace.scala 69:18]
  assign FullAdder_1025_io_b = io_pp_10[32]; // @[wallace.scala 70:18]
  assign FullAdder_1025_io_ci = io_pp_11[31]; // @[wallace.scala 71:19]
  assign FullAdder_1026_io_a = io_pp_12[30]; // @[wallace.scala 69:18]
  assign FullAdder_1026_io_b = io_pp_13[29]; // @[wallace.scala 70:18]
  assign FullAdder_1026_io_ci = io_pp_14[28]; // @[wallace.scala 71:19]
  assign FullAdder_1027_io_a = io_pp_15[27]; // @[wallace.scala 69:18]
  assign FullAdder_1027_io_b = io_pp_16[26]; // @[wallace.scala 70:18]
  assign FullAdder_1027_io_ci = io_pp_17[25]; // @[wallace.scala 71:19]
  assign FullAdder_1028_io_a = io_pp_18[24]; // @[wallace.scala 69:18]
  assign FullAdder_1028_io_b = io_pp_19[23]; // @[wallace.scala 70:18]
  assign FullAdder_1028_io_ci = io_pp_20[22]; // @[wallace.scala 71:19]
  assign FullAdder_1029_io_a = io_pp_21[21]; // @[wallace.scala 69:18]
  assign FullAdder_1029_io_b = io_pp_22[20]; // @[wallace.scala 70:18]
  assign FullAdder_1029_io_ci = io_pp_23[19]; // @[wallace.scala 71:19]
  assign FullAdder_1030_io_a = io_pp_24[18]; // @[wallace.scala 69:18]
  assign FullAdder_1030_io_b = io_pp_25[17]; // @[wallace.scala 70:18]
  assign FullAdder_1030_io_ci = io_pp_26[16]; // @[wallace.scala 71:19]
  assign FullAdder_1031_io_a = io_pp_27[15]; // @[wallace.scala 69:18]
  assign FullAdder_1031_io_b = io_pp_28[14]; // @[wallace.scala 70:18]
  assign FullAdder_1031_io_ci = io_pp_29[13]; // @[wallace.scala 71:19]
  assign FullAdder_1032_io_a = io_pp_30[12]; // @[wallace.scala 69:18]
  assign FullAdder_1032_io_b = io_pp_31[11]; // @[wallace.scala 70:18]
  assign FullAdder_1032_io_ci = io_pp_32[10]; // @[wallace.scala 71:19]
  assign FullAdder_1033_io_a = io_pp_33[9]; // @[wallace.scala 69:18]
  assign FullAdder_1033_io_b = io_pp_34[8]; // @[wallace.scala 70:18]
  assign FullAdder_1033_io_ci = io_pp_35[7]; // @[wallace.scala 71:19]
  assign FullAdder_1034_io_a = io_pp_36[6]; // @[wallace.scala 69:18]
  assign FullAdder_1034_io_b = io_pp_37[5]; // @[wallace.scala 70:18]
  assign FullAdder_1034_io_ci = io_pp_38[4]; // @[wallace.scala 71:19]
  assign FullAdder_1035_io_a = io_pp_39[3]; // @[wallace.scala 69:18]
  assign FullAdder_1035_io_b = io_pp_40[2]; // @[wallace.scala 70:18]
  assign FullAdder_1035_io_ci = io_pp_41[1]; // @[wallace.scala 71:19]
  assign FullAdder_1036_io_a = io_pp_0[41]; // @[wallace.scala 69:18]
  assign FullAdder_1036_io_b = io_pp_1[40]; // @[wallace.scala 70:18]
  assign FullAdder_1036_io_ci = io_pp_2[39]; // @[wallace.scala 71:19]
  assign FullAdder_1037_io_a = io_pp_3[38]; // @[wallace.scala 69:18]
  assign FullAdder_1037_io_b = io_pp_4[37]; // @[wallace.scala 70:18]
  assign FullAdder_1037_io_ci = io_pp_5[36]; // @[wallace.scala 71:19]
  assign FullAdder_1038_io_a = io_pp_6[35]; // @[wallace.scala 69:18]
  assign FullAdder_1038_io_b = io_pp_7[34]; // @[wallace.scala 70:18]
  assign FullAdder_1038_io_ci = io_pp_8[33]; // @[wallace.scala 71:19]
  assign FullAdder_1039_io_a = io_pp_9[32]; // @[wallace.scala 69:18]
  assign FullAdder_1039_io_b = io_pp_10[31]; // @[wallace.scala 70:18]
  assign FullAdder_1039_io_ci = io_pp_11[30]; // @[wallace.scala 71:19]
  assign FullAdder_1040_io_a = io_pp_12[29]; // @[wallace.scala 69:18]
  assign FullAdder_1040_io_b = io_pp_13[28]; // @[wallace.scala 70:18]
  assign FullAdder_1040_io_ci = io_pp_14[27]; // @[wallace.scala 71:19]
  assign FullAdder_1041_io_a = io_pp_15[26]; // @[wallace.scala 69:18]
  assign FullAdder_1041_io_b = io_pp_16[25]; // @[wallace.scala 70:18]
  assign FullAdder_1041_io_ci = io_pp_17[24]; // @[wallace.scala 71:19]
  assign FullAdder_1042_io_a = io_pp_18[23]; // @[wallace.scala 69:18]
  assign FullAdder_1042_io_b = io_pp_19[22]; // @[wallace.scala 70:18]
  assign FullAdder_1042_io_ci = io_pp_20[21]; // @[wallace.scala 71:19]
  assign FullAdder_1043_io_a = io_pp_21[20]; // @[wallace.scala 69:18]
  assign FullAdder_1043_io_b = io_pp_22[19]; // @[wallace.scala 70:18]
  assign FullAdder_1043_io_ci = io_pp_23[18]; // @[wallace.scala 71:19]
  assign FullAdder_1044_io_a = io_pp_24[17]; // @[wallace.scala 69:18]
  assign FullAdder_1044_io_b = io_pp_25[16]; // @[wallace.scala 70:18]
  assign FullAdder_1044_io_ci = io_pp_26[15]; // @[wallace.scala 71:19]
  assign FullAdder_1045_io_a = io_pp_27[14]; // @[wallace.scala 69:18]
  assign FullAdder_1045_io_b = io_pp_28[13]; // @[wallace.scala 70:18]
  assign FullAdder_1045_io_ci = io_pp_29[12]; // @[wallace.scala 71:19]
  assign FullAdder_1046_io_a = io_pp_30[11]; // @[wallace.scala 69:18]
  assign FullAdder_1046_io_b = io_pp_31[10]; // @[wallace.scala 70:18]
  assign FullAdder_1046_io_ci = io_pp_32[9]; // @[wallace.scala 71:19]
  assign FullAdder_1047_io_a = io_pp_33[8]; // @[wallace.scala 69:18]
  assign FullAdder_1047_io_b = io_pp_34[7]; // @[wallace.scala 70:18]
  assign FullAdder_1047_io_ci = io_pp_35[6]; // @[wallace.scala 71:19]
  assign FullAdder_1048_io_a = io_pp_36[5]; // @[wallace.scala 69:18]
  assign FullAdder_1048_io_b = io_pp_37[4]; // @[wallace.scala 70:18]
  assign FullAdder_1048_io_ci = io_pp_38[3]; // @[wallace.scala 71:19]
  assign FullAdder_1049_io_a = io_pp_39[2]; // @[wallace.scala 69:18]
  assign FullAdder_1049_io_b = io_pp_40[1]; // @[wallace.scala 70:18]
  assign FullAdder_1049_io_ci = io_pp_41[0]; // @[wallace.scala 71:19]
  assign FullAdder_1050_io_a = io_pp_0[40]; // @[wallace.scala 69:18]
  assign FullAdder_1050_io_b = io_pp_1[39]; // @[wallace.scala 70:18]
  assign FullAdder_1050_io_ci = io_pp_2[38]; // @[wallace.scala 71:19]
  assign FullAdder_1051_io_a = io_pp_3[37]; // @[wallace.scala 69:18]
  assign FullAdder_1051_io_b = io_pp_4[36]; // @[wallace.scala 70:18]
  assign FullAdder_1051_io_ci = io_pp_5[35]; // @[wallace.scala 71:19]
  assign FullAdder_1052_io_a = io_pp_6[34]; // @[wallace.scala 69:18]
  assign FullAdder_1052_io_b = io_pp_7[33]; // @[wallace.scala 70:18]
  assign FullAdder_1052_io_ci = io_pp_8[32]; // @[wallace.scala 71:19]
  assign FullAdder_1053_io_a = io_pp_9[31]; // @[wallace.scala 69:18]
  assign FullAdder_1053_io_b = io_pp_10[30]; // @[wallace.scala 70:18]
  assign FullAdder_1053_io_ci = io_pp_11[29]; // @[wallace.scala 71:19]
  assign FullAdder_1054_io_a = io_pp_12[28]; // @[wallace.scala 69:18]
  assign FullAdder_1054_io_b = io_pp_13[27]; // @[wallace.scala 70:18]
  assign FullAdder_1054_io_ci = io_pp_14[26]; // @[wallace.scala 71:19]
  assign FullAdder_1055_io_a = io_pp_15[25]; // @[wallace.scala 69:18]
  assign FullAdder_1055_io_b = io_pp_16[24]; // @[wallace.scala 70:18]
  assign FullAdder_1055_io_ci = io_pp_17[23]; // @[wallace.scala 71:19]
  assign FullAdder_1056_io_a = io_pp_18[22]; // @[wallace.scala 69:18]
  assign FullAdder_1056_io_b = io_pp_19[21]; // @[wallace.scala 70:18]
  assign FullAdder_1056_io_ci = io_pp_20[20]; // @[wallace.scala 71:19]
  assign FullAdder_1057_io_a = io_pp_21[19]; // @[wallace.scala 69:18]
  assign FullAdder_1057_io_b = io_pp_22[18]; // @[wallace.scala 70:18]
  assign FullAdder_1057_io_ci = io_pp_23[17]; // @[wallace.scala 71:19]
  assign FullAdder_1058_io_a = io_pp_24[16]; // @[wallace.scala 69:18]
  assign FullAdder_1058_io_b = io_pp_25[15]; // @[wallace.scala 70:18]
  assign FullAdder_1058_io_ci = io_pp_26[14]; // @[wallace.scala 71:19]
  assign FullAdder_1059_io_a = io_pp_27[13]; // @[wallace.scala 69:18]
  assign FullAdder_1059_io_b = io_pp_28[12]; // @[wallace.scala 70:18]
  assign FullAdder_1059_io_ci = io_pp_29[11]; // @[wallace.scala 71:19]
  assign FullAdder_1060_io_a = io_pp_30[10]; // @[wallace.scala 69:18]
  assign FullAdder_1060_io_b = io_pp_31[9]; // @[wallace.scala 70:18]
  assign FullAdder_1060_io_ci = io_pp_32[8]; // @[wallace.scala 71:19]
  assign FullAdder_1061_io_a = io_pp_33[7]; // @[wallace.scala 69:18]
  assign FullAdder_1061_io_b = io_pp_34[6]; // @[wallace.scala 70:18]
  assign FullAdder_1061_io_ci = io_pp_35[5]; // @[wallace.scala 71:19]
  assign FullAdder_1062_io_a = io_pp_36[4]; // @[wallace.scala 69:18]
  assign FullAdder_1062_io_b = io_pp_37[3]; // @[wallace.scala 70:18]
  assign FullAdder_1062_io_ci = io_pp_38[2]; // @[wallace.scala 71:19]
  assign FullAdder_1063_io_a = io_pp_0[39]; // @[wallace.scala 69:18]
  assign FullAdder_1063_io_b = io_pp_1[38]; // @[wallace.scala 70:18]
  assign FullAdder_1063_io_ci = io_pp_2[37]; // @[wallace.scala 71:19]
  assign FullAdder_1064_io_a = io_pp_3[36]; // @[wallace.scala 69:18]
  assign FullAdder_1064_io_b = io_pp_4[35]; // @[wallace.scala 70:18]
  assign FullAdder_1064_io_ci = io_pp_5[34]; // @[wallace.scala 71:19]
  assign FullAdder_1065_io_a = io_pp_6[33]; // @[wallace.scala 69:18]
  assign FullAdder_1065_io_b = io_pp_7[32]; // @[wallace.scala 70:18]
  assign FullAdder_1065_io_ci = io_pp_8[31]; // @[wallace.scala 71:19]
  assign FullAdder_1066_io_a = io_pp_9[30]; // @[wallace.scala 69:18]
  assign FullAdder_1066_io_b = io_pp_10[29]; // @[wallace.scala 70:18]
  assign FullAdder_1066_io_ci = io_pp_11[28]; // @[wallace.scala 71:19]
  assign FullAdder_1067_io_a = io_pp_12[27]; // @[wallace.scala 69:18]
  assign FullAdder_1067_io_b = io_pp_13[26]; // @[wallace.scala 70:18]
  assign FullAdder_1067_io_ci = io_pp_14[25]; // @[wallace.scala 71:19]
  assign FullAdder_1068_io_a = io_pp_15[24]; // @[wallace.scala 69:18]
  assign FullAdder_1068_io_b = io_pp_16[23]; // @[wallace.scala 70:18]
  assign FullAdder_1068_io_ci = io_pp_17[22]; // @[wallace.scala 71:19]
  assign FullAdder_1069_io_a = io_pp_18[21]; // @[wallace.scala 69:18]
  assign FullAdder_1069_io_b = io_pp_19[20]; // @[wallace.scala 70:18]
  assign FullAdder_1069_io_ci = io_pp_20[19]; // @[wallace.scala 71:19]
  assign FullAdder_1070_io_a = io_pp_21[18]; // @[wallace.scala 69:18]
  assign FullAdder_1070_io_b = io_pp_22[17]; // @[wallace.scala 70:18]
  assign FullAdder_1070_io_ci = io_pp_23[16]; // @[wallace.scala 71:19]
  assign FullAdder_1071_io_a = io_pp_24[15]; // @[wallace.scala 69:18]
  assign FullAdder_1071_io_b = io_pp_25[14]; // @[wallace.scala 70:18]
  assign FullAdder_1071_io_ci = io_pp_26[13]; // @[wallace.scala 71:19]
  assign FullAdder_1072_io_a = io_pp_27[12]; // @[wallace.scala 69:18]
  assign FullAdder_1072_io_b = io_pp_28[11]; // @[wallace.scala 70:18]
  assign FullAdder_1072_io_ci = io_pp_29[10]; // @[wallace.scala 71:19]
  assign FullAdder_1073_io_a = io_pp_30[9]; // @[wallace.scala 69:18]
  assign FullAdder_1073_io_b = io_pp_31[8]; // @[wallace.scala 70:18]
  assign FullAdder_1073_io_ci = io_pp_32[7]; // @[wallace.scala 71:19]
  assign FullAdder_1074_io_a = io_pp_33[6]; // @[wallace.scala 69:18]
  assign FullAdder_1074_io_b = io_pp_34[5]; // @[wallace.scala 70:18]
  assign FullAdder_1074_io_ci = io_pp_35[4]; // @[wallace.scala 71:19]
  assign FullAdder_1075_io_a = io_pp_36[3]; // @[wallace.scala 69:18]
  assign FullAdder_1075_io_b = io_pp_37[2]; // @[wallace.scala 70:18]
  assign FullAdder_1075_io_ci = io_pp_38[1]; // @[wallace.scala 71:19]
  assign FullAdder_1076_io_a = io_pp_0[38]; // @[wallace.scala 69:18]
  assign FullAdder_1076_io_b = io_pp_1[37]; // @[wallace.scala 70:18]
  assign FullAdder_1076_io_ci = io_pp_2[36]; // @[wallace.scala 71:19]
  assign FullAdder_1077_io_a = io_pp_3[35]; // @[wallace.scala 69:18]
  assign FullAdder_1077_io_b = io_pp_4[34]; // @[wallace.scala 70:18]
  assign FullAdder_1077_io_ci = io_pp_5[33]; // @[wallace.scala 71:19]
  assign FullAdder_1078_io_a = io_pp_6[32]; // @[wallace.scala 69:18]
  assign FullAdder_1078_io_b = io_pp_7[31]; // @[wallace.scala 70:18]
  assign FullAdder_1078_io_ci = io_pp_8[30]; // @[wallace.scala 71:19]
  assign FullAdder_1079_io_a = io_pp_9[29]; // @[wallace.scala 69:18]
  assign FullAdder_1079_io_b = io_pp_10[28]; // @[wallace.scala 70:18]
  assign FullAdder_1079_io_ci = io_pp_11[27]; // @[wallace.scala 71:19]
  assign FullAdder_1080_io_a = io_pp_12[26]; // @[wallace.scala 69:18]
  assign FullAdder_1080_io_b = io_pp_13[25]; // @[wallace.scala 70:18]
  assign FullAdder_1080_io_ci = io_pp_14[24]; // @[wallace.scala 71:19]
  assign FullAdder_1081_io_a = io_pp_15[23]; // @[wallace.scala 69:18]
  assign FullAdder_1081_io_b = io_pp_16[22]; // @[wallace.scala 70:18]
  assign FullAdder_1081_io_ci = io_pp_17[21]; // @[wallace.scala 71:19]
  assign FullAdder_1082_io_a = io_pp_18[20]; // @[wallace.scala 69:18]
  assign FullAdder_1082_io_b = io_pp_19[19]; // @[wallace.scala 70:18]
  assign FullAdder_1082_io_ci = io_pp_20[18]; // @[wallace.scala 71:19]
  assign FullAdder_1083_io_a = io_pp_21[17]; // @[wallace.scala 69:18]
  assign FullAdder_1083_io_b = io_pp_22[16]; // @[wallace.scala 70:18]
  assign FullAdder_1083_io_ci = io_pp_23[15]; // @[wallace.scala 71:19]
  assign FullAdder_1084_io_a = io_pp_24[14]; // @[wallace.scala 69:18]
  assign FullAdder_1084_io_b = io_pp_25[13]; // @[wallace.scala 70:18]
  assign FullAdder_1084_io_ci = io_pp_26[12]; // @[wallace.scala 71:19]
  assign FullAdder_1085_io_a = io_pp_27[11]; // @[wallace.scala 69:18]
  assign FullAdder_1085_io_b = io_pp_28[10]; // @[wallace.scala 70:18]
  assign FullAdder_1085_io_ci = io_pp_29[9]; // @[wallace.scala 71:19]
  assign FullAdder_1086_io_a = io_pp_30[8]; // @[wallace.scala 69:18]
  assign FullAdder_1086_io_b = io_pp_31[7]; // @[wallace.scala 70:18]
  assign FullAdder_1086_io_ci = io_pp_32[6]; // @[wallace.scala 71:19]
  assign FullAdder_1087_io_a = io_pp_33[5]; // @[wallace.scala 69:18]
  assign FullAdder_1087_io_b = io_pp_34[4]; // @[wallace.scala 70:18]
  assign FullAdder_1087_io_ci = io_pp_35[3]; // @[wallace.scala 71:19]
  assign FullAdder_1088_io_a = io_pp_36[2]; // @[wallace.scala 69:18]
  assign FullAdder_1088_io_b = io_pp_37[1]; // @[wallace.scala 70:18]
  assign FullAdder_1088_io_ci = io_pp_38[0]; // @[wallace.scala 71:19]
  assign FullAdder_1089_io_a = io_pp_0[37]; // @[wallace.scala 69:18]
  assign FullAdder_1089_io_b = io_pp_1[36]; // @[wallace.scala 70:18]
  assign FullAdder_1089_io_ci = io_pp_2[35]; // @[wallace.scala 71:19]
  assign FullAdder_1090_io_a = io_pp_3[34]; // @[wallace.scala 69:18]
  assign FullAdder_1090_io_b = io_pp_4[33]; // @[wallace.scala 70:18]
  assign FullAdder_1090_io_ci = io_pp_5[32]; // @[wallace.scala 71:19]
  assign FullAdder_1091_io_a = io_pp_6[31]; // @[wallace.scala 69:18]
  assign FullAdder_1091_io_b = io_pp_7[30]; // @[wallace.scala 70:18]
  assign FullAdder_1091_io_ci = io_pp_8[29]; // @[wallace.scala 71:19]
  assign FullAdder_1092_io_a = io_pp_9[28]; // @[wallace.scala 69:18]
  assign FullAdder_1092_io_b = io_pp_10[27]; // @[wallace.scala 70:18]
  assign FullAdder_1092_io_ci = io_pp_11[26]; // @[wallace.scala 71:19]
  assign FullAdder_1093_io_a = io_pp_12[25]; // @[wallace.scala 69:18]
  assign FullAdder_1093_io_b = io_pp_13[24]; // @[wallace.scala 70:18]
  assign FullAdder_1093_io_ci = io_pp_14[23]; // @[wallace.scala 71:19]
  assign FullAdder_1094_io_a = io_pp_15[22]; // @[wallace.scala 69:18]
  assign FullAdder_1094_io_b = io_pp_16[21]; // @[wallace.scala 70:18]
  assign FullAdder_1094_io_ci = io_pp_17[20]; // @[wallace.scala 71:19]
  assign FullAdder_1095_io_a = io_pp_18[19]; // @[wallace.scala 69:18]
  assign FullAdder_1095_io_b = io_pp_19[18]; // @[wallace.scala 70:18]
  assign FullAdder_1095_io_ci = io_pp_20[17]; // @[wallace.scala 71:19]
  assign FullAdder_1096_io_a = io_pp_21[16]; // @[wallace.scala 69:18]
  assign FullAdder_1096_io_b = io_pp_22[15]; // @[wallace.scala 70:18]
  assign FullAdder_1096_io_ci = io_pp_23[14]; // @[wallace.scala 71:19]
  assign FullAdder_1097_io_a = io_pp_24[13]; // @[wallace.scala 69:18]
  assign FullAdder_1097_io_b = io_pp_25[12]; // @[wallace.scala 70:18]
  assign FullAdder_1097_io_ci = io_pp_26[11]; // @[wallace.scala 71:19]
  assign FullAdder_1098_io_a = io_pp_27[10]; // @[wallace.scala 69:18]
  assign FullAdder_1098_io_b = io_pp_28[9]; // @[wallace.scala 70:18]
  assign FullAdder_1098_io_ci = io_pp_29[8]; // @[wallace.scala 71:19]
  assign FullAdder_1099_io_a = io_pp_30[7]; // @[wallace.scala 69:18]
  assign FullAdder_1099_io_b = io_pp_31[6]; // @[wallace.scala 70:18]
  assign FullAdder_1099_io_ci = io_pp_32[5]; // @[wallace.scala 71:19]
  assign FullAdder_1100_io_a = io_pp_33[4]; // @[wallace.scala 69:18]
  assign FullAdder_1100_io_b = io_pp_34[3]; // @[wallace.scala 70:18]
  assign FullAdder_1100_io_ci = io_pp_35[2]; // @[wallace.scala 71:19]
  assign HalfAdder_22_io_a = io_pp_36[1]; // @[wallace.scala 59:18]
  assign HalfAdder_22_io_b = io_pp_37[0]; // @[wallace.scala 60:18]
  assign FullAdder_1101_io_a = io_pp_0[36]; // @[wallace.scala 69:18]
  assign FullAdder_1101_io_b = io_pp_1[35]; // @[wallace.scala 70:18]
  assign FullAdder_1101_io_ci = io_pp_2[34]; // @[wallace.scala 71:19]
  assign FullAdder_1102_io_a = io_pp_3[33]; // @[wallace.scala 69:18]
  assign FullAdder_1102_io_b = io_pp_4[32]; // @[wallace.scala 70:18]
  assign FullAdder_1102_io_ci = io_pp_5[31]; // @[wallace.scala 71:19]
  assign FullAdder_1103_io_a = io_pp_6[30]; // @[wallace.scala 69:18]
  assign FullAdder_1103_io_b = io_pp_7[29]; // @[wallace.scala 70:18]
  assign FullAdder_1103_io_ci = io_pp_8[28]; // @[wallace.scala 71:19]
  assign FullAdder_1104_io_a = io_pp_9[27]; // @[wallace.scala 69:18]
  assign FullAdder_1104_io_b = io_pp_10[26]; // @[wallace.scala 70:18]
  assign FullAdder_1104_io_ci = io_pp_11[25]; // @[wallace.scala 71:19]
  assign FullAdder_1105_io_a = io_pp_12[24]; // @[wallace.scala 69:18]
  assign FullAdder_1105_io_b = io_pp_13[23]; // @[wallace.scala 70:18]
  assign FullAdder_1105_io_ci = io_pp_14[22]; // @[wallace.scala 71:19]
  assign FullAdder_1106_io_a = io_pp_15[21]; // @[wallace.scala 69:18]
  assign FullAdder_1106_io_b = io_pp_16[20]; // @[wallace.scala 70:18]
  assign FullAdder_1106_io_ci = io_pp_17[19]; // @[wallace.scala 71:19]
  assign FullAdder_1107_io_a = io_pp_18[18]; // @[wallace.scala 69:18]
  assign FullAdder_1107_io_b = io_pp_19[17]; // @[wallace.scala 70:18]
  assign FullAdder_1107_io_ci = io_pp_20[16]; // @[wallace.scala 71:19]
  assign FullAdder_1108_io_a = io_pp_21[15]; // @[wallace.scala 69:18]
  assign FullAdder_1108_io_b = io_pp_22[14]; // @[wallace.scala 70:18]
  assign FullAdder_1108_io_ci = io_pp_23[13]; // @[wallace.scala 71:19]
  assign FullAdder_1109_io_a = io_pp_24[12]; // @[wallace.scala 69:18]
  assign FullAdder_1109_io_b = io_pp_25[11]; // @[wallace.scala 70:18]
  assign FullAdder_1109_io_ci = io_pp_26[10]; // @[wallace.scala 71:19]
  assign FullAdder_1110_io_a = io_pp_27[9]; // @[wallace.scala 69:18]
  assign FullAdder_1110_io_b = io_pp_28[8]; // @[wallace.scala 70:18]
  assign FullAdder_1110_io_ci = io_pp_29[7]; // @[wallace.scala 71:19]
  assign FullAdder_1111_io_a = io_pp_30[6]; // @[wallace.scala 69:18]
  assign FullAdder_1111_io_b = io_pp_31[5]; // @[wallace.scala 70:18]
  assign FullAdder_1111_io_ci = io_pp_32[4]; // @[wallace.scala 71:19]
  assign FullAdder_1112_io_a = io_pp_33[3]; // @[wallace.scala 69:18]
  assign FullAdder_1112_io_b = io_pp_34[2]; // @[wallace.scala 70:18]
  assign FullAdder_1112_io_ci = io_pp_35[1]; // @[wallace.scala 71:19]
  assign FullAdder_1113_io_a = io_pp_0[35]; // @[wallace.scala 69:18]
  assign FullAdder_1113_io_b = io_pp_1[34]; // @[wallace.scala 70:18]
  assign FullAdder_1113_io_ci = io_pp_2[33]; // @[wallace.scala 71:19]
  assign FullAdder_1114_io_a = io_pp_3[32]; // @[wallace.scala 69:18]
  assign FullAdder_1114_io_b = io_pp_4[31]; // @[wallace.scala 70:18]
  assign FullAdder_1114_io_ci = io_pp_5[30]; // @[wallace.scala 71:19]
  assign FullAdder_1115_io_a = io_pp_6[29]; // @[wallace.scala 69:18]
  assign FullAdder_1115_io_b = io_pp_7[28]; // @[wallace.scala 70:18]
  assign FullAdder_1115_io_ci = io_pp_8[27]; // @[wallace.scala 71:19]
  assign FullAdder_1116_io_a = io_pp_9[26]; // @[wallace.scala 69:18]
  assign FullAdder_1116_io_b = io_pp_10[25]; // @[wallace.scala 70:18]
  assign FullAdder_1116_io_ci = io_pp_11[24]; // @[wallace.scala 71:19]
  assign FullAdder_1117_io_a = io_pp_12[23]; // @[wallace.scala 69:18]
  assign FullAdder_1117_io_b = io_pp_13[22]; // @[wallace.scala 70:18]
  assign FullAdder_1117_io_ci = io_pp_14[21]; // @[wallace.scala 71:19]
  assign FullAdder_1118_io_a = io_pp_15[20]; // @[wallace.scala 69:18]
  assign FullAdder_1118_io_b = io_pp_16[19]; // @[wallace.scala 70:18]
  assign FullAdder_1118_io_ci = io_pp_17[18]; // @[wallace.scala 71:19]
  assign FullAdder_1119_io_a = io_pp_18[17]; // @[wallace.scala 69:18]
  assign FullAdder_1119_io_b = io_pp_19[16]; // @[wallace.scala 70:18]
  assign FullAdder_1119_io_ci = io_pp_20[15]; // @[wallace.scala 71:19]
  assign FullAdder_1120_io_a = io_pp_21[14]; // @[wallace.scala 69:18]
  assign FullAdder_1120_io_b = io_pp_22[13]; // @[wallace.scala 70:18]
  assign FullAdder_1120_io_ci = io_pp_23[12]; // @[wallace.scala 71:19]
  assign FullAdder_1121_io_a = io_pp_24[11]; // @[wallace.scala 69:18]
  assign FullAdder_1121_io_b = io_pp_25[10]; // @[wallace.scala 70:18]
  assign FullAdder_1121_io_ci = io_pp_26[9]; // @[wallace.scala 71:19]
  assign FullAdder_1122_io_a = io_pp_27[8]; // @[wallace.scala 69:18]
  assign FullAdder_1122_io_b = io_pp_28[7]; // @[wallace.scala 70:18]
  assign FullAdder_1122_io_ci = io_pp_29[6]; // @[wallace.scala 71:19]
  assign FullAdder_1123_io_a = io_pp_30[5]; // @[wallace.scala 69:18]
  assign FullAdder_1123_io_b = io_pp_31[4]; // @[wallace.scala 70:18]
  assign FullAdder_1123_io_ci = io_pp_32[3]; // @[wallace.scala 71:19]
  assign FullAdder_1124_io_a = io_pp_33[2]; // @[wallace.scala 69:18]
  assign FullAdder_1124_io_b = io_pp_34[1]; // @[wallace.scala 70:18]
  assign FullAdder_1124_io_ci = io_pp_35[0]; // @[wallace.scala 71:19]
  assign FullAdder_1125_io_a = io_pp_0[34]; // @[wallace.scala 69:18]
  assign FullAdder_1125_io_b = io_pp_1[33]; // @[wallace.scala 70:18]
  assign FullAdder_1125_io_ci = io_pp_2[32]; // @[wallace.scala 71:19]
  assign FullAdder_1126_io_a = io_pp_3[31]; // @[wallace.scala 69:18]
  assign FullAdder_1126_io_b = io_pp_4[30]; // @[wallace.scala 70:18]
  assign FullAdder_1126_io_ci = io_pp_5[29]; // @[wallace.scala 71:19]
  assign FullAdder_1127_io_a = io_pp_6[28]; // @[wallace.scala 69:18]
  assign FullAdder_1127_io_b = io_pp_7[27]; // @[wallace.scala 70:18]
  assign FullAdder_1127_io_ci = io_pp_8[26]; // @[wallace.scala 71:19]
  assign FullAdder_1128_io_a = io_pp_9[25]; // @[wallace.scala 69:18]
  assign FullAdder_1128_io_b = io_pp_10[24]; // @[wallace.scala 70:18]
  assign FullAdder_1128_io_ci = io_pp_11[23]; // @[wallace.scala 71:19]
  assign FullAdder_1129_io_a = io_pp_12[22]; // @[wallace.scala 69:18]
  assign FullAdder_1129_io_b = io_pp_13[21]; // @[wallace.scala 70:18]
  assign FullAdder_1129_io_ci = io_pp_14[20]; // @[wallace.scala 71:19]
  assign FullAdder_1130_io_a = io_pp_15[19]; // @[wallace.scala 69:18]
  assign FullAdder_1130_io_b = io_pp_16[18]; // @[wallace.scala 70:18]
  assign FullAdder_1130_io_ci = io_pp_17[17]; // @[wallace.scala 71:19]
  assign FullAdder_1131_io_a = io_pp_18[16]; // @[wallace.scala 69:18]
  assign FullAdder_1131_io_b = io_pp_19[15]; // @[wallace.scala 70:18]
  assign FullAdder_1131_io_ci = io_pp_20[14]; // @[wallace.scala 71:19]
  assign FullAdder_1132_io_a = io_pp_21[13]; // @[wallace.scala 69:18]
  assign FullAdder_1132_io_b = io_pp_22[12]; // @[wallace.scala 70:18]
  assign FullAdder_1132_io_ci = io_pp_23[11]; // @[wallace.scala 71:19]
  assign FullAdder_1133_io_a = io_pp_24[10]; // @[wallace.scala 69:18]
  assign FullAdder_1133_io_b = io_pp_25[9]; // @[wallace.scala 70:18]
  assign FullAdder_1133_io_ci = io_pp_26[8]; // @[wallace.scala 71:19]
  assign FullAdder_1134_io_a = io_pp_27[7]; // @[wallace.scala 69:18]
  assign FullAdder_1134_io_b = io_pp_28[6]; // @[wallace.scala 70:18]
  assign FullAdder_1134_io_ci = io_pp_29[5]; // @[wallace.scala 71:19]
  assign FullAdder_1135_io_a = io_pp_30[4]; // @[wallace.scala 69:18]
  assign FullAdder_1135_io_b = io_pp_31[3]; // @[wallace.scala 70:18]
  assign FullAdder_1135_io_ci = io_pp_32[2]; // @[wallace.scala 71:19]
  assign HalfAdder_23_io_a = io_pp_33[1]; // @[wallace.scala 59:18]
  assign HalfAdder_23_io_b = io_pp_34[0]; // @[wallace.scala 60:18]
  assign FullAdder_1136_io_a = io_pp_0[33]; // @[wallace.scala 69:18]
  assign FullAdder_1136_io_b = io_pp_1[32]; // @[wallace.scala 70:18]
  assign FullAdder_1136_io_ci = io_pp_2[31]; // @[wallace.scala 71:19]
  assign FullAdder_1137_io_a = io_pp_3[30]; // @[wallace.scala 69:18]
  assign FullAdder_1137_io_b = io_pp_4[29]; // @[wallace.scala 70:18]
  assign FullAdder_1137_io_ci = io_pp_5[28]; // @[wallace.scala 71:19]
  assign FullAdder_1138_io_a = io_pp_6[27]; // @[wallace.scala 69:18]
  assign FullAdder_1138_io_b = io_pp_7[26]; // @[wallace.scala 70:18]
  assign FullAdder_1138_io_ci = io_pp_8[25]; // @[wallace.scala 71:19]
  assign FullAdder_1139_io_a = io_pp_9[24]; // @[wallace.scala 69:18]
  assign FullAdder_1139_io_b = io_pp_10[23]; // @[wallace.scala 70:18]
  assign FullAdder_1139_io_ci = io_pp_11[22]; // @[wallace.scala 71:19]
  assign FullAdder_1140_io_a = io_pp_12[21]; // @[wallace.scala 69:18]
  assign FullAdder_1140_io_b = io_pp_13[20]; // @[wallace.scala 70:18]
  assign FullAdder_1140_io_ci = io_pp_14[19]; // @[wallace.scala 71:19]
  assign FullAdder_1141_io_a = io_pp_15[18]; // @[wallace.scala 69:18]
  assign FullAdder_1141_io_b = io_pp_16[17]; // @[wallace.scala 70:18]
  assign FullAdder_1141_io_ci = io_pp_17[16]; // @[wallace.scala 71:19]
  assign FullAdder_1142_io_a = io_pp_18[15]; // @[wallace.scala 69:18]
  assign FullAdder_1142_io_b = io_pp_19[14]; // @[wallace.scala 70:18]
  assign FullAdder_1142_io_ci = io_pp_20[13]; // @[wallace.scala 71:19]
  assign FullAdder_1143_io_a = io_pp_21[12]; // @[wallace.scala 69:18]
  assign FullAdder_1143_io_b = io_pp_22[11]; // @[wallace.scala 70:18]
  assign FullAdder_1143_io_ci = io_pp_23[10]; // @[wallace.scala 71:19]
  assign FullAdder_1144_io_a = io_pp_24[9]; // @[wallace.scala 69:18]
  assign FullAdder_1144_io_b = io_pp_25[8]; // @[wallace.scala 70:18]
  assign FullAdder_1144_io_ci = io_pp_26[7]; // @[wallace.scala 71:19]
  assign FullAdder_1145_io_a = io_pp_27[6]; // @[wallace.scala 69:18]
  assign FullAdder_1145_io_b = io_pp_28[5]; // @[wallace.scala 70:18]
  assign FullAdder_1145_io_ci = io_pp_29[4]; // @[wallace.scala 71:19]
  assign FullAdder_1146_io_a = io_pp_30[3]; // @[wallace.scala 69:18]
  assign FullAdder_1146_io_b = io_pp_31[2]; // @[wallace.scala 70:18]
  assign FullAdder_1146_io_ci = io_pp_32[1]; // @[wallace.scala 71:19]
  assign FullAdder_1147_io_a = io_pp_0[32]; // @[wallace.scala 69:18]
  assign FullAdder_1147_io_b = io_pp_1[31]; // @[wallace.scala 70:18]
  assign FullAdder_1147_io_ci = io_pp_2[30]; // @[wallace.scala 71:19]
  assign FullAdder_1148_io_a = io_pp_3[29]; // @[wallace.scala 69:18]
  assign FullAdder_1148_io_b = io_pp_4[28]; // @[wallace.scala 70:18]
  assign FullAdder_1148_io_ci = io_pp_5[27]; // @[wallace.scala 71:19]
  assign FullAdder_1149_io_a = io_pp_6[26]; // @[wallace.scala 69:18]
  assign FullAdder_1149_io_b = io_pp_7[25]; // @[wallace.scala 70:18]
  assign FullAdder_1149_io_ci = io_pp_8[24]; // @[wallace.scala 71:19]
  assign FullAdder_1150_io_a = io_pp_9[23]; // @[wallace.scala 69:18]
  assign FullAdder_1150_io_b = io_pp_10[22]; // @[wallace.scala 70:18]
  assign FullAdder_1150_io_ci = io_pp_11[21]; // @[wallace.scala 71:19]
  assign FullAdder_1151_io_a = io_pp_12[20]; // @[wallace.scala 69:18]
  assign FullAdder_1151_io_b = io_pp_13[19]; // @[wallace.scala 70:18]
  assign FullAdder_1151_io_ci = io_pp_14[18]; // @[wallace.scala 71:19]
  assign FullAdder_1152_io_a = io_pp_15[17]; // @[wallace.scala 69:18]
  assign FullAdder_1152_io_b = io_pp_16[16]; // @[wallace.scala 70:18]
  assign FullAdder_1152_io_ci = io_pp_17[15]; // @[wallace.scala 71:19]
  assign FullAdder_1153_io_a = io_pp_18[14]; // @[wallace.scala 69:18]
  assign FullAdder_1153_io_b = io_pp_19[13]; // @[wallace.scala 70:18]
  assign FullAdder_1153_io_ci = io_pp_20[12]; // @[wallace.scala 71:19]
  assign FullAdder_1154_io_a = io_pp_21[11]; // @[wallace.scala 69:18]
  assign FullAdder_1154_io_b = io_pp_22[10]; // @[wallace.scala 70:18]
  assign FullAdder_1154_io_ci = io_pp_23[9]; // @[wallace.scala 71:19]
  assign FullAdder_1155_io_a = io_pp_24[8]; // @[wallace.scala 69:18]
  assign FullAdder_1155_io_b = io_pp_25[7]; // @[wallace.scala 70:18]
  assign FullAdder_1155_io_ci = io_pp_26[6]; // @[wallace.scala 71:19]
  assign FullAdder_1156_io_a = io_pp_27[5]; // @[wallace.scala 69:18]
  assign FullAdder_1156_io_b = io_pp_28[4]; // @[wallace.scala 70:18]
  assign FullAdder_1156_io_ci = io_pp_29[3]; // @[wallace.scala 71:19]
  assign FullAdder_1157_io_a = io_pp_30[2]; // @[wallace.scala 69:18]
  assign FullAdder_1157_io_b = io_pp_31[1]; // @[wallace.scala 70:18]
  assign FullAdder_1157_io_ci = io_pp_32[0]; // @[wallace.scala 71:19]
  assign FullAdder_1158_io_a = io_pp_0[31]; // @[wallace.scala 69:18]
  assign FullAdder_1158_io_b = io_pp_1[30]; // @[wallace.scala 70:18]
  assign FullAdder_1158_io_ci = io_pp_2[29]; // @[wallace.scala 71:19]
  assign FullAdder_1159_io_a = io_pp_3[28]; // @[wallace.scala 69:18]
  assign FullAdder_1159_io_b = io_pp_4[27]; // @[wallace.scala 70:18]
  assign FullAdder_1159_io_ci = io_pp_5[26]; // @[wallace.scala 71:19]
  assign FullAdder_1160_io_a = io_pp_6[25]; // @[wallace.scala 69:18]
  assign FullAdder_1160_io_b = io_pp_7[24]; // @[wallace.scala 70:18]
  assign FullAdder_1160_io_ci = io_pp_8[23]; // @[wallace.scala 71:19]
  assign FullAdder_1161_io_a = io_pp_9[22]; // @[wallace.scala 69:18]
  assign FullAdder_1161_io_b = io_pp_10[21]; // @[wallace.scala 70:18]
  assign FullAdder_1161_io_ci = io_pp_11[20]; // @[wallace.scala 71:19]
  assign FullAdder_1162_io_a = io_pp_12[19]; // @[wallace.scala 69:18]
  assign FullAdder_1162_io_b = io_pp_13[18]; // @[wallace.scala 70:18]
  assign FullAdder_1162_io_ci = io_pp_14[17]; // @[wallace.scala 71:19]
  assign FullAdder_1163_io_a = io_pp_15[16]; // @[wallace.scala 69:18]
  assign FullAdder_1163_io_b = io_pp_16[15]; // @[wallace.scala 70:18]
  assign FullAdder_1163_io_ci = io_pp_17[14]; // @[wallace.scala 71:19]
  assign FullAdder_1164_io_a = io_pp_18[13]; // @[wallace.scala 69:18]
  assign FullAdder_1164_io_b = io_pp_19[12]; // @[wallace.scala 70:18]
  assign FullAdder_1164_io_ci = io_pp_20[11]; // @[wallace.scala 71:19]
  assign FullAdder_1165_io_a = io_pp_21[10]; // @[wallace.scala 69:18]
  assign FullAdder_1165_io_b = io_pp_22[9]; // @[wallace.scala 70:18]
  assign FullAdder_1165_io_ci = io_pp_23[8]; // @[wallace.scala 71:19]
  assign FullAdder_1166_io_a = io_pp_24[7]; // @[wallace.scala 69:18]
  assign FullAdder_1166_io_b = io_pp_25[6]; // @[wallace.scala 70:18]
  assign FullAdder_1166_io_ci = io_pp_26[5]; // @[wallace.scala 71:19]
  assign FullAdder_1167_io_a = io_pp_27[4]; // @[wallace.scala 69:18]
  assign FullAdder_1167_io_b = io_pp_28[3]; // @[wallace.scala 70:18]
  assign FullAdder_1167_io_ci = io_pp_29[2]; // @[wallace.scala 71:19]
  assign HalfAdder_24_io_a = io_pp_30[1]; // @[wallace.scala 59:18]
  assign HalfAdder_24_io_b = io_pp_31[0]; // @[wallace.scala 60:18]
  assign FullAdder_1168_io_a = io_pp_0[30]; // @[wallace.scala 69:18]
  assign FullAdder_1168_io_b = io_pp_1[29]; // @[wallace.scala 70:18]
  assign FullAdder_1168_io_ci = io_pp_2[28]; // @[wallace.scala 71:19]
  assign FullAdder_1169_io_a = io_pp_3[27]; // @[wallace.scala 69:18]
  assign FullAdder_1169_io_b = io_pp_4[26]; // @[wallace.scala 70:18]
  assign FullAdder_1169_io_ci = io_pp_5[25]; // @[wallace.scala 71:19]
  assign FullAdder_1170_io_a = io_pp_6[24]; // @[wallace.scala 69:18]
  assign FullAdder_1170_io_b = io_pp_7[23]; // @[wallace.scala 70:18]
  assign FullAdder_1170_io_ci = io_pp_8[22]; // @[wallace.scala 71:19]
  assign FullAdder_1171_io_a = io_pp_9[21]; // @[wallace.scala 69:18]
  assign FullAdder_1171_io_b = io_pp_10[20]; // @[wallace.scala 70:18]
  assign FullAdder_1171_io_ci = io_pp_11[19]; // @[wallace.scala 71:19]
  assign FullAdder_1172_io_a = io_pp_12[18]; // @[wallace.scala 69:18]
  assign FullAdder_1172_io_b = io_pp_13[17]; // @[wallace.scala 70:18]
  assign FullAdder_1172_io_ci = io_pp_14[16]; // @[wallace.scala 71:19]
  assign FullAdder_1173_io_a = io_pp_15[15]; // @[wallace.scala 69:18]
  assign FullAdder_1173_io_b = io_pp_16[14]; // @[wallace.scala 70:18]
  assign FullAdder_1173_io_ci = io_pp_17[13]; // @[wallace.scala 71:19]
  assign FullAdder_1174_io_a = io_pp_18[12]; // @[wallace.scala 69:18]
  assign FullAdder_1174_io_b = io_pp_19[11]; // @[wallace.scala 70:18]
  assign FullAdder_1174_io_ci = io_pp_20[10]; // @[wallace.scala 71:19]
  assign FullAdder_1175_io_a = io_pp_21[9]; // @[wallace.scala 69:18]
  assign FullAdder_1175_io_b = io_pp_22[8]; // @[wallace.scala 70:18]
  assign FullAdder_1175_io_ci = io_pp_23[7]; // @[wallace.scala 71:19]
  assign FullAdder_1176_io_a = io_pp_24[6]; // @[wallace.scala 69:18]
  assign FullAdder_1176_io_b = io_pp_25[5]; // @[wallace.scala 70:18]
  assign FullAdder_1176_io_ci = io_pp_26[4]; // @[wallace.scala 71:19]
  assign FullAdder_1177_io_a = io_pp_27[3]; // @[wallace.scala 69:18]
  assign FullAdder_1177_io_b = io_pp_28[2]; // @[wallace.scala 70:18]
  assign FullAdder_1177_io_ci = io_pp_29[1]; // @[wallace.scala 71:19]
  assign FullAdder_1178_io_a = io_pp_0[29]; // @[wallace.scala 69:18]
  assign FullAdder_1178_io_b = io_pp_1[28]; // @[wallace.scala 70:18]
  assign FullAdder_1178_io_ci = io_pp_2[27]; // @[wallace.scala 71:19]
  assign FullAdder_1179_io_a = io_pp_3[26]; // @[wallace.scala 69:18]
  assign FullAdder_1179_io_b = io_pp_4[25]; // @[wallace.scala 70:18]
  assign FullAdder_1179_io_ci = io_pp_5[24]; // @[wallace.scala 71:19]
  assign FullAdder_1180_io_a = io_pp_6[23]; // @[wallace.scala 69:18]
  assign FullAdder_1180_io_b = io_pp_7[22]; // @[wallace.scala 70:18]
  assign FullAdder_1180_io_ci = io_pp_8[21]; // @[wallace.scala 71:19]
  assign FullAdder_1181_io_a = io_pp_9[20]; // @[wallace.scala 69:18]
  assign FullAdder_1181_io_b = io_pp_10[19]; // @[wallace.scala 70:18]
  assign FullAdder_1181_io_ci = io_pp_11[18]; // @[wallace.scala 71:19]
  assign FullAdder_1182_io_a = io_pp_12[17]; // @[wallace.scala 69:18]
  assign FullAdder_1182_io_b = io_pp_13[16]; // @[wallace.scala 70:18]
  assign FullAdder_1182_io_ci = io_pp_14[15]; // @[wallace.scala 71:19]
  assign FullAdder_1183_io_a = io_pp_15[14]; // @[wallace.scala 69:18]
  assign FullAdder_1183_io_b = io_pp_16[13]; // @[wallace.scala 70:18]
  assign FullAdder_1183_io_ci = io_pp_17[12]; // @[wallace.scala 71:19]
  assign FullAdder_1184_io_a = io_pp_18[11]; // @[wallace.scala 69:18]
  assign FullAdder_1184_io_b = io_pp_19[10]; // @[wallace.scala 70:18]
  assign FullAdder_1184_io_ci = io_pp_20[9]; // @[wallace.scala 71:19]
  assign FullAdder_1185_io_a = io_pp_21[8]; // @[wallace.scala 69:18]
  assign FullAdder_1185_io_b = io_pp_22[7]; // @[wallace.scala 70:18]
  assign FullAdder_1185_io_ci = io_pp_23[6]; // @[wallace.scala 71:19]
  assign FullAdder_1186_io_a = io_pp_24[5]; // @[wallace.scala 69:18]
  assign FullAdder_1186_io_b = io_pp_25[4]; // @[wallace.scala 70:18]
  assign FullAdder_1186_io_ci = io_pp_26[3]; // @[wallace.scala 71:19]
  assign FullAdder_1187_io_a = io_pp_27[2]; // @[wallace.scala 69:18]
  assign FullAdder_1187_io_b = io_pp_28[1]; // @[wallace.scala 70:18]
  assign FullAdder_1187_io_ci = io_pp_29[0]; // @[wallace.scala 71:19]
  assign FullAdder_1188_io_a = io_pp_0[28]; // @[wallace.scala 69:18]
  assign FullAdder_1188_io_b = io_pp_1[27]; // @[wallace.scala 70:18]
  assign FullAdder_1188_io_ci = io_pp_2[26]; // @[wallace.scala 71:19]
  assign FullAdder_1189_io_a = io_pp_3[25]; // @[wallace.scala 69:18]
  assign FullAdder_1189_io_b = io_pp_4[24]; // @[wallace.scala 70:18]
  assign FullAdder_1189_io_ci = io_pp_5[23]; // @[wallace.scala 71:19]
  assign FullAdder_1190_io_a = io_pp_6[22]; // @[wallace.scala 69:18]
  assign FullAdder_1190_io_b = io_pp_7[21]; // @[wallace.scala 70:18]
  assign FullAdder_1190_io_ci = io_pp_8[20]; // @[wallace.scala 71:19]
  assign FullAdder_1191_io_a = io_pp_9[19]; // @[wallace.scala 69:18]
  assign FullAdder_1191_io_b = io_pp_10[18]; // @[wallace.scala 70:18]
  assign FullAdder_1191_io_ci = io_pp_11[17]; // @[wallace.scala 71:19]
  assign FullAdder_1192_io_a = io_pp_12[16]; // @[wallace.scala 69:18]
  assign FullAdder_1192_io_b = io_pp_13[15]; // @[wallace.scala 70:18]
  assign FullAdder_1192_io_ci = io_pp_14[14]; // @[wallace.scala 71:19]
  assign FullAdder_1193_io_a = io_pp_15[13]; // @[wallace.scala 69:18]
  assign FullAdder_1193_io_b = io_pp_16[12]; // @[wallace.scala 70:18]
  assign FullAdder_1193_io_ci = io_pp_17[11]; // @[wallace.scala 71:19]
  assign FullAdder_1194_io_a = io_pp_18[10]; // @[wallace.scala 69:18]
  assign FullAdder_1194_io_b = io_pp_19[9]; // @[wallace.scala 70:18]
  assign FullAdder_1194_io_ci = io_pp_20[8]; // @[wallace.scala 71:19]
  assign FullAdder_1195_io_a = io_pp_21[7]; // @[wallace.scala 69:18]
  assign FullAdder_1195_io_b = io_pp_22[6]; // @[wallace.scala 70:18]
  assign FullAdder_1195_io_ci = io_pp_23[5]; // @[wallace.scala 71:19]
  assign FullAdder_1196_io_a = io_pp_24[4]; // @[wallace.scala 69:18]
  assign FullAdder_1196_io_b = io_pp_25[3]; // @[wallace.scala 70:18]
  assign FullAdder_1196_io_ci = io_pp_26[2]; // @[wallace.scala 71:19]
  assign HalfAdder_25_io_a = io_pp_27[1]; // @[wallace.scala 59:18]
  assign HalfAdder_25_io_b = io_pp_28[0]; // @[wallace.scala 60:18]
  assign FullAdder_1197_io_a = io_pp_0[27]; // @[wallace.scala 69:18]
  assign FullAdder_1197_io_b = io_pp_1[26]; // @[wallace.scala 70:18]
  assign FullAdder_1197_io_ci = io_pp_2[25]; // @[wallace.scala 71:19]
  assign FullAdder_1198_io_a = io_pp_3[24]; // @[wallace.scala 69:18]
  assign FullAdder_1198_io_b = io_pp_4[23]; // @[wallace.scala 70:18]
  assign FullAdder_1198_io_ci = io_pp_5[22]; // @[wallace.scala 71:19]
  assign FullAdder_1199_io_a = io_pp_6[21]; // @[wallace.scala 69:18]
  assign FullAdder_1199_io_b = io_pp_7[20]; // @[wallace.scala 70:18]
  assign FullAdder_1199_io_ci = io_pp_8[19]; // @[wallace.scala 71:19]
  assign FullAdder_1200_io_a = io_pp_9[18]; // @[wallace.scala 69:18]
  assign FullAdder_1200_io_b = io_pp_10[17]; // @[wallace.scala 70:18]
  assign FullAdder_1200_io_ci = io_pp_11[16]; // @[wallace.scala 71:19]
  assign FullAdder_1201_io_a = io_pp_12[15]; // @[wallace.scala 69:18]
  assign FullAdder_1201_io_b = io_pp_13[14]; // @[wallace.scala 70:18]
  assign FullAdder_1201_io_ci = io_pp_14[13]; // @[wallace.scala 71:19]
  assign FullAdder_1202_io_a = io_pp_15[12]; // @[wallace.scala 69:18]
  assign FullAdder_1202_io_b = io_pp_16[11]; // @[wallace.scala 70:18]
  assign FullAdder_1202_io_ci = io_pp_17[10]; // @[wallace.scala 71:19]
  assign FullAdder_1203_io_a = io_pp_18[9]; // @[wallace.scala 69:18]
  assign FullAdder_1203_io_b = io_pp_19[8]; // @[wallace.scala 70:18]
  assign FullAdder_1203_io_ci = io_pp_20[7]; // @[wallace.scala 71:19]
  assign FullAdder_1204_io_a = io_pp_21[6]; // @[wallace.scala 69:18]
  assign FullAdder_1204_io_b = io_pp_22[5]; // @[wallace.scala 70:18]
  assign FullAdder_1204_io_ci = io_pp_23[4]; // @[wallace.scala 71:19]
  assign FullAdder_1205_io_a = io_pp_24[3]; // @[wallace.scala 69:18]
  assign FullAdder_1205_io_b = io_pp_25[2]; // @[wallace.scala 70:18]
  assign FullAdder_1205_io_ci = io_pp_26[1]; // @[wallace.scala 71:19]
  assign FullAdder_1206_io_a = io_pp_0[26]; // @[wallace.scala 69:18]
  assign FullAdder_1206_io_b = io_pp_1[25]; // @[wallace.scala 70:18]
  assign FullAdder_1206_io_ci = io_pp_2[24]; // @[wallace.scala 71:19]
  assign FullAdder_1207_io_a = io_pp_3[23]; // @[wallace.scala 69:18]
  assign FullAdder_1207_io_b = io_pp_4[22]; // @[wallace.scala 70:18]
  assign FullAdder_1207_io_ci = io_pp_5[21]; // @[wallace.scala 71:19]
  assign FullAdder_1208_io_a = io_pp_6[20]; // @[wallace.scala 69:18]
  assign FullAdder_1208_io_b = io_pp_7[19]; // @[wallace.scala 70:18]
  assign FullAdder_1208_io_ci = io_pp_8[18]; // @[wallace.scala 71:19]
  assign FullAdder_1209_io_a = io_pp_9[17]; // @[wallace.scala 69:18]
  assign FullAdder_1209_io_b = io_pp_10[16]; // @[wallace.scala 70:18]
  assign FullAdder_1209_io_ci = io_pp_11[15]; // @[wallace.scala 71:19]
  assign FullAdder_1210_io_a = io_pp_12[14]; // @[wallace.scala 69:18]
  assign FullAdder_1210_io_b = io_pp_13[13]; // @[wallace.scala 70:18]
  assign FullAdder_1210_io_ci = io_pp_14[12]; // @[wallace.scala 71:19]
  assign FullAdder_1211_io_a = io_pp_15[11]; // @[wallace.scala 69:18]
  assign FullAdder_1211_io_b = io_pp_16[10]; // @[wallace.scala 70:18]
  assign FullAdder_1211_io_ci = io_pp_17[9]; // @[wallace.scala 71:19]
  assign FullAdder_1212_io_a = io_pp_18[8]; // @[wallace.scala 69:18]
  assign FullAdder_1212_io_b = io_pp_19[7]; // @[wallace.scala 70:18]
  assign FullAdder_1212_io_ci = io_pp_20[6]; // @[wallace.scala 71:19]
  assign FullAdder_1213_io_a = io_pp_21[5]; // @[wallace.scala 69:18]
  assign FullAdder_1213_io_b = io_pp_22[4]; // @[wallace.scala 70:18]
  assign FullAdder_1213_io_ci = io_pp_23[3]; // @[wallace.scala 71:19]
  assign FullAdder_1214_io_a = io_pp_24[2]; // @[wallace.scala 69:18]
  assign FullAdder_1214_io_b = io_pp_25[1]; // @[wallace.scala 70:18]
  assign FullAdder_1214_io_ci = io_pp_26[0]; // @[wallace.scala 71:19]
  assign FullAdder_1215_io_a = io_pp_0[25]; // @[wallace.scala 69:18]
  assign FullAdder_1215_io_b = io_pp_1[24]; // @[wallace.scala 70:18]
  assign FullAdder_1215_io_ci = io_pp_2[23]; // @[wallace.scala 71:19]
  assign FullAdder_1216_io_a = io_pp_3[22]; // @[wallace.scala 69:18]
  assign FullAdder_1216_io_b = io_pp_4[21]; // @[wallace.scala 70:18]
  assign FullAdder_1216_io_ci = io_pp_5[20]; // @[wallace.scala 71:19]
  assign FullAdder_1217_io_a = io_pp_6[19]; // @[wallace.scala 69:18]
  assign FullAdder_1217_io_b = io_pp_7[18]; // @[wallace.scala 70:18]
  assign FullAdder_1217_io_ci = io_pp_8[17]; // @[wallace.scala 71:19]
  assign FullAdder_1218_io_a = io_pp_9[16]; // @[wallace.scala 69:18]
  assign FullAdder_1218_io_b = io_pp_10[15]; // @[wallace.scala 70:18]
  assign FullAdder_1218_io_ci = io_pp_11[14]; // @[wallace.scala 71:19]
  assign FullAdder_1219_io_a = io_pp_12[13]; // @[wallace.scala 69:18]
  assign FullAdder_1219_io_b = io_pp_13[12]; // @[wallace.scala 70:18]
  assign FullAdder_1219_io_ci = io_pp_14[11]; // @[wallace.scala 71:19]
  assign FullAdder_1220_io_a = io_pp_15[10]; // @[wallace.scala 69:18]
  assign FullAdder_1220_io_b = io_pp_16[9]; // @[wallace.scala 70:18]
  assign FullAdder_1220_io_ci = io_pp_17[8]; // @[wallace.scala 71:19]
  assign FullAdder_1221_io_a = io_pp_18[7]; // @[wallace.scala 69:18]
  assign FullAdder_1221_io_b = io_pp_19[6]; // @[wallace.scala 70:18]
  assign FullAdder_1221_io_ci = io_pp_20[5]; // @[wallace.scala 71:19]
  assign FullAdder_1222_io_a = io_pp_21[4]; // @[wallace.scala 69:18]
  assign FullAdder_1222_io_b = io_pp_22[3]; // @[wallace.scala 70:18]
  assign FullAdder_1222_io_ci = io_pp_23[2]; // @[wallace.scala 71:19]
  assign FullAdder_1223_io_a = io_pp_0[24]; // @[wallace.scala 69:18]
  assign FullAdder_1223_io_b = io_pp_1[23]; // @[wallace.scala 70:18]
  assign FullAdder_1223_io_ci = io_pp_2[22]; // @[wallace.scala 71:19]
  assign FullAdder_1224_io_a = io_pp_3[21]; // @[wallace.scala 69:18]
  assign FullAdder_1224_io_b = io_pp_4[20]; // @[wallace.scala 70:18]
  assign FullAdder_1224_io_ci = io_pp_5[19]; // @[wallace.scala 71:19]
  assign FullAdder_1225_io_a = io_pp_6[18]; // @[wallace.scala 69:18]
  assign FullAdder_1225_io_b = io_pp_7[17]; // @[wallace.scala 70:18]
  assign FullAdder_1225_io_ci = io_pp_8[16]; // @[wallace.scala 71:19]
  assign FullAdder_1226_io_a = io_pp_9[15]; // @[wallace.scala 69:18]
  assign FullAdder_1226_io_b = io_pp_10[14]; // @[wallace.scala 70:18]
  assign FullAdder_1226_io_ci = io_pp_11[13]; // @[wallace.scala 71:19]
  assign FullAdder_1227_io_a = io_pp_12[12]; // @[wallace.scala 69:18]
  assign FullAdder_1227_io_b = io_pp_13[11]; // @[wallace.scala 70:18]
  assign FullAdder_1227_io_ci = io_pp_14[10]; // @[wallace.scala 71:19]
  assign FullAdder_1228_io_a = io_pp_15[9]; // @[wallace.scala 69:18]
  assign FullAdder_1228_io_b = io_pp_16[8]; // @[wallace.scala 70:18]
  assign FullAdder_1228_io_ci = io_pp_17[7]; // @[wallace.scala 71:19]
  assign FullAdder_1229_io_a = io_pp_18[6]; // @[wallace.scala 69:18]
  assign FullAdder_1229_io_b = io_pp_19[5]; // @[wallace.scala 70:18]
  assign FullAdder_1229_io_ci = io_pp_20[4]; // @[wallace.scala 71:19]
  assign FullAdder_1230_io_a = io_pp_21[3]; // @[wallace.scala 69:18]
  assign FullAdder_1230_io_b = io_pp_22[2]; // @[wallace.scala 70:18]
  assign FullAdder_1230_io_ci = io_pp_23[1]; // @[wallace.scala 71:19]
  assign FullAdder_1231_io_a = io_pp_0[23]; // @[wallace.scala 69:18]
  assign FullAdder_1231_io_b = io_pp_1[22]; // @[wallace.scala 70:18]
  assign FullAdder_1231_io_ci = io_pp_2[21]; // @[wallace.scala 71:19]
  assign FullAdder_1232_io_a = io_pp_3[20]; // @[wallace.scala 69:18]
  assign FullAdder_1232_io_b = io_pp_4[19]; // @[wallace.scala 70:18]
  assign FullAdder_1232_io_ci = io_pp_5[18]; // @[wallace.scala 71:19]
  assign FullAdder_1233_io_a = io_pp_6[17]; // @[wallace.scala 69:18]
  assign FullAdder_1233_io_b = io_pp_7[16]; // @[wallace.scala 70:18]
  assign FullAdder_1233_io_ci = io_pp_8[15]; // @[wallace.scala 71:19]
  assign FullAdder_1234_io_a = io_pp_9[14]; // @[wallace.scala 69:18]
  assign FullAdder_1234_io_b = io_pp_10[13]; // @[wallace.scala 70:18]
  assign FullAdder_1234_io_ci = io_pp_11[12]; // @[wallace.scala 71:19]
  assign FullAdder_1235_io_a = io_pp_12[11]; // @[wallace.scala 69:18]
  assign FullAdder_1235_io_b = io_pp_13[10]; // @[wallace.scala 70:18]
  assign FullAdder_1235_io_ci = io_pp_14[9]; // @[wallace.scala 71:19]
  assign FullAdder_1236_io_a = io_pp_15[8]; // @[wallace.scala 69:18]
  assign FullAdder_1236_io_b = io_pp_16[7]; // @[wallace.scala 70:18]
  assign FullAdder_1236_io_ci = io_pp_17[6]; // @[wallace.scala 71:19]
  assign FullAdder_1237_io_a = io_pp_18[5]; // @[wallace.scala 69:18]
  assign FullAdder_1237_io_b = io_pp_19[4]; // @[wallace.scala 70:18]
  assign FullAdder_1237_io_ci = io_pp_20[3]; // @[wallace.scala 71:19]
  assign FullAdder_1238_io_a = io_pp_21[2]; // @[wallace.scala 69:18]
  assign FullAdder_1238_io_b = io_pp_22[1]; // @[wallace.scala 70:18]
  assign FullAdder_1238_io_ci = io_pp_23[0]; // @[wallace.scala 71:19]
  assign FullAdder_1239_io_a = io_pp_0[22]; // @[wallace.scala 69:18]
  assign FullAdder_1239_io_b = io_pp_1[21]; // @[wallace.scala 70:18]
  assign FullAdder_1239_io_ci = io_pp_2[20]; // @[wallace.scala 71:19]
  assign FullAdder_1240_io_a = io_pp_3[19]; // @[wallace.scala 69:18]
  assign FullAdder_1240_io_b = io_pp_4[18]; // @[wallace.scala 70:18]
  assign FullAdder_1240_io_ci = io_pp_5[17]; // @[wallace.scala 71:19]
  assign FullAdder_1241_io_a = io_pp_6[16]; // @[wallace.scala 69:18]
  assign FullAdder_1241_io_b = io_pp_7[15]; // @[wallace.scala 70:18]
  assign FullAdder_1241_io_ci = io_pp_8[14]; // @[wallace.scala 71:19]
  assign FullAdder_1242_io_a = io_pp_9[13]; // @[wallace.scala 69:18]
  assign FullAdder_1242_io_b = io_pp_10[12]; // @[wallace.scala 70:18]
  assign FullAdder_1242_io_ci = io_pp_11[11]; // @[wallace.scala 71:19]
  assign FullAdder_1243_io_a = io_pp_12[10]; // @[wallace.scala 69:18]
  assign FullAdder_1243_io_b = io_pp_13[9]; // @[wallace.scala 70:18]
  assign FullAdder_1243_io_ci = io_pp_14[8]; // @[wallace.scala 71:19]
  assign FullAdder_1244_io_a = io_pp_15[7]; // @[wallace.scala 69:18]
  assign FullAdder_1244_io_b = io_pp_16[6]; // @[wallace.scala 70:18]
  assign FullAdder_1244_io_ci = io_pp_17[5]; // @[wallace.scala 71:19]
  assign FullAdder_1245_io_a = io_pp_18[4]; // @[wallace.scala 69:18]
  assign FullAdder_1245_io_b = io_pp_19[3]; // @[wallace.scala 70:18]
  assign FullAdder_1245_io_ci = io_pp_20[2]; // @[wallace.scala 71:19]
  assign HalfAdder_26_io_a = io_pp_21[1]; // @[wallace.scala 59:18]
  assign HalfAdder_26_io_b = io_pp_22[0]; // @[wallace.scala 60:18]
  assign FullAdder_1246_io_a = io_pp_0[21]; // @[wallace.scala 69:18]
  assign FullAdder_1246_io_b = io_pp_1[20]; // @[wallace.scala 70:18]
  assign FullAdder_1246_io_ci = io_pp_2[19]; // @[wallace.scala 71:19]
  assign FullAdder_1247_io_a = io_pp_3[18]; // @[wallace.scala 69:18]
  assign FullAdder_1247_io_b = io_pp_4[17]; // @[wallace.scala 70:18]
  assign FullAdder_1247_io_ci = io_pp_5[16]; // @[wallace.scala 71:19]
  assign FullAdder_1248_io_a = io_pp_6[15]; // @[wallace.scala 69:18]
  assign FullAdder_1248_io_b = io_pp_7[14]; // @[wallace.scala 70:18]
  assign FullAdder_1248_io_ci = io_pp_8[13]; // @[wallace.scala 71:19]
  assign FullAdder_1249_io_a = io_pp_9[12]; // @[wallace.scala 69:18]
  assign FullAdder_1249_io_b = io_pp_10[11]; // @[wallace.scala 70:18]
  assign FullAdder_1249_io_ci = io_pp_11[10]; // @[wallace.scala 71:19]
  assign FullAdder_1250_io_a = io_pp_12[9]; // @[wallace.scala 69:18]
  assign FullAdder_1250_io_b = io_pp_13[8]; // @[wallace.scala 70:18]
  assign FullAdder_1250_io_ci = io_pp_14[7]; // @[wallace.scala 71:19]
  assign FullAdder_1251_io_a = io_pp_15[6]; // @[wallace.scala 69:18]
  assign FullAdder_1251_io_b = io_pp_16[5]; // @[wallace.scala 70:18]
  assign FullAdder_1251_io_ci = io_pp_17[4]; // @[wallace.scala 71:19]
  assign FullAdder_1252_io_a = io_pp_18[3]; // @[wallace.scala 69:18]
  assign FullAdder_1252_io_b = io_pp_19[2]; // @[wallace.scala 70:18]
  assign FullAdder_1252_io_ci = io_pp_20[1]; // @[wallace.scala 71:19]
  assign FullAdder_1253_io_a = io_pp_0[20]; // @[wallace.scala 69:18]
  assign FullAdder_1253_io_b = io_pp_1[19]; // @[wallace.scala 70:18]
  assign FullAdder_1253_io_ci = io_pp_2[18]; // @[wallace.scala 71:19]
  assign FullAdder_1254_io_a = io_pp_3[17]; // @[wallace.scala 69:18]
  assign FullAdder_1254_io_b = io_pp_4[16]; // @[wallace.scala 70:18]
  assign FullAdder_1254_io_ci = io_pp_5[15]; // @[wallace.scala 71:19]
  assign FullAdder_1255_io_a = io_pp_6[14]; // @[wallace.scala 69:18]
  assign FullAdder_1255_io_b = io_pp_7[13]; // @[wallace.scala 70:18]
  assign FullAdder_1255_io_ci = io_pp_8[12]; // @[wallace.scala 71:19]
  assign FullAdder_1256_io_a = io_pp_9[11]; // @[wallace.scala 69:18]
  assign FullAdder_1256_io_b = io_pp_10[10]; // @[wallace.scala 70:18]
  assign FullAdder_1256_io_ci = io_pp_11[9]; // @[wallace.scala 71:19]
  assign FullAdder_1257_io_a = io_pp_12[8]; // @[wallace.scala 69:18]
  assign FullAdder_1257_io_b = io_pp_13[7]; // @[wallace.scala 70:18]
  assign FullAdder_1257_io_ci = io_pp_14[6]; // @[wallace.scala 71:19]
  assign FullAdder_1258_io_a = io_pp_15[5]; // @[wallace.scala 69:18]
  assign FullAdder_1258_io_b = io_pp_16[4]; // @[wallace.scala 70:18]
  assign FullAdder_1258_io_ci = io_pp_17[3]; // @[wallace.scala 71:19]
  assign FullAdder_1259_io_a = io_pp_18[2]; // @[wallace.scala 69:18]
  assign FullAdder_1259_io_b = io_pp_19[1]; // @[wallace.scala 70:18]
  assign FullAdder_1259_io_ci = io_pp_20[0]; // @[wallace.scala 71:19]
  assign FullAdder_1260_io_a = io_pp_0[19]; // @[wallace.scala 69:18]
  assign FullAdder_1260_io_b = io_pp_1[18]; // @[wallace.scala 70:18]
  assign FullAdder_1260_io_ci = io_pp_2[17]; // @[wallace.scala 71:19]
  assign FullAdder_1261_io_a = io_pp_3[16]; // @[wallace.scala 69:18]
  assign FullAdder_1261_io_b = io_pp_4[15]; // @[wallace.scala 70:18]
  assign FullAdder_1261_io_ci = io_pp_5[14]; // @[wallace.scala 71:19]
  assign FullAdder_1262_io_a = io_pp_6[13]; // @[wallace.scala 69:18]
  assign FullAdder_1262_io_b = io_pp_7[12]; // @[wallace.scala 70:18]
  assign FullAdder_1262_io_ci = io_pp_8[11]; // @[wallace.scala 71:19]
  assign FullAdder_1263_io_a = io_pp_9[10]; // @[wallace.scala 69:18]
  assign FullAdder_1263_io_b = io_pp_10[9]; // @[wallace.scala 70:18]
  assign FullAdder_1263_io_ci = io_pp_11[8]; // @[wallace.scala 71:19]
  assign FullAdder_1264_io_a = io_pp_12[7]; // @[wallace.scala 69:18]
  assign FullAdder_1264_io_b = io_pp_13[6]; // @[wallace.scala 70:18]
  assign FullAdder_1264_io_ci = io_pp_14[5]; // @[wallace.scala 71:19]
  assign FullAdder_1265_io_a = io_pp_15[4]; // @[wallace.scala 69:18]
  assign FullAdder_1265_io_b = io_pp_16[3]; // @[wallace.scala 70:18]
  assign FullAdder_1265_io_ci = io_pp_17[2]; // @[wallace.scala 71:19]
  assign HalfAdder_27_io_a = io_pp_18[1]; // @[wallace.scala 59:18]
  assign HalfAdder_27_io_b = io_pp_19[0]; // @[wallace.scala 60:18]
  assign FullAdder_1266_io_a = io_pp_0[18]; // @[wallace.scala 69:18]
  assign FullAdder_1266_io_b = io_pp_1[17]; // @[wallace.scala 70:18]
  assign FullAdder_1266_io_ci = io_pp_2[16]; // @[wallace.scala 71:19]
  assign FullAdder_1267_io_a = io_pp_3[15]; // @[wallace.scala 69:18]
  assign FullAdder_1267_io_b = io_pp_4[14]; // @[wallace.scala 70:18]
  assign FullAdder_1267_io_ci = io_pp_5[13]; // @[wallace.scala 71:19]
  assign FullAdder_1268_io_a = io_pp_6[12]; // @[wallace.scala 69:18]
  assign FullAdder_1268_io_b = io_pp_7[11]; // @[wallace.scala 70:18]
  assign FullAdder_1268_io_ci = io_pp_8[10]; // @[wallace.scala 71:19]
  assign FullAdder_1269_io_a = io_pp_9[9]; // @[wallace.scala 69:18]
  assign FullAdder_1269_io_b = io_pp_10[8]; // @[wallace.scala 70:18]
  assign FullAdder_1269_io_ci = io_pp_11[7]; // @[wallace.scala 71:19]
  assign FullAdder_1270_io_a = io_pp_12[6]; // @[wallace.scala 69:18]
  assign FullAdder_1270_io_b = io_pp_13[5]; // @[wallace.scala 70:18]
  assign FullAdder_1270_io_ci = io_pp_14[4]; // @[wallace.scala 71:19]
  assign FullAdder_1271_io_a = io_pp_15[3]; // @[wallace.scala 69:18]
  assign FullAdder_1271_io_b = io_pp_16[2]; // @[wallace.scala 70:18]
  assign FullAdder_1271_io_ci = io_pp_17[1]; // @[wallace.scala 71:19]
  assign FullAdder_1272_io_a = io_pp_0[17]; // @[wallace.scala 69:18]
  assign FullAdder_1272_io_b = io_pp_1[16]; // @[wallace.scala 70:18]
  assign FullAdder_1272_io_ci = io_pp_2[15]; // @[wallace.scala 71:19]
  assign FullAdder_1273_io_a = io_pp_3[14]; // @[wallace.scala 69:18]
  assign FullAdder_1273_io_b = io_pp_4[13]; // @[wallace.scala 70:18]
  assign FullAdder_1273_io_ci = io_pp_5[12]; // @[wallace.scala 71:19]
  assign FullAdder_1274_io_a = io_pp_6[11]; // @[wallace.scala 69:18]
  assign FullAdder_1274_io_b = io_pp_7[10]; // @[wallace.scala 70:18]
  assign FullAdder_1274_io_ci = io_pp_8[9]; // @[wallace.scala 71:19]
  assign FullAdder_1275_io_a = io_pp_9[8]; // @[wallace.scala 69:18]
  assign FullAdder_1275_io_b = io_pp_10[7]; // @[wallace.scala 70:18]
  assign FullAdder_1275_io_ci = io_pp_11[6]; // @[wallace.scala 71:19]
  assign FullAdder_1276_io_a = io_pp_12[5]; // @[wallace.scala 69:18]
  assign FullAdder_1276_io_b = io_pp_13[4]; // @[wallace.scala 70:18]
  assign FullAdder_1276_io_ci = io_pp_14[3]; // @[wallace.scala 71:19]
  assign FullAdder_1277_io_a = io_pp_15[2]; // @[wallace.scala 69:18]
  assign FullAdder_1277_io_b = io_pp_16[1]; // @[wallace.scala 70:18]
  assign FullAdder_1277_io_ci = io_pp_17[0]; // @[wallace.scala 71:19]
  assign FullAdder_1278_io_a = io_pp_0[16]; // @[wallace.scala 69:18]
  assign FullAdder_1278_io_b = io_pp_1[15]; // @[wallace.scala 70:18]
  assign FullAdder_1278_io_ci = io_pp_2[14]; // @[wallace.scala 71:19]
  assign FullAdder_1279_io_a = io_pp_3[13]; // @[wallace.scala 69:18]
  assign FullAdder_1279_io_b = io_pp_4[12]; // @[wallace.scala 70:18]
  assign FullAdder_1279_io_ci = io_pp_5[11]; // @[wallace.scala 71:19]
  assign FullAdder_1280_io_a = io_pp_6[10]; // @[wallace.scala 69:18]
  assign FullAdder_1280_io_b = io_pp_7[9]; // @[wallace.scala 70:18]
  assign FullAdder_1280_io_ci = io_pp_8[8]; // @[wallace.scala 71:19]
  assign FullAdder_1281_io_a = io_pp_9[7]; // @[wallace.scala 69:18]
  assign FullAdder_1281_io_b = io_pp_10[6]; // @[wallace.scala 70:18]
  assign FullAdder_1281_io_ci = io_pp_11[5]; // @[wallace.scala 71:19]
  assign FullAdder_1282_io_a = io_pp_12[4]; // @[wallace.scala 69:18]
  assign FullAdder_1282_io_b = io_pp_13[3]; // @[wallace.scala 70:18]
  assign FullAdder_1282_io_ci = io_pp_14[2]; // @[wallace.scala 71:19]
  assign HalfAdder_28_io_a = io_pp_15[1]; // @[wallace.scala 59:18]
  assign HalfAdder_28_io_b = io_pp_16[0]; // @[wallace.scala 60:18]
  assign FullAdder_1283_io_a = io_pp_0[15]; // @[wallace.scala 69:18]
  assign FullAdder_1283_io_b = io_pp_1[14]; // @[wallace.scala 70:18]
  assign FullAdder_1283_io_ci = io_pp_2[13]; // @[wallace.scala 71:19]
  assign FullAdder_1284_io_a = io_pp_3[12]; // @[wallace.scala 69:18]
  assign FullAdder_1284_io_b = io_pp_4[11]; // @[wallace.scala 70:18]
  assign FullAdder_1284_io_ci = io_pp_5[10]; // @[wallace.scala 71:19]
  assign FullAdder_1285_io_a = io_pp_6[9]; // @[wallace.scala 69:18]
  assign FullAdder_1285_io_b = io_pp_7[8]; // @[wallace.scala 70:18]
  assign FullAdder_1285_io_ci = io_pp_8[7]; // @[wallace.scala 71:19]
  assign FullAdder_1286_io_a = io_pp_9[6]; // @[wallace.scala 69:18]
  assign FullAdder_1286_io_b = io_pp_10[5]; // @[wallace.scala 70:18]
  assign FullAdder_1286_io_ci = io_pp_11[4]; // @[wallace.scala 71:19]
  assign FullAdder_1287_io_a = io_pp_12[3]; // @[wallace.scala 69:18]
  assign FullAdder_1287_io_b = io_pp_13[2]; // @[wallace.scala 70:18]
  assign FullAdder_1287_io_ci = io_pp_14[1]; // @[wallace.scala 71:19]
  assign FullAdder_1288_io_a = io_pp_0[14]; // @[wallace.scala 69:18]
  assign FullAdder_1288_io_b = io_pp_1[13]; // @[wallace.scala 70:18]
  assign FullAdder_1288_io_ci = io_pp_2[12]; // @[wallace.scala 71:19]
  assign FullAdder_1289_io_a = io_pp_3[11]; // @[wallace.scala 69:18]
  assign FullAdder_1289_io_b = io_pp_4[10]; // @[wallace.scala 70:18]
  assign FullAdder_1289_io_ci = io_pp_5[9]; // @[wallace.scala 71:19]
  assign FullAdder_1290_io_a = io_pp_6[8]; // @[wallace.scala 69:18]
  assign FullAdder_1290_io_b = io_pp_7[7]; // @[wallace.scala 70:18]
  assign FullAdder_1290_io_ci = io_pp_8[6]; // @[wallace.scala 71:19]
  assign FullAdder_1291_io_a = io_pp_9[5]; // @[wallace.scala 69:18]
  assign FullAdder_1291_io_b = io_pp_10[4]; // @[wallace.scala 70:18]
  assign FullAdder_1291_io_ci = io_pp_11[3]; // @[wallace.scala 71:19]
  assign FullAdder_1292_io_a = io_pp_12[2]; // @[wallace.scala 69:18]
  assign FullAdder_1292_io_b = io_pp_13[1]; // @[wallace.scala 70:18]
  assign FullAdder_1292_io_ci = io_pp_14[0]; // @[wallace.scala 71:19]
  assign FullAdder_1293_io_a = io_pp_0[13]; // @[wallace.scala 69:18]
  assign FullAdder_1293_io_b = io_pp_1[12]; // @[wallace.scala 70:18]
  assign FullAdder_1293_io_ci = io_pp_2[11]; // @[wallace.scala 71:19]
  assign FullAdder_1294_io_a = io_pp_3[10]; // @[wallace.scala 69:18]
  assign FullAdder_1294_io_b = io_pp_4[9]; // @[wallace.scala 70:18]
  assign FullAdder_1294_io_ci = io_pp_5[8]; // @[wallace.scala 71:19]
  assign FullAdder_1295_io_a = io_pp_6[7]; // @[wallace.scala 69:18]
  assign FullAdder_1295_io_b = io_pp_7[6]; // @[wallace.scala 70:18]
  assign FullAdder_1295_io_ci = io_pp_8[5]; // @[wallace.scala 71:19]
  assign FullAdder_1296_io_a = io_pp_9[4]; // @[wallace.scala 69:18]
  assign FullAdder_1296_io_b = io_pp_10[3]; // @[wallace.scala 70:18]
  assign FullAdder_1296_io_ci = io_pp_11[2]; // @[wallace.scala 71:19]
  assign HalfAdder_29_io_a = io_pp_12[1]; // @[wallace.scala 59:18]
  assign HalfAdder_29_io_b = io_pp_13[0]; // @[wallace.scala 60:18]
  assign FullAdder_1297_io_a = io_pp_0[12]; // @[wallace.scala 69:18]
  assign FullAdder_1297_io_b = io_pp_1[11]; // @[wallace.scala 70:18]
  assign FullAdder_1297_io_ci = io_pp_2[10]; // @[wallace.scala 71:19]
  assign FullAdder_1298_io_a = io_pp_3[9]; // @[wallace.scala 69:18]
  assign FullAdder_1298_io_b = io_pp_4[8]; // @[wallace.scala 70:18]
  assign FullAdder_1298_io_ci = io_pp_5[7]; // @[wallace.scala 71:19]
  assign FullAdder_1299_io_a = io_pp_6[6]; // @[wallace.scala 69:18]
  assign FullAdder_1299_io_b = io_pp_7[5]; // @[wallace.scala 70:18]
  assign FullAdder_1299_io_ci = io_pp_8[4]; // @[wallace.scala 71:19]
  assign FullAdder_1300_io_a = io_pp_9[3]; // @[wallace.scala 69:18]
  assign FullAdder_1300_io_b = io_pp_10[2]; // @[wallace.scala 70:18]
  assign FullAdder_1300_io_ci = io_pp_11[1]; // @[wallace.scala 71:19]
  assign FullAdder_1301_io_a = io_pp_0[11]; // @[wallace.scala 69:18]
  assign FullAdder_1301_io_b = io_pp_1[10]; // @[wallace.scala 70:18]
  assign FullAdder_1301_io_ci = io_pp_2[9]; // @[wallace.scala 71:19]
  assign FullAdder_1302_io_a = io_pp_3[8]; // @[wallace.scala 69:18]
  assign FullAdder_1302_io_b = io_pp_4[7]; // @[wallace.scala 70:18]
  assign FullAdder_1302_io_ci = io_pp_5[6]; // @[wallace.scala 71:19]
  assign FullAdder_1303_io_a = io_pp_6[5]; // @[wallace.scala 69:18]
  assign FullAdder_1303_io_b = io_pp_7[4]; // @[wallace.scala 70:18]
  assign FullAdder_1303_io_ci = io_pp_8[3]; // @[wallace.scala 71:19]
  assign FullAdder_1304_io_a = io_pp_9[2]; // @[wallace.scala 69:18]
  assign FullAdder_1304_io_b = io_pp_10[1]; // @[wallace.scala 70:18]
  assign FullAdder_1304_io_ci = io_pp_11[0]; // @[wallace.scala 71:19]
  assign FullAdder_1305_io_a = io_pp_0[10]; // @[wallace.scala 69:18]
  assign FullAdder_1305_io_b = io_pp_1[9]; // @[wallace.scala 70:18]
  assign FullAdder_1305_io_ci = io_pp_2[8]; // @[wallace.scala 71:19]
  assign FullAdder_1306_io_a = io_pp_3[7]; // @[wallace.scala 69:18]
  assign FullAdder_1306_io_b = io_pp_4[6]; // @[wallace.scala 70:18]
  assign FullAdder_1306_io_ci = io_pp_5[5]; // @[wallace.scala 71:19]
  assign FullAdder_1307_io_a = io_pp_6[4]; // @[wallace.scala 69:18]
  assign FullAdder_1307_io_b = io_pp_7[3]; // @[wallace.scala 70:18]
  assign FullAdder_1307_io_ci = io_pp_8[2]; // @[wallace.scala 71:19]
  assign HalfAdder_30_io_a = io_pp_9[1]; // @[wallace.scala 59:18]
  assign HalfAdder_30_io_b = io_pp_10[0]; // @[wallace.scala 60:18]
  assign FullAdder_1308_io_a = io_pp_0[9]; // @[wallace.scala 69:18]
  assign FullAdder_1308_io_b = io_pp_1[8]; // @[wallace.scala 70:18]
  assign FullAdder_1308_io_ci = io_pp_2[7]; // @[wallace.scala 71:19]
  assign FullAdder_1309_io_a = io_pp_3[6]; // @[wallace.scala 69:18]
  assign FullAdder_1309_io_b = io_pp_4[5]; // @[wallace.scala 70:18]
  assign FullAdder_1309_io_ci = io_pp_5[4]; // @[wallace.scala 71:19]
  assign FullAdder_1310_io_a = io_pp_6[3]; // @[wallace.scala 69:18]
  assign FullAdder_1310_io_b = io_pp_7[2]; // @[wallace.scala 70:18]
  assign FullAdder_1310_io_ci = io_pp_8[1]; // @[wallace.scala 71:19]
  assign FullAdder_1311_io_a = io_pp_0[8]; // @[wallace.scala 69:18]
  assign FullAdder_1311_io_b = io_pp_1[7]; // @[wallace.scala 70:18]
  assign FullAdder_1311_io_ci = io_pp_2[6]; // @[wallace.scala 71:19]
  assign FullAdder_1312_io_a = io_pp_3[5]; // @[wallace.scala 69:18]
  assign FullAdder_1312_io_b = io_pp_4[4]; // @[wallace.scala 70:18]
  assign FullAdder_1312_io_ci = io_pp_5[3]; // @[wallace.scala 71:19]
  assign FullAdder_1313_io_a = io_pp_6[2]; // @[wallace.scala 69:18]
  assign FullAdder_1313_io_b = io_pp_7[1]; // @[wallace.scala 70:18]
  assign FullAdder_1313_io_ci = io_pp_8[0]; // @[wallace.scala 71:19]
  assign FullAdder_1314_io_a = io_pp_0[7]; // @[wallace.scala 69:18]
  assign FullAdder_1314_io_b = io_pp_1[6]; // @[wallace.scala 70:18]
  assign FullAdder_1314_io_ci = io_pp_2[5]; // @[wallace.scala 71:19]
  assign FullAdder_1315_io_a = io_pp_3[4]; // @[wallace.scala 69:18]
  assign FullAdder_1315_io_b = io_pp_4[3]; // @[wallace.scala 70:18]
  assign FullAdder_1315_io_ci = io_pp_5[2]; // @[wallace.scala 71:19]
  assign HalfAdder_31_io_a = io_pp_6[1]; // @[wallace.scala 59:18]
  assign HalfAdder_31_io_b = io_pp_7[0]; // @[wallace.scala 60:18]
  assign FullAdder_1316_io_a = io_pp_0[6]; // @[wallace.scala 69:18]
  assign FullAdder_1316_io_b = io_pp_1[5]; // @[wallace.scala 70:18]
  assign FullAdder_1316_io_ci = io_pp_2[4]; // @[wallace.scala 71:19]
  assign FullAdder_1317_io_a = io_pp_3[3]; // @[wallace.scala 69:18]
  assign FullAdder_1317_io_b = io_pp_4[2]; // @[wallace.scala 70:18]
  assign FullAdder_1317_io_ci = io_pp_5[1]; // @[wallace.scala 71:19]
  assign FullAdder_1318_io_a = io_pp_0[5]; // @[wallace.scala 69:18]
  assign FullAdder_1318_io_b = io_pp_1[4]; // @[wallace.scala 70:18]
  assign FullAdder_1318_io_ci = io_pp_2[3]; // @[wallace.scala 71:19]
  assign FullAdder_1319_io_a = io_pp_3[2]; // @[wallace.scala 69:18]
  assign FullAdder_1319_io_b = io_pp_4[1]; // @[wallace.scala 70:18]
  assign FullAdder_1319_io_ci = io_pp_5[0]; // @[wallace.scala 71:19]
  assign FullAdder_1320_io_a = io_pp_0[4]; // @[wallace.scala 69:18]
  assign FullAdder_1320_io_b = io_pp_1[3]; // @[wallace.scala 70:18]
  assign FullAdder_1320_io_ci = io_pp_2[2]; // @[wallace.scala 71:19]
  assign HalfAdder_32_io_a = io_pp_3[1]; // @[wallace.scala 59:18]
  assign HalfAdder_32_io_b = io_pp_4[0]; // @[wallace.scala 60:18]
  assign FullAdder_1321_io_a = io_pp_0[3]; // @[wallace.scala 69:18]
  assign FullAdder_1321_io_b = io_pp_1[2]; // @[wallace.scala 70:18]
  assign FullAdder_1321_io_ci = io_pp_2[1]; // @[wallace.scala 71:19]
  assign HalfAdder_33_io_a = io_pp_0[2]; // @[wallace.scala 59:18]
  assign HalfAdder_33_io_b = io_pp_1[1]; // @[wallace.scala 60:18]
  assign HalfAdder_34_io_a = io_pp_63[63]; // @[wallace.scala 59:18]
  assign HalfAdder_34_io_b = HalfAdder_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_35_io_a = HalfAdder_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_35_io_b = FullAdder_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_36_io_a = FullAdder_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_36_io_b = FullAdder_1_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1322_io_a = io_pp_63[60]; // @[wallace.scala 69:18]
  assign FullAdder_1322_io_b = FullAdder_1_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1322_io_ci = FullAdder_2_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1323_io_a = FullAdder_2_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1323_io_b = HalfAdder_1_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1323_io_ci = FullAdder_3_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1324_io_a = FullAdder_3_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1324_io_b = FullAdder_4_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1324_io_ci = FullAdder_5_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1325_io_a = io_pp_63[57]; // @[wallace.scala 69:18]
  assign FullAdder_1325_io_b = FullAdder_5_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1325_io_ci = FullAdder_6_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1326_io_a = FullAdder_7_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1326_io_b = FullAdder_8_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1326_io_ci = HalfAdder_2_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1327_io_a = FullAdder_7_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1327_io_b = FullAdder_8_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1327_io_ci = HalfAdder_2_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1328_io_a = FullAdder_9_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1328_io_b = FullAdder_10_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1328_io_ci = FullAdder_11_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1329_io_a = FullAdder_9_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1329_io_b = FullAdder_10_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1329_io_ci = FullAdder_11_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1330_io_a = FullAdder_12_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1330_io_b = FullAdder_13_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1330_io_ci = FullAdder_14_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1331_io_a = io_pp_63[54]; // @[wallace.scala 69:18]
  assign FullAdder_1331_io_b = FullAdder_12_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1331_io_ci = FullAdder_13_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1332_io_a = FullAdder_14_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1332_io_b = FullAdder_15_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1332_io_ci = FullAdder_16_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1333_io_a = FullAdder_15_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1333_io_b = FullAdder_16_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1333_io_ci = FullAdder_17_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1334_io_a = HalfAdder_3_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1334_io_b = FullAdder_18_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1334_io_ci = FullAdder_19_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_37_io_a = FullAdder_20_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_37_io_b = FullAdder_21_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1335_io_a = FullAdder_18_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1335_io_b = FullAdder_19_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1335_io_ci = FullAdder_20_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1336_io_a = FullAdder_21_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1336_io_b = FullAdder_22_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1336_io_ci = FullAdder_23_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_38_io_a = FullAdder_24_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_38_io_b = FullAdder_25_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1337_io_a = io_pp_63[51]; // @[wallace.scala 69:18]
  assign FullAdder_1337_io_b = FullAdder_22_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1337_io_ci = FullAdder_23_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1338_io_a = FullAdder_24_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1338_io_b = FullAdder_25_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1338_io_ci = FullAdder_26_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1339_io_a = FullAdder_27_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1339_io_b = FullAdder_28_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1339_io_ci = FullAdder_29_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1340_io_a = io_pp_62[51]; // @[wallace.scala 69:18]
  assign FullAdder_1340_io_b = io_pp_63[50]; // @[wallace.scala 70:18]
  assign FullAdder_1340_io_ci = FullAdder_26_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1341_io_a = FullAdder_27_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1341_io_b = FullAdder_28_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1341_io_ci = FullAdder_29_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1342_io_a = FullAdder_30_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1342_io_b = FullAdder_31_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1342_io_ci = FullAdder_32_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1343_io_a = FullAdder_30_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1343_io_b = FullAdder_31_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1343_io_ci = FullAdder_32_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1344_io_a = FullAdder_33_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1344_io_b = FullAdder_34_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1344_io_ci = FullAdder_35_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1345_io_a = FullAdder_36_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1345_io_b = FullAdder_37_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1345_io_ci = FullAdder_38_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1346_io_a = io_pp_63[48]; // @[wallace.scala 69:18]
  assign FullAdder_1346_io_b = FullAdder_35_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1346_io_ci = FullAdder_36_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1347_io_a = FullAdder_37_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1347_io_b = FullAdder_38_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1347_io_ci = FullAdder_39_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1348_io_a = FullAdder_40_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1348_io_b = FullAdder_41_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1348_io_ci = FullAdder_42_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1349_io_a = FullAdder_43_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1349_io_b = FullAdder_44_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1349_io_ci = HalfAdder_4_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1350_io_a = FullAdder_40_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1350_io_b = FullAdder_41_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1350_io_ci = FullAdder_42_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1351_io_a = FullAdder_43_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1351_io_b = FullAdder_44_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1351_io_ci = HalfAdder_4_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1352_io_a = FullAdder_45_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1352_io_b = FullAdder_46_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1352_io_ci = FullAdder_47_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1353_io_a = FullAdder_48_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1353_io_b = FullAdder_49_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1353_io_ci = FullAdder_50_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1354_io_a = FullAdder_45_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1354_io_b = FullAdder_46_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1354_io_ci = FullAdder_47_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1355_io_a = FullAdder_48_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1355_io_b = FullAdder_49_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1355_io_ci = FullAdder_50_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1356_io_a = FullAdder_51_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1356_io_b = FullAdder_52_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1356_io_ci = FullAdder_53_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1357_io_a = FullAdder_54_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1357_io_b = FullAdder_55_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1357_io_ci = FullAdder_56_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1358_io_a = io_pp_63[45]; // @[wallace.scala 69:18]
  assign FullAdder_1358_io_b = FullAdder_51_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1358_io_ci = FullAdder_52_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1359_io_a = FullAdder_53_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1359_io_b = FullAdder_54_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1359_io_ci = FullAdder_55_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1360_io_a = FullAdder_56_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1360_io_b = FullAdder_57_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1360_io_ci = FullAdder_58_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1361_io_a = FullAdder_59_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1361_io_b = FullAdder_60_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1361_io_ci = FullAdder_61_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_39_io_a = FullAdder_62_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_39_io_b = HalfAdder_5_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1362_io_a = FullAdder_57_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1362_io_b = FullAdder_58_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1362_io_ci = FullAdder_59_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1363_io_a = FullAdder_60_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1363_io_b = FullAdder_61_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1363_io_ci = FullAdder_62_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1364_io_a = HalfAdder_5_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1364_io_b = FullAdder_63_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1364_io_ci = FullAdder_64_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1365_io_a = FullAdder_65_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1365_io_b = FullAdder_66_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1365_io_ci = FullAdder_67_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_40_io_a = FullAdder_68_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_40_io_b = FullAdder_69_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1366_io_a = FullAdder_63_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1366_io_b = FullAdder_64_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1366_io_ci = FullAdder_65_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1367_io_a = FullAdder_66_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1367_io_b = FullAdder_67_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1367_io_ci = FullAdder_68_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1368_io_a = FullAdder_69_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1368_io_b = FullAdder_70_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1368_io_ci = FullAdder_71_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1369_io_a = FullAdder_72_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1369_io_b = FullAdder_73_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1369_io_ci = FullAdder_74_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_41_io_a = FullAdder_75_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_41_io_b = FullAdder_76_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1370_io_a = io_pp_63[42]; // @[wallace.scala 69:18]
  assign FullAdder_1370_io_b = FullAdder_70_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1370_io_ci = FullAdder_71_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1371_io_a = FullAdder_72_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1371_io_b = FullAdder_73_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1371_io_ci = FullAdder_74_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1372_io_a = FullAdder_75_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1372_io_b = FullAdder_76_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1372_io_ci = FullAdder_77_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1373_io_a = FullAdder_78_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1373_io_b = FullAdder_79_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1373_io_ci = FullAdder_80_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1374_io_a = FullAdder_81_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1374_io_b = FullAdder_82_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1374_io_ci = FullAdder_83_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1375_io_a = FullAdder_77_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1375_io_b = FullAdder_78_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1375_io_ci = FullAdder_79_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1376_io_a = FullAdder_80_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1376_io_b = FullAdder_81_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1376_io_ci = FullAdder_82_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1377_io_a = FullAdder_83_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1377_io_b = HalfAdder_6_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1377_io_ci = FullAdder_84_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1378_io_a = FullAdder_85_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1378_io_b = FullAdder_86_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1378_io_ci = FullAdder_87_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1379_io_a = FullAdder_88_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1379_io_b = FullAdder_89_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1379_io_ci = FullAdder_90_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1380_io_a = FullAdder_84_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1380_io_b = FullAdder_85_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1380_io_ci = FullAdder_86_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1381_io_a = FullAdder_87_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1381_io_b = FullAdder_88_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1381_io_ci = FullAdder_89_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1382_io_a = FullAdder_90_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1382_io_b = FullAdder_91_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1382_io_ci = FullAdder_92_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1383_io_a = FullAdder_93_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1383_io_b = FullAdder_94_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1383_io_ci = FullAdder_95_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1384_io_a = FullAdder_96_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1384_io_b = FullAdder_97_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1384_io_ci = FullAdder_98_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1385_io_a = io_pp_63[39]; // @[wallace.scala 69:18]
  assign FullAdder_1385_io_b = FullAdder_92_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1385_io_ci = FullAdder_93_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1386_io_a = FullAdder_94_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1386_io_b = FullAdder_95_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1386_io_ci = FullAdder_96_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1387_io_a = FullAdder_97_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1387_io_b = FullAdder_98_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1387_io_ci = FullAdder_99_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1388_io_a = FullAdder_100_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1388_io_b = FullAdder_101_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1388_io_ci = FullAdder_102_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1389_io_a = FullAdder_103_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1389_io_b = FullAdder_104_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1389_io_ci = FullAdder_105_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1390_io_a = io_pp_62[39]; // @[wallace.scala 69:18]
  assign FullAdder_1390_io_b = io_pp_63[38]; // @[wallace.scala 70:18]
  assign FullAdder_1390_io_ci = FullAdder_100_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1391_io_a = FullAdder_101_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1391_io_b = FullAdder_102_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1391_io_ci = FullAdder_103_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1392_io_a = FullAdder_104_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1392_io_b = FullAdder_105_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1392_io_ci = FullAdder_106_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1393_io_a = FullAdder_107_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1393_io_b = FullAdder_108_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1393_io_ci = FullAdder_109_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1394_io_a = FullAdder_110_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1394_io_b = FullAdder_111_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1394_io_ci = FullAdder_112_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1395_io_a = FullAdder_113_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1395_io_b = FullAdder_114_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1395_io_ci = FullAdder_115_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1396_io_a = FullAdder_108_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1396_io_b = FullAdder_109_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1396_io_ci = FullAdder_110_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1397_io_a = FullAdder_111_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1397_io_b = FullAdder_112_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1397_io_ci = FullAdder_113_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1398_io_a = FullAdder_114_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1398_io_b = FullAdder_115_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1398_io_ci = FullAdder_116_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1399_io_a = FullAdder_117_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1399_io_b = FullAdder_118_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1399_io_ci = FullAdder_119_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1400_io_a = FullAdder_120_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1400_io_b = FullAdder_121_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1400_io_ci = FullAdder_122_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1401_io_a = FullAdder_123_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1401_io_b = FullAdder_124_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1401_io_ci = FullAdder_125_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1402_io_a = io_pp_63[36]; // @[wallace.scala 69:18]
  assign FullAdder_1402_io_b = FullAdder_117_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1402_io_ci = FullAdder_118_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1403_io_a = FullAdder_119_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1403_io_b = FullAdder_120_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1403_io_ci = FullAdder_121_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1404_io_a = FullAdder_122_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1404_io_b = FullAdder_123_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1404_io_ci = FullAdder_124_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1405_io_a = FullAdder_125_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1405_io_b = FullAdder_126_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1405_io_ci = FullAdder_127_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1406_io_a = FullAdder_128_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1406_io_b = FullAdder_129_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1406_io_ci = FullAdder_130_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1407_io_a = FullAdder_131_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1407_io_b = FullAdder_132_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1407_io_ci = FullAdder_133_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1408_io_a = io_pp_62[36]; // @[wallace.scala 69:18]
  assign FullAdder_1408_io_b = io_pp_63[35]; // @[wallace.scala 70:18]
  assign FullAdder_1408_io_ci = FullAdder_126_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1409_io_a = FullAdder_127_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1409_io_b = FullAdder_128_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1409_io_ci = FullAdder_129_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1410_io_a = FullAdder_130_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1410_io_b = FullAdder_131_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1410_io_ci = FullAdder_132_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1411_io_a = FullAdder_133_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1411_io_b = FullAdder_134_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1411_io_ci = FullAdder_135_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1412_io_a = FullAdder_136_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1412_io_b = FullAdder_137_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1412_io_ci = FullAdder_138_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1413_io_a = FullAdder_139_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1413_io_b = FullAdder_140_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1413_io_ci = FullAdder_141_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1414_io_a = FullAdder_142_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1414_io_b = FullAdder_143_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1414_io_ci = FullAdder_144_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1415_io_a = FullAdder_135_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1415_io_b = FullAdder_136_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1415_io_ci = FullAdder_137_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1416_io_a = FullAdder_138_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1416_io_b = FullAdder_139_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1416_io_ci = FullAdder_140_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1417_io_a = FullAdder_141_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1417_io_b = FullAdder_142_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1417_io_ci = FullAdder_143_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1418_io_a = FullAdder_144_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1418_io_b = FullAdder_145_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1418_io_ci = FullAdder_146_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1419_io_a = FullAdder_147_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1419_io_b = FullAdder_148_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1419_io_ci = FullAdder_149_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1420_io_a = FullAdder_150_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1420_io_b = FullAdder_151_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1420_io_ci = FullAdder_152_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_42_io_a = FullAdder_153_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_42_io_b = FullAdder_154_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1421_io_a = io_pp_63[33]; // @[wallace.scala 69:18]
  assign FullAdder_1421_io_b = FullAdder_145_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1421_io_ci = FullAdder_146_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1422_io_a = FullAdder_147_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1422_io_b = FullAdder_148_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1422_io_ci = FullAdder_149_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1423_io_a = FullAdder_150_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1423_io_b = FullAdder_151_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1423_io_ci = FullAdder_152_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1424_io_a = FullAdder_153_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1424_io_b = FullAdder_154_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1424_io_ci = FullAdder_155_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1425_io_a = FullAdder_156_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1425_io_b = FullAdder_157_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1425_io_ci = FullAdder_158_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1426_io_a = FullAdder_159_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1426_io_b = FullAdder_160_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1426_io_ci = FullAdder_161_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1427_io_a = FullAdder_162_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1427_io_b = FullAdder_163_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1427_io_ci = FullAdder_164_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1428_io_a = FullAdder_155_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1428_io_b = FullAdder_156_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1428_io_ci = FullAdder_157_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1429_io_a = FullAdder_158_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1429_io_b = FullAdder_159_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1429_io_ci = FullAdder_160_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1430_io_a = FullAdder_161_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1430_io_b = FullAdder_162_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1430_io_ci = FullAdder_163_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1431_io_a = FullAdder_164_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1431_io_b = HalfAdder_7_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1431_io_ci = FullAdder_165_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1432_io_a = FullAdder_166_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1432_io_b = FullAdder_167_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1432_io_ci = FullAdder_168_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1433_io_a = FullAdder_169_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1433_io_b = FullAdder_170_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1433_io_ci = FullAdder_171_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1434_io_a = FullAdder_172_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1434_io_b = FullAdder_173_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1434_io_ci = FullAdder_174_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1435_io_a = FullAdder_165_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1435_io_b = FullAdder_166_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1435_io_ci = FullAdder_167_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1436_io_a = FullAdder_168_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1436_io_b = FullAdder_169_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1436_io_ci = FullAdder_170_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1437_io_a = FullAdder_171_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1437_io_b = FullAdder_172_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1437_io_ci = FullAdder_173_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1438_io_a = FullAdder_174_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1438_io_b = FullAdder_175_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1438_io_ci = FullAdder_176_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1439_io_a = FullAdder_177_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1439_io_b = FullAdder_178_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1439_io_ci = FullAdder_179_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1440_io_a = FullAdder_180_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1440_io_b = FullAdder_181_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1440_io_ci = FullAdder_182_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1441_io_a = FullAdder_183_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1441_io_b = FullAdder_184_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1441_io_ci = FullAdder_185_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1442_io_a = io_pp_63[30]; // @[wallace.scala 69:18]
  assign FullAdder_1442_io_b = FullAdder_176_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1442_io_ci = FullAdder_177_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1443_io_a = FullAdder_178_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1443_io_b = FullAdder_179_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1443_io_ci = FullAdder_180_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1444_io_a = FullAdder_181_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1444_io_b = FullAdder_182_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1444_io_ci = FullAdder_183_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1445_io_a = FullAdder_184_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1445_io_b = FullAdder_185_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1445_io_ci = FullAdder_186_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1446_io_a = FullAdder_187_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1446_io_b = FullAdder_188_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1446_io_ci = FullAdder_189_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1447_io_a = FullAdder_190_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1447_io_b = FullAdder_191_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1447_io_ci = FullAdder_192_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1448_io_a = FullAdder_193_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1448_io_b = FullAdder_194_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1448_io_ci = FullAdder_195_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1449_io_a = FullAdder_196_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1449_io_b = FullAdder_197_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1449_io_ci = HalfAdder_8_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1450_io_a = FullAdder_187_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1450_io_b = FullAdder_188_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1450_io_ci = FullAdder_189_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1451_io_a = FullAdder_190_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1451_io_b = FullAdder_191_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1451_io_ci = FullAdder_192_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1452_io_a = FullAdder_193_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1452_io_b = FullAdder_194_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1452_io_ci = FullAdder_195_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1453_io_a = FullAdder_196_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1453_io_b = FullAdder_197_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1453_io_ci = HalfAdder_8_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1454_io_a = FullAdder_198_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1454_io_b = FullAdder_199_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1454_io_ci = FullAdder_200_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1455_io_a = FullAdder_201_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1455_io_b = FullAdder_202_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1455_io_ci = FullAdder_203_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1456_io_a = FullAdder_204_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1456_io_b = FullAdder_205_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1456_io_ci = FullAdder_206_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1457_io_a = FullAdder_207_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1457_io_b = FullAdder_208_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1457_io_ci = FullAdder_209_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1458_io_a = FullAdder_198_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1458_io_b = FullAdder_199_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1458_io_ci = FullAdder_200_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1459_io_a = FullAdder_201_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1459_io_b = FullAdder_202_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1459_io_ci = FullAdder_203_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1460_io_a = FullAdder_204_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1460_io_b = FullAdder_205_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1460_io_ci = FullAdder_206_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1461_io_a = FullAdder_207_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1461_io_b = FullAdder_208_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1461_io_ci = FullAdder_209_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1462_io_a = FullAdder_210_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1462_io_b = FullAdder_211_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1462_io_ci = FullAdder_212_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1463_io_a = FullAdder_213_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1463_io_b = FullAdder_214_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1463_io_ci = FullAdder_215_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1464_io_a = FullAdder_216_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1464_io_b = FullAdder_217_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1464_io_ci = FullAdder_218_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1465_io_a = FullAdder_219_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1465_io_b = FullAdder_220_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1465_io_ci = FullAdder_221_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1466_io_a = io_pp_63[27]; // @[wallace.scala 69:18]
  assign FullAdder_1466_io_b = FullAdder_210_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1466_io_ci = FullAdder_211_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1467_io_a = FullAdder_212_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1467_io_b = FullAdder_213_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1467_io_ci = FullAdder_214_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1468_io_a = FullAdder_215_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1468_io_b = FullAdder_216_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1468_io_ci = FullAdder_217_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1469_io_a = FullAdder_218_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1469_io_b = FullAdder_219_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1469_io_ci = FullAdder_220_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1470_io_a = FullAdder_221_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1470_io_b = FullAdder_222_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1470_io_ci = FullAdder_223_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1471_io_a = FullAdder_224_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1471_io_b = FullAdder_225_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1471_io_ci = FullAdder_226_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1472_io_a = FullAdder_227_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1472_io_b = FullAdder_228_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1472_io_ci = FullAdder_229_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1473_io_a = FullAdder_230_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1473_io_b = FullAdder_231_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1473_io_ci = FullAdder_232_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_43_io_a = FullAdder_233_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_43_io_b = HalfAdder_9_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1474_io_a = FullAdder_222_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1474_io_b = FullAdder_223_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1474_io_ci = FullAdder_224_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1475_io_a = FullAdder_225_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1475_io_b = FullAdder_226_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1475_io_ci = FullAdder_227_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1476_io_a = FullAdder_228_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1476_io_b = FullAdder_229_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1476_io_ci = FullAdder_230_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1477_io_a = FullAdder_231_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1477_io_b = FullAdder_232_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1477_io_ci = FullAdder_233_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1478_io_a = HalfAdder_9_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1478_io_b = FullAdder_234_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1478_io_ci = FullAdder_235_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1479_io_a = FullAdder_236_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1479_io_b = FullAdder_237_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1479_io_ci = FullAdder_238_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1480_io_a = FullAdder_239_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1480_io_b = FullAdder_240_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1480_io_ci = FullAdder_241_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1481_io_a = FullAdder_242_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1481_io_b = FullAdder_243_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1481_io_ci = FullAdder_244_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_44_io_a = FullAdder_245_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_44_io_b = FullAdder_246_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1482_io_a = FullAdder_234_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1482_io_b = FullAdder_235_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1482_io_ci = FullAdder_236_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1483_io_a = FullAdder_237_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1483_io_b = FullAdder_238_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1483_io_ci = FullAdder_239_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1484_io_a = FullAdder_240_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1484_io_b = FullAdder_241_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1484_io_ci = FullAdder_242_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1485_io_a = FullAdder_243_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1485_io_b = FullAdder_244_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1485_io_ci = FullAdder_245_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1486_io_a = FullAdder_246_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1486_io_b = FullAdder_247_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1486_io_ci = FullAdder_248_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1487_io_a = FullAdder_249_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1487_io_b = FullAdder_250_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1487_io_ci = FullAdder_251_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1488_io_a = FullAdder_252_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1488_io_b = FullAdder_253_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1488_io_ci = FullAdder_254_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1489_io_a = FullAdder_255_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1489_io_b = FullAdder_256_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1489_io_ci = FullAdder_257_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_45_io_a = FullAdder_258_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_45_io_b = FullAdder_259_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1490_io_a = io_pp_63[24]; // @[wallace.scala 69:18]
  assign FullAdder_1490_io_b = FullAdder_247_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1490_io_ci = FullAdder_248_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1491_io_a = FullAdder_249_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1491_io_b = FullAdder_250_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1491_io_ci = FullAdder_251_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1492_io_a = FullAdder_252_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1492_io_b = FullAdder_253_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1492_io_ci = FullAdder_254_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1493_io_a = FullAdder_255_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1493_io_b = FullAdder_256_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1493_io_ci = FullAdder_257_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1494_io_a = FullAdder_258_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1494_io_b = FullAdder_259_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1494_io_ci = FullAdder_260_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1495_io_a = FullAdder_261_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1495_io_b = FullAdder_262_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1495_io_ci = FullAdder_263_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1496_io_a = FullAdder_264_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1496_io_b = FullAdder_265_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1496_io_ci = FullAdder_266_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1497_io_a = FullAdder_267_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1497_io_b = FullAdder_268_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1497_io_ci = FullAdder_269_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1498_io_a = FullAdder_270_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1498_io_b = FullAdder_271_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1498_io_ci = FullAdder_272_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1499_io_a = FullAdder_260_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1499_io_b = FullAdder_261_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1499_io_ci = FullAdder_262_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1500_io_a = FullAdder_263_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1500_io_b = FullAdder_264_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1500_io_ci = FullAdder_265_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1501_io_a = FullAdder_266_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1501_io_b = FullAdder_267_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1501_io_ci = FullAdder_268_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1502_io_a = FullAdder_269_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1502_io_b = FullAdder_270_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1502_io_ci = FullAdder_271_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1503_io_a = FullAdder_272_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1503_io_b = HalfAdder_10_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1503_io_ci = FullAdder_273_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1504_io_a = FullAdder_274_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1504_io_b = FullAdder_275_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1504_io_ci = FullAdder_276_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1505_io_a = FullAdder_277_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1505_io_b = FullAdder_278_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1505_io_ci = FullAdder_279_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1506_io_a = FullAdder_280_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1506_io_b = FullAdder_281_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1506_io_ci = FullAdder_282_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1507_io_a = FullAdder_283_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1507_io_b = FullAdder_284_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1507_io_ci = FullAdder_285_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1508_io_a = FullAdder_273_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1508_io_b = FullAdder_274_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1508_io_ci = FullAdder_275_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1509_io_a = FullAdder_276_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1509_io_b = FullAdder_277_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1509_io_ci = FullAdder_278_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1510_io_a = FullAdder_279_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1510_io_b = FullAdder_280_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1510_io_ci = FullAdder_281_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1511_io_a = FullAdder_282_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1511_io_b = FullAdder_283_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1511_io_ci = FullAdder_284_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1512_io_a = FullAdder_285_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1512_io_b = FullAdder_286_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1512_io_ci = FullAdder_287_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1513_io_a = FullAdder_288_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1513_io_b = FullAdder_289_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1513_io_ci = FullAdder_290_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1514_io_a = FullAdder_291_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1514_io_b = FullAdder_292_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1514_io_ci = FullAdder_293_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1515_io_a = FullAdder_294_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1515_io_b = FullAdder_295_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1515_io_ci = FullAdder_296_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1516_io_a = FullAdder_297_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1516_io_b = FullAdder_298_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1516_io_ci = FullAdder_299_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1517_io_a = io_pp_63[21]; // @[wallace.scala 69:18]
  assign FullAdder_1517_io_b = FullAdder_287_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1517_io_ci = FullAdder_288_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1518_io_a = FullAdder_289_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1518_io_b = FullAdder_290_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1518_io_ci = FullAdder_291_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1519_io_a = FullAdder_292_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1519_io_b = FullAdder_293_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1519_io_ci = FullAdder_294_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1520_io_a = FullAdder_295_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1520_io_b = FullAdder_296_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1520_io_ci = FullAdder_297_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1521_io_a = FullAdder_298_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1521_io_b = FullAdder_299_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1521_io_ci = FullAdder_300_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1522_io_a = FullAdder_301_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1522_io_b = FullAdder_302_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1522_io_ci = FullAdder_303_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1523_io_a = FullAdder_304_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1523_io_b = FullAdder_305_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1523_io_ci = FullAdder_306_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1524_io_a = FullAdder_307_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1524_io_b = FullAdder_308_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1524_io_ci = FullAdder_309_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1525_io_a = FullAdder_310_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1525_io_b = FullAdder_311_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1525_io_ci = FullAdder_312_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1526_io_a = FullAdder_313_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1526_io_b = FullAdder_314_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1526_io_ci = HalfAdder_11_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1527_io_a = FullAdder_301_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1527_io_b = FullAdder_302_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1527_io_ci = FullAdder_303_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1528_io_a = FullAdder_304_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1528_io_b = FullAdder_305_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1528_io_ci = FullAdder_306_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1529_io_a = FullAdder_307_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1529_io_b = FullAdder_308_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1529_io_ci = FullAdder_309_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1530_io_a = FullAdder_310_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1530_io_b = FullAdder_311_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1530_io_ci = FullAdder_312_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1531_io_a = FullAdder_313_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1531_io_b = FullAdder_314_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1531_io_ci = HalfAdder_11_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1532_io_a = FullAdder_315_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1532_io_b = FullAdder_316_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1532_io_ci = FullAdder_317_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1533_io_a = FullAdder_318_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1533_io_b = FullAdder_319_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1533_io_ci = FullAdder_320_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1534_io_a = FullAdder_321_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1534_io_b = FullAdder_322_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1534_io_ci = FullAdder_323_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1535_io_a = FullAdder_324_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1535_io_b = FullAdder_325_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1535_io_ci = FullAdder_326_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1536_io_a = FullAdder_327_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1536_io_b = FullAdder_328_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1536_io_ci = FullAdder_329_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1537_io_a = FullAdder_315_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1537_io_b = FullAdder_316_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1537_io_ci = FullAdder_317_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1538_io_a = FullAdder_318_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1538_io_b = FullAdder_319_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1538_io_ci = FullAdder_320_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1539_io_a = FullAdder_321_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1539_io_b = FullAdder_322_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1539_io_ci = FullAdder_323_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1540_io_a = FullAdder_324_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1540_io_b = FullAdder_325_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1540_io_ci = FullAdder_326_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1541_io_a = FullAdder_327_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1541_io_b = FullAdder_328_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1541_io_ci = FullAdder_329_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1542_io_a = FullAdder_330_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1542_io_b = FullAdder_331_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1542_io_ci = FullAdder_332_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1543_io_a = FullAdder_333_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1543_io_b = FullAdder_334_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1543_io_ci = FullAdder_335_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1544_io_a = FullAdder_336_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1544_io_b = FullAdder_337_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1544_io_ci = FullAdder_338_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1545_io_a = FullAdder_339_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1545_io_b = FullAdder_340_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1545_io_ci = FullAdder_341_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1546_io_a = FullAdder_342_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1546_io_b = FullAdder_343_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1546_io_ci = FullAdder_344_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1547_io_a = io_pp_63[18]; // @[wallace.scala 69:18]
  assign FullAdder_1547_io_b = FullAdder_330_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1547_io_ci = FullAdder_331_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1548_io_a = FullAdder_332_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1548_io_b = FullAdder_333_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1548_io_ci = FullAdder_334_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1549_io_a = FullAdder_335_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1549_io_b = FullAdder_336_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1549_io_ci = FullAdder_337_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1550_io_a = FullAdder_338_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1550_io_b = FullAdder_339_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1550_io_ci = FullAdder_340_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1551_io_a = FullAdder_341_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1551_io_b = FullAdder_342_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1551_io_ci = FullAdder_343_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1552_io_a = FullAdder_344_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1552_io_b = FullAdder_345_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1552_io_ci = FullAdder_346_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1553_io_a = FullAdder_347_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1553_io_b = FullAdder_348_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1553_io_ci = FullAdder_349_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1554_io_a = FullAdder_350_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1554_io_b = FullAdder_351_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1554_io_ci = FullAdder_352_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1555_io_a = FullAdder_353_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1555_io_b = FullAdder_354_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1555_io_ci = FullAdder_355_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1556_io_a = FullAdder_356_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1556_io_b = FullAdder_357_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1556_io_ci = FullAdder_358_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1557_io_a = FullAdder_345_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1557_io_b = FullAdder_346_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1557_io_ci = FullAdder_347_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1558_io_a = FullAdder_348_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1558_io_b = FullAdder_349_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1558_io_ci = FullAdder_350_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1559_io_a = FullAdder_351_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1559_io_b = FullAdder_352_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1559_io_ci = FullAdder_353_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1560_io_a = FullAdder_354_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1560_io_b = FullAdder_355_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1560_io_ci = FullAdder_356_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1561_io_a = FullAdder_357_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1561_io_b = FullAdder_358_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1561_io_ci = FullAdder_359_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1562_io_a = HalfAdder_12_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1562_io_b = FullAdder_360_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1562_io_ci = FullAdder_361_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1563_io_a = FullAdder_362_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1563_io_b = FullAdder_363_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1563_io_ci = FullAdder_364_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1564_io_a = FullAdder_365_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1564_io_b = FullAdder_366_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1564_io_ci = FullAdder_367_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1565_io_a = FullAdder_368_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1565_io_b = FullAdder_369_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1565_io_ci = FullAdder_370_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1566_io_a = FullAdder_371_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1566_io_b = FullAdder_372_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1566_io_ci = FullAdder_373_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1567_io_a = FullAdder_360_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1567_io_b = FullAdder_361_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1567_io_ci = FullAdder_362_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1568_io_a = FullAdder_363_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1568_io_b = FullAdder_364_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1568_io_ci = FullAdder_365_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1569_io_a = FullAdder_366_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1569_io_b = FullAdder_367_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1569_io_ci = FullAdder_368_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1570_io_a = FullAdder_369_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1570_io_b = FullAdder_370_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1570_io_ci = FullAdder_371_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1571_io_a = FullAdder_372_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1571_io_b = FullAdder_373_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1571_io_ci = FullAdder_374_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1572_io_a = FullAdder_375_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1572_io_b = FullAdder_376_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1572_io_ci = FullAdder_377_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1573_io_a = FullAdder_378_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1573_io_b = FullAdder_379_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1573_io_ci = FullAdder_380_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1574_io_a = FullAdder_381_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1574_io_b = FullAdder_382_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1574_io_ci = FullAdder_383_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1575_io_a = FullAdder_384_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1575_io_b = FullAdder_385_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1575_io_ci = FullAdder_386_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1576_io_a = FullAdder_387_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1576_io_b = FullAdder_388_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1576_io_ci = FullAdder_389_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_46_io_a = FullAdder_390_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_46_io_b = FullAdder_391_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1577_io_a = io_pp_63[15]; // @[wallace.scala 69:18]
  assign FullAdder_1577_io_b = FullAdder_376_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1577_io_ci = FullAdder_377_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1578_io_a = FullAdder_378_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1578_io_b = FullAdder_379_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1578_io_ci = FullAdder_380_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1579_io_a = FullAdder_381_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1579_io_b = FullAdder_382_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1579_io_ci = FullAdder_383_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1580_io_a = FullAdder_384_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1580_io_b = FullAdder_385_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1580_io_ci = FullAdder_386_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1581_io_a = FullAdder_387_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1581_io_b = FullAdder_388_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1581_io_ci = FullAdder_389_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1582_io_a = FullAdder_390_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1582_io_b = FullAdder_391_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1582_io_ci = FullAdder_392_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1583_io_a = FullAdder_393_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1583_io_b = FullAdder_394_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1583_io_ci = FullAdder_395_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1584_io_a = FullAdder_396_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1584_io_b = FullAdder_397_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1584_io_ci = FullAdder_398_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1585_io_a = FullAdder_399_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1585_io_b = FullAdder_400_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1585_io_ci = FullAdder_401_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1586_io_a = FullAdder_402_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1586_io_b = FullAdder_403_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1586_io_ci = FullAdder_404_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1587_io_a = FullAdder_405_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1587_io_b = FullAdder_406_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1587_io_ci = FullAdder_407_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1588_io_a = FullAdder_392_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1588_io_b = FullAdder_393_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1588_io_ci = FullAdder_394_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1589_io_a = FullAdder_395_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1589_io_b = FullAdder_396_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1589_io_ci = FullAdder_397_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1590_io_a = FullAdder_398_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1590_io_b = FullAdder_399_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1590_io_ci = FullAdder_400_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1591_io_a = FullAdder_401_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1591_io_b = FullAdder_402_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1591_io_ci = FullAdder_403_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1592_io_a = FullAdder_404_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1592_io_b = FullAdder_405_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1592_io_ci = FullAdder_406_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1593_io_a = FullAdder_407_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1593_io_b = HalfAdder_13_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1593_io_ci = FullAdder_408_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1594_io_a = FullAdder_409_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1594_io_b = FullAdder_410_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1594_io_ci = FullAdder_411_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1595_io_a = FullAdder_412_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1595_io_b = FullAdder_413_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1595_io_ci = FullAdder_414_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1596_io_a = FullAdder_415_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1596_io_b = FullAdder_416_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1596_io_ci = FullAdder_417_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1597_io_a = FullAdder_418_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1597_io_b = FullAdder_419_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1597_io_ci = FullAdder_420_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1598_io_a = FullAdder_421_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1598_io_b = FullAdder_422_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1598_io_ci = FullAdder_423_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1599_io_a = FullAdder_408_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1599_io_b = FullAdder_409_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1599_io_ci = FullAdder_410_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1600_io_a = FullAdder_411_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1600_io_b = FullAdder_412_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1600_io_ci = FullAdder_413_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1601_io_a = FullAdder_414_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1601_io_b = FullAdder_415_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1601_io_ci = FullAdder_416_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1602_io_a = FullAdder_417_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1602_io_b = FullAdder_418_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1602_io_ci = FullAdder_419_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1603_io_a = FullAdder_420_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1603_io_b = FullAdder_421_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1603_io_ci = FullAdder_422_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1604_io_a = FullAdder_423_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1604_io_b = FullAdder_424_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1604_io_ci = FullAdder_425_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1605_io_a = FullAdder_426_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1605_io_b = FullAdder_427_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1605_io_ci = FullAdder_428_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1606_io_a = FullAdder_429_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1606_io_b = FullAdder_430_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1606_io_ci = FullAdder_431_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1607_io_a = FullAdder_432_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1607_io_b = FullAdder_433_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1607_io_ci = FullAdder_434_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1608_io_a = FullAdder_435_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1608_io_b = FullAdder_436_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1608_io_ci = FullAdder_437_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1609_io_a = FullAdder_438_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1609_io_b = FullAdder_439_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1609_io_ci = FullAdder_440_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1610_io_a = io_pp_63[12]; // @[wallace.scala 69:18]
  assign FullAdder_1610_io_b = FullAdder_425_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1610_io_ci = FullAdder_426_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1611_io_a = FullAdder_427_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1611_io_b = FullAdder_428_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1611_io_ci = FullAdder_429_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1612_io_a = FullAdder_430_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1612_io_b = FullAdder_431_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1612_io_ci = FullAdder_432_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1613_io_a = FullAdder_433_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1613_io_b = FullAdder_434_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1613_io_ci = FullAdder_435_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1614_io_a = FullAdder_436_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1614_io_b = FullAdder_437_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1614_io_ci = FullAdder_438_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1615_io_a = FullAdder_439_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1615_io_b = FullAdder_440_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1615_io_ci = FullAdder_441_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1616_io_a = FullAdder_442_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1616_io_b = FullAdder_443_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1616_io_ci = FullAdder_444_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1617_io_a = FullAdder_445_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1617_io_b = FullAdder_446_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1617_io_ci = FullAdder_447_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1618_io_a = FullAdder_448_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1618_io_b = FullAdder_449_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1618_io_ci = FullAdder_450_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1619_io_a = FullAdder_451_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1619_io_b = FullAdder_452_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1619_io_ci = FullAdder_453_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1620_io_a = FullAdder_454_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1620_io_b = FullAdder_455_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1620_io_ci = FullAdder_456_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1621_io_a = FullAdder_457_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1621_io_b = FullAdder_458_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1621_io_ci = HalfAdder_14_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1622_io_a = FullAdder_442_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1622_io_b = FullAdder_443_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1622_io_ci = FullAdder_444_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1623_io_a = FullAdder_445_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1623_io_b = FullAdder_446_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1623_io_ci = FullAdder_447_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1624_io_a = FullAdder_448_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1624_io_b = FullAdder_449_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1624_io_ci = FullAdder_450_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1625_io_a = FullAdder_451_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1625_io_b = FullAdder_452_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1625_io_ci = FullAdder_453_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1626_io_a = FullAdder_454_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1626_io_b = FullAdder_455_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1626_io_ci = FullAdder_456_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1627_io_a = FullAdder_457_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1627_io_b = FullAdder_458_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1627_io_ci = HalfAdder_14_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1628_io_a = FullAdder_459_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1628_io_b = FullAdder_460_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1628_io_ci = FullAdder_461_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1629_io_a = FullAdder_462_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1629_io_b = FullAdder_463_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1629_io_ci = FullAdder_464_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1630_io_a = FullAdder_465_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1630_io_b = FullAdder_466_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1630_io_ci = FullAdder_467_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1631_io_a = FullAdder_468_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1631_io_b = FullAdder_469_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1631_io_ci = FullAdder_470_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1632_io_a = FullAdder_471_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1632_io_b = FullAdder_472_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1632_io_ci = FullAdder_473_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1633_io_a = FullAdder_474_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1633_io_b = FullAdder_475_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1633_io_ci = FullAdder_476_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1634_io_a = FullAdder_459_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1634_io_b = FullAdder_460_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1634_io_ci = FullAdder_461_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1635_io_a = FullAdder_462_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1635_io_b = FullAdder_463_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1635_io_ci = FullAdder_464_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1636_io_a = FullAdder_465_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1636_io_b = FullAdder_466_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1636_io_ci = FullAdder_467_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1637_io_a = FullAdder_468_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1637_io_b = FullAdder_469_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1637_io_ci = FullAdder_470_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1638_io_a = FullAdder_471_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1638_io_b = FullAdder_472_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1638_io_ci = FullAdder_473_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1639_io_a = FullAdder_474_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1639_io_b = FullAdder_475_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1639_io_ci = FullAdder_476_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1640_io_a = FullAdder_477_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1640_io_b = FullAdder_478_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1640_io_ci = FullAdder_479_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1641_io_a = FullAdder_480_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1641_io_b = FullAdder_481_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1641_io_ci = FullAdder_482_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1642_io_a = FullAdder_483_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1642_io_b = FullAdder_484_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1642_io_ci = FullAdder_485_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1643_io_a = FullAdder_486_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1643_io_b = FullAdder_487_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1643_io_ci = FullAdder_488_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1644_io_a = FullAdder_489_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1644_io_b = FullAdder_490_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1644_io_ci = FullAdder_491_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1645_io_a = FullAdder_492_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1645_io_b = FullAdder_493_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1645_io_ci = FullAdder_494_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1646_io_a = io_pp_63[9]; // @[wallace.scala 69:18]
  assign FullAdder_1646_io_b = FullAdder_477_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1646_io_ci = FullAdder_478_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1647_io_a = FullAdder_479_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1647_io_b = FullAdder_480_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1647_io_ci = FullAdder_481_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1648_io_a = FullAdder_482_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1648_io_b = FullAdder_483_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1648_io_ci = FullAdder_484_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1649_io_a = FullAdder_485_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1649_io_b = FullAdder_486_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1649_io_ci = FullAdder_487_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1650_io_a = FullAdder_488_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1650_io_b = FullAdder_489_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1650_io_ci = FullAdder_490_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1651_io_a = FullAdder_491_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1651_io_b = FullAdder_492_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1651_io_ci = FullAdder_493_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1652_io_a = FullAdder_494_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1652_io_b = FullAdder_495_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1652_io_ci = FullAdder_496_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1653_io_a = FullAdder_497_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1653_io_b = FullAdder_498_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1653_io_ci = FullAdder_499_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1654_io_a = FullAdder_500_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1654_io_b = FullAdder_501_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1654_io_ci = FullAdder_502_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1655_io_a = FullAdder_503_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1655_io_b = FullAdder_504_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1655_io_ci = FullAdder_505_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1656_io_a = FullAdder_506_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1656_io_b = FullAdder_507_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1656_io_ci = FullAdder_508_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1657_io_a = FullAdder_509_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1657_io_b = FullAdder_510_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1657_io_ci = FullAdder_511_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_47_io_a = FullAdder_512_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_47_io_b = HalfAdder_15_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1658_io_a = FullAdder_495_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1658_io_b = FullAdder_496_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1658_io_ci = FullAdder_497_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1659_io_a = FullAdder_498_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1659_io_b = FullAdder_499_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1659_io_ci = FullAdder_500_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1660_io_a = FullAdder_501_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1660_io_b = FullAdder_502_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1660_io_ci = FullAdder_503_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1661_io_a = FullAdder_504_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1661_io_b = FullAdder_505_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1661_io_ci = FullAdder_506_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1662_io_a = FullAdder_507_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1662_io_b = FullAdder_508_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1662_io_ci = FullAdder_509_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1663_io_a = FullAdder_510_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1663_io_b = FullAdder_511_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1663_io_ci = FullAdder_512_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1664_io_a = HalfAdder_15_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1664_io_b = FullAdder_513_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1664_io_ci = FullAdder_514_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1665_io_a = FullAdder_515_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1665_io_b = FullAdder_516_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1665_io_ci = FullAdder_517_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1666_io_a = FullAdder_518_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1666_io_b = FullAdder_519_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1666_io_ci = FullAdder_520_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1667_io_a = FullAdder_521_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1667_io_b = FullAdder_522_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1667_io_ci = FullAdder_523_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1668_io_a = FullAdder_524_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1668_io_b = FullAdder_525_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1668_io_ci = FullAdder_526_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1669_io_a = FullAdder_527_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1669_io_b = FullAdder_528_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1669_io_ci = FullAdder_529_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_48_io_a = FullAdder_530_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_48_io_b = FullAdder_531_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1670_io_a = FullAdder_513_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1670_io_b = FullAdder_514_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1670_io_ci = FullAdder_515_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1671_io_a = FullAdder_516_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1671_io_b = FullAdder_517_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1671_io_ci = FullAdder_518_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1672_io_a = FullAdder_519_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1672_io_b = FullAdder_520_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1672_io_ci = FullAdder_521_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1673_io_a = FullAdder_522_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1673_io_b = FullAdder_523_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1673_io_ci = FullAdder_524_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1674_io_a = FullAdder_525_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1674_io_b = FullAdder_526_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1674_io_ci = FullAdder_527_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1675_io_a = FullAdder_528_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1675_io_b = FullAdder_529_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1675_io_ci = FullAdder_530_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1676_io_a = FullAdder_531_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1676_io_b = FullAdder_532_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1676_io_ci = FullAdder_533_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1677_io_a = FullAdder_534_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1677_io_b = FullAdder_535_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1677_io_ci = FullAdder_536_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1678_io_a = FullAdder_537_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1678_io_b = FullAdder_538_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1678_io_ci = FullAdder_539_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1679_io_a = FullAdder_540_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1679_io_b = FullAdder_541_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1679_io_ci = FullAdder_542_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1680_io_a = FullAdder_543_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1680_io_b = FullAdder_544_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1680_io_ci = FullAdder_545_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1681_io_a = FullAdder_546_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1681_io_b = FullAdder_547_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1681_io_ci = FullAdder_548_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1682_io_a = io_pp_63[6]; // @[wallace.scala 69:18]
  assign FullAdder_1682_io_b = FullAdder_532_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1682_io_ci = FullAdder_533_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1683_io_a = FullAdder_534_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1683_io_b = FullAdder_535_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1683_io_ci = FullAdder_536_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1684_io_a = FullAdder_537_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1684_io_b = FullAdder_538_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1684_io_ci = FullAdder_539_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1685_io_a = FullAdder_540_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1685_io_b = FullAdder_541_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1685_io_ci = FullAdder_542_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1686_io_a = FullAdder_543_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1686_io_b = FullAdder_544_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1686_io_ci = FullAdder_545_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1687_io_a = FullAdder_546_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1687_io_b = FullAdder_547_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1687_io_ci = FullAdder_548_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1688_io_a = FullAdder_549_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1688_io_b = FullAdder_550_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1688_io_ci = FullAdder_551_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1689_io_a = FullAdder_552_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1689_io_b = FullAdder_553_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1689_io_ci = FullAdder_554_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1690_io_a = FullAdder_555_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1690_io_b = FullAdder_556_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1690_io_ci = FullAdder_557_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1691_io_a = FullAdder_558_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1691_io_b = FullAdder_559_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1691_io_ci = FullAdder_560_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1692_io_a = FullAdder_561_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1692_io_b = FullAdder_562_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1692_io_ci = FullAdder_563_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1693_io_a = FullAdder_564_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1693_io_b = FullAdder_565_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1693_io_ci = FullAdder_566_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1694_io_a = FullAdder_567_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1694_io_b = FullAdder_568_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1694_io_ci = FullAdder_569_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1695_io_a = FullAdder_551_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1695_io_b = FullAdder_552_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1695_io_ci = FullAdder_553_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1696_io_a = FullAdder_554_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1696_io_b = FullAdder_555_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1696_io_ci = FullAdder_556_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1697_io_a = FullAdder_557_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1697_io_b = FullAdder_558_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1697_io_ci = FullAdder_559_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1698_io_a = FullAdder_560_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1698_io_b = FullAdder_561_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1698_io_ci = FullAdder_562_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1699_io_a = FullAdder_563_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1699_io_b = FullAdder_564_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1699_io_ci = FullAdder_565_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1700_io_a = FullAdder_566_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1700_io_b = FullAdder_567_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1700_io_ci = FullAdder_568_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1701_io_a = FullAdder_569_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1701_io_b = HalfAdder_16_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1701_io_ci = FullAdder_570_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1702_io_a = FullAdder_571_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1702_io_b = FullAdder_572_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1702_io_ci = FullAdder_573_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1703_io_a = FullAdder_574_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1703_io_b = FullAdder_575_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1703_io_ci = FullAdder_576_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1704_io_a = FullAdder_577_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1704_io_b = FullAdder_578_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1704_io_ci = FullAdder_579_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1705_io_a = FullAdder_580_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1705_io_b = FullAdder_581_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1705_io_ci = FullAdder_582_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1706_io_a = FullAdder_583_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1706_io_b = FullAdder_584_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1706_io_ci = FullAdder_585_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1707_io_a = FullAdder_586_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1707_io_b = FullAdder_587_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1707_io_ci = FullAdder_588_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1708_io_a = FullAdder_570_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1708_io_b = FullAdder_571_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1708_io_ci = FullAdder_572_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1709_io_a = FullAdder_573_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1709_io_b = FullAdder_574_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1709_io_ci = FullAdder_575_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1710_io_a = FullAdder_576_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1710_io_b = FullAdder_577_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1710_io_ci = FullAdder_578_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1711_io_a = FullAdder_579_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1711_io_b = FullAdder_580_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1711_io_ci = FullAdder_581_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1712_io_a = FullAdder_582_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1712_io_b = FullAdder_583_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1712_io_ci = FullAdder_584_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1713_io_a = FullAdder_585_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1713_io_b = FullAdder_586_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1713_io_ci = FullAdder_587_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1714_io_a = FullAdder_588_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1714_io_b = FullAdder_589_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1714_io_ci = FullAdder_590_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1715_io_a = FullAdder_591_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1715_io_b = FullAdder_592_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1715_io_ci = FullAdder_593_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1716_io_a = FullAdder_594_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1716_io_b = FullAdder_595_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1716_io_ci = FullAdder_596_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1717_io_a = FullAdder_597_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1717_io_b = FullAdder_598_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1717_io_ci = FullAdder_599_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1718_io_a = FullAdder_600_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1718_io_b = FullAdder_601_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1718_io_ci = FullAdder_602_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1719_io_a = FullAdder_603_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1719_io_b = FullAdder_604_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1719_io_ci = FullAdder_605_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1720_io_a = FullAdder_606_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1720_io_b = FullAdder_607_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1720_io_ci = FullAdder_608_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1721_io_a = io_pp_63[3]; // @[wallace.scala 69:18]
  assign FullAdder_1721_io_b = FullAdder_590_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1721_io_ci = FullAdder_591_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1722_io_a = FullAdder_592_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1722_io_b = FullAdder_593_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1722_io_ci = FullAdder_594_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1723_io_a = FullAdder_595_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1723_io_b = FullAdder_596_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1723_io_ci = FullAdder_597_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1724_io_a = FullAdder_598_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1724_io_b = FullAdder_599_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1724_io_ci = FullAdder_600_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1725_io_a = FullAdder_601_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1725_io_b = FullAdder_602_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1725_io_ci = FullAdder_603_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1726_io_a = FullAdder_604_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1726_io_b = FullAdder_605_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1726_io_ci = FullAdder_606_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1727_io_a = FullAdder_607_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1727_io_b = FullAdder_608_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1727_io_ci = FullAdder_609_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1728_io_a = FullAdder_610_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1728_io_b = FullAdder_611_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1728_io_ci = FullAdder_612_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1729_io_a = FullAdder_613_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1729_io_b = FullAdder_614_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1729_io_ci = FullAdder_615_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1730_io_a = FullAdder_616_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1730_io_b = FullAdder_617_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1730_io_ci = FullAdder_618_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1731_io_a = FullAdder_619_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1731_io_b = FullAdder_620_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1731_io_ci = FullAdder_621_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1732_io_a = FullAdder_622_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1732_io_b = FullAdder_623_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1732_io_ci = FullAdder_624_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1733_io_a = FullAdder_625_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1733_io_b = FullAdder_626_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1733_io_ci = FullAdder_627_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1734_io_a = FullAdder_628_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1734_io_b = FullAdder_629_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1734_io_ci = HalfAdder_17_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1735_io_a = FullAdder_610_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1735_io_b = FullAdder_611_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1735_io_ci = FullAdder_612_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1736_io_a = FullAdder_613_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1736_io_b = FullAdder_614_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1736_io_ci = FullAdder_615_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1737_io_a = FullAdder_616_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1737_io_b = FullAdder_617_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1737_io_ci = FullAdder_618_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1738_io_a = FullAdder_619_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1738_io_b = FullAdder_620_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1738_io_ci = FullAdder_621_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1739_io_a = FullAdder_622_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1739_io_b = FullAdder_623_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1739_io_ci = FullAdder_624_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1740_io_a = FullAdder_625_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1740_io_b = FullAdder_626_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1740_io_ci = FullAdder_627_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1741_io_a = FullAdder_628_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1741_io_b = FullAdder_629_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1741_io_ci = HalfAdder_17_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1742_io_a = FullAdder_630_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1742_io_b = FullAdder_631_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1742_io_ci = FullAdder_632_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1743_io_a = FullAdder_633_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1743_io_b = FullAdder_634_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1743_io_ci = FullAdder_635_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1744_io_a = FullAdder_636_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1744_io_b = FullAdder_637_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1744_io_ci = FullAdder_638_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1745_io_a = FullAdder_639_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1745_io_b = FullAdder_640_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1745_io_ci = FullAdder_641_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1746_io_a = FullAdder_642_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1746_io_b = FullAdder_643_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1746_io_ci = FullAdder_644_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1747_io_a = FullAdder_645_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1747_io_b = FullAdder_646_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1747_io_ci = FullAdder_647_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1748_io_a = FullAdder_648_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1748_io_b = FullAdder_649_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1748_io_ci = FullAdder_650_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1749_io_a = FullAdder_630_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1749_io_b = FullAdder_631_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1749_io_ci = FullAdder_632_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1750_io_a = FullAdder_633_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1750_io_b = FullAdder_634_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1750_io_ci = FullAdder_635_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1751_io_a = FullAdder_636_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1751_io_b = FullAdder_637_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1751_io_ci = FullAdder_638_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1752_io_a = FullAdder_639_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1752_io_b = FullAdder_640_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1752_io_ci = FullAdder_641_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1753_io_a = FullAdder_642_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1753_io_b = FullAdder_643_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1753_io_ci = FullAdder_644_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1754_io_a = FullAdder_645_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1754_io_b = FullAdder_646_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1754_io_ci = FullAdder_647_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1755_io_a = FullAdder_648_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1755_io_b = FullAdder_649_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1755_io_ci = FullAdder_650_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1756_io_a = FullAdder_651_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1756_io_b = FullAdder_652_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1756_io_ci = FullAdder_653_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1757_io_a = FullAdder_654_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1757_io_b = FullAdder_655_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1757_io_ci = FullAdder_656_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1758_io_a = FullAdder_657_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1758_io_b = FullAdder_658_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1758_io_ci = FullAdder_659_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1759_io_a = FullAdder_660_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1759_io_b = FullAdder_661_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1759_io_ci = FullAdder_662_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1760_io_a = FullAdder_663_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1760_io_b = FullAdder_664_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1760_io_ci = FullAdder_665_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1761_io_a = FullAdder_666_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1761_io_b = FullAdder_667_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1761_io_ci = FullAdder_668_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1762_io_a = FullAdder_669_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1762_io_b = FullAdder_670_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1762_io_ci = FullAdder_671_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1763_io_a = io_pp_63[0]; // @[wallace.scala 69:18]
  assign FullAdder_1763_io_b = FullAdder_651_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1763_io_ci = FullAdder_652_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1764_io_a = FullAdder_653_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1764_io_b = FullAdder_654_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1764_io_ci = FullAdder_655_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1765_io_a = FullAdder_656_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1765_io_b = FullAdder_657_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1765_io_ci = FullAdder_658_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1766_io_a = FullAdder_659_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1766_io_b = FullAdder_660_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1766_io_ci = FullAdder_661_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1767_io_a = FullAdder_662_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1767_io_b = FullAdder_663_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1767_io_ci = FullAdder_664_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1768_io_a = FullAdder_665_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1768_io_b = FullAdder_666_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1768_io_ci = FullAdder_667_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1769_io_a = FullAdder_668_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1769_io_b = FullAdder_669_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1769_io_ci = FullAdder_670_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1770_io_a = FullAdder_671_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1770_io_b = FullAdder_672_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1770_io_ci = FullAdder_673_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1771_io_a = FullAdder_674_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1771_io_b = FullAdder_675_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1771_io_ci = FullAdder_676_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1772_io_a = FullAdder_677_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1772_io_b = FullAdder_678_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1772_io_ci = FullAdder_679_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1773_io_a = FullAdder_680_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1773_io_b = FullAdder_681_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1773_io_ci = FullAdder_682_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1774_io_a = FullAdder_683_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1774_io_b = FullAdder_684_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1774_io_ci = FullAdder_685_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1775_io_a = FullAdder_686_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1775_io_b = FullAdder_687_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1775_io_ci = FullAdder_688_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1776_io_a = FullAdder_689_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1776_io_b = FullAdder_690_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1776_io_ci = FullAdder_691_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1777_io_a = FullAdder_672_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1777_io_b = FullAdder_673_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1777_io_ci = FullAdder_674_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1778_io_a = FullAdder_675_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1778_io_b = FullAdder_676_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1778_io_ci = FullAdder_677_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1779_io_a = FullAdder_678_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1779_io_b = FullAdder_679_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1779_io_ci = FullAdder_680_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1780_io_a = FullAdder_681_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1780_io_b = FullAdder_682_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1780_io_ci = FullAdder_683_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1781_io_a = FullAdder_684_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1781_io_b = FullAdder_685_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1781_io_ci = FullAdder_686_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1782_io_a = FullAdder_687_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1782_io_b = FullAdder_688_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1782_io_ci = FullAdder_689_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1783_io_a = FullAdder_690_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1783_io_b = FullAdder_691_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1783_io_ci = FullAdder_692_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1784_io_a = FullAdder_693_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1784_io_b = FullAdder_694_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1784_io_ci = FullAdder_695_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1785_io_a = FullAdder_696_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1785_io_b = FullAdder_697_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1785_io_ci = FullAdder_698_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1786_io_a = FullAdder_699_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1786_io_b = FullAdder_700_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1786_io_ci = FullAdder_701_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1787_io_a = FullAdder_702_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1787_io_b = FullAdder_703_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1787_io_ci = FullAdder_704_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1788_io_a = FullAdder_705_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1788_io_b = FullAdder_706_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1788_io_ci = FullAdder_707_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1789_io_a = FullAdder_708_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1789_io_b = FullAdder_709_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1789_io_ci = FullAdder_710_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1790_io_a = FullAdder_711_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1790_io_b = FullAdder_712_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1790_io_ci = HalfAdder_18_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1791_io_a = FullAdder_693_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1791_io_b = FullAdder_694_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1791_io_ci = FullAdder_695_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1792_io_a = FullAdder_696_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1792_io_b = FullAdder_697_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1792_io_ci = FullAdder_698_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1793_io_a = FullAdder_699_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1793_io_b = FullAdder_700_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1793_io_ci = FullAdder_701_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1794_io_a = FullAdder_702_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1794_io_b = FullAdder_703_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1794_io_ci = FullAdder_704_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1795_io_a = FullAdder_705_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1795_io_b = FullAdder_706_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1795_io_ci = FullAdder_707_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1796_io_a = FullAdder_708_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1796_io_b = FullAdder_709_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1796_io_ci = FullAdder_710_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1797_io_a = FullAdder_711_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1797_io_b = FullAdder_712_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1797_io_ci = HalfAdder_18_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1798_io_a = FullAdder_713_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1798_io_b = FullAdder_714_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1798_io_ci = FullAdder_715_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1799_io_a = FullAdder_716_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1799_io_b = FullAdder_717_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1799_io_ci = FullAdder_718_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1800_io_a = FullAdder_719_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1800_io_b = FullAdder_720_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1800_io_ci = FullAdder_721_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1801_io_a = FullAdder_722_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1801_io_b = FullAdder_723_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1801_io_ci = FullAdder_724_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1802_io_a = FullAdder_725_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1802_io_b = FullAdder_726_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1802_io_ci = FullAdder_727_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1803_io_a = FullAdder_728_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1803_io_b = FullAdder_729_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1803_io_ci = FullAdder_730_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_49_io_a = FullAdder_731_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_49_io_b = FullAdder_732_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1804_io_a = io_pp_60[0]; // @[wallace.scala 69:18]
  assign FullAdder_1804_io_b = FullAdder_713_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1804_io_ci = FullAdder_714_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1805_io_a = FullAdder_715_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1805_io_b = FullAdder_716_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1805_io_ci = FullAdder_717_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1806_io_a = FullAdder_718_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1806_io_b = FullAdder_719_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1806_io_ci = FullAdder_720_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1807_io_a = FullAdder_721_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1807_io_b = FullAdder_722_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1807_io_ci = FullAdder_723_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1808_io_a = FullAdder_724_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1808_io_b = FullAdder_725_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1808_io_ci = FullAdder_726_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1809_io_a = FullAdder_727_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1809_io_b = FullAdder_728_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1809_io_ci = FullAdder_729_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1810_io_a = FullAdder_730_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1810_io_b = FullAdder_731_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1810_io_ci = FullAdder_732_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1811_io_a = FullAdder_733_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1811_io_b = FullAdder_734_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1811_io_ci = FullAdder_735_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1812_io_a = FullAdder_736_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1812_io_b = FullAdder_737_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1812_io_ci = FullAdder_738_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1813_io_a = FullAdder_739_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1813_io_b = FullAdder_740_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1813_io_ci = FullAdder_741_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1814_io_a = FullAdder_742_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1814_io_b = FullAdder_743_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1814_io_ci = FullAdder_744_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1815_io_a = FullAdder_745_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1815_io_b = FullAdder_746_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1815_io_ci = FullAdder_747_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1816_io_a = FullAdder_748_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1816_io_b = FullAdder_749_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1816_io_ci = FullAdder_750_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1817_io_a = FullAdder_733_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1817_io_b = FullAdder_734_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1817_io_ci = FullAdder_735_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1818_io_a = FullAdder_736_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1818_io_b = FullAdder_737_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1818_io_ci = FullAdder_738_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1819_io_a = FullAdder_739_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1819_io_b = FullAdder_740_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1819_io_ci = FullAdder_741_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1820_io_a = FullAdder_742_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1820_io_b = FullAdder_743_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1820_io_ci = FullAdder_744_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1821_io_a = FullAdder_745_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1821_io_b = FullAdder_746_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1821_io_ci = FullAdder_747_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1822_io_a = FullAdder_748_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1822_io_b = FullAdder_749_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1822_io_ci = FullAdder_750_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1823_io_a = FullAdder_751_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1823_io_b = FullAdder_752_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1823_io_ci = FullAdder_753_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1824_io_a = FullAdder_754_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1824_io_b = FullAdder_755_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1824_io_ci = FullAdder_756_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1825_io_a = FullAdder_757_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1825_io_b = FullAdder_758_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1825_io_ci = FullAdder_759_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1826_io_a = FullAdder_760_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1826_io_b = FullAdder_761_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1826_io_ci = FullAdder_762_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1827_io_a = FullAdder_763_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1827_io_b = FullAdder_764_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1827_io_ci = FullAdder_765_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1828_io_a = FullAdder_766_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1828_io_b = FullAdder_767_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1828_io_ci = FullAdder_768_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1829_io_a = FullAdder_769_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1829_io_b = FullAdder_770_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1829_io_ci = FullAdder_771_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1830_io_a = FullAdder_753_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1830_io_b = FullAdder_754_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1830_io_ci = FullAdder_755_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1831_io_a = FullAdder_756_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1831_io_b = FullAdder_757_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1831_io_ci = FullAdder_758_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1832_io_a = FullAdder_759_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1832_io_b = FullAdder_760_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1832_io_ci = FullAdder_761_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1833_io_a = FullAdder_762_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1833_io_b = FullAdder_763_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1833_io_ci = FullAdder_764_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1834_io_a = FullAdder_765_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1834_io_b = FullAdder_766_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1834_io_ci = FullAdder_767_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1835_io_a = FullAdder_768_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1835_io_b = FullAdder_769_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1835_io_ci = FullAdder_770_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1836_io_a = FullAdder_771_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1836_io_b = HalfAdder_19_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1836_io_ci = FullAdder_772_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1837_io_a = FullAdder_773_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1837_io_b = FullAdder_774_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1837_io_ci = FullAdder_775_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1838_io_a = FullAdder_776_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1838_io_b = FullAdder_777_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1838_io_ci = FullAdder_778_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1839_io_a = FullAdder_779_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1839_io_b = FullAdder_780_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1839_io_ci = FullAdder_781_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1840_io_a = FullAdder_782_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1840_io_b = FullAdder_783_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1840_io_ci = FullAdder_784_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1841_io_a = FullAdder_785_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1841_io_b = FullAdder_786_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1841_io_ci = FullAdder_787_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1842_io_a = FullAdder_788_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1842_io_b = FullAdder_789_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1842_io_ci = FullAdder_790_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1843_io_a = io_pp_57[0]; // @[wallace.scala 69:18]
  assign FullAdder_1843_io_b = FullAdder_772_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1843_io_ci = FullAdder_773_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1844_io_a = FullAdder_774_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1844_io_b = FullAdder_775_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1844_io_ci = FullAdder_776_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1845_io_a = FullAdder_777_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1845_io_b = FullAdder_778_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1845_io_ci = FullAdder_779_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1846_io_a = FullAdder_780_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1846_io_b = FullAdder_781_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1846_io_ci = FullAdder_782_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1847_io_a = FullAdder_783_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1847_io_b = FullAdder_784_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1847_io_ci = FullAdder_785_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1848_io_a = FullAdder_786_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1848_io_b = FullAdder_787_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1848_io_ci = FullAdder_788_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1849_io_a = FullAdder_789_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1849_io_b = FullAdder_790_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1849_io_ci = FullAdder_791_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1850_io_a = FullAdder_792_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1850_io_b = FullAdder_793_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1850_io_ci = FullAdder_794_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1851_io_a = FullAdder_795_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1851_io_b = FullAdder_796_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1851_io_ci = FullAdder_797_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1852_io_a = FullAdder_798_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1852_io_b = FullAdder_799_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1852_io_ci = FullAdder_800_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1853_io_a = FullAdder_801_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1853_io_b = FullAdder_802_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1853_io_ci = FullAdder_803_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1854_io_a = FullAdder_804_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1854_io_b = FullAdder_805_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1854_io_ci = FullAdder_806_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1855_io_a = FullAdder_807_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1855_io_b = FullAdder_808_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1855_io_ci = FullAdder_809_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1856_io_a = FullAdder_791_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1856_io_b = FullAdder_792_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1856_io_ci = FullAdder_793_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1857_io_a = FullAdder_794_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1857_io_b = FullAdder_795_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1857_io_ci = FullAdder_796_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1858_io_a = FullAdder_797_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1858_io_b = FullAdder_798_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1858_io_ci = FullAdder_799_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1859_io_a = FullAdder_800_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1859_io_b = FullAdder_801_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1859_io_ci = FullAdder_802_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1860_io_a = FullAdder_803_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1860_io_b = FullAdder_804_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1860_io_ci = FullAdder_805_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1861_io_a = FullAdder_806_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1861_io_b = FullAdder_807_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1861_io_ci = FullAdder_808_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1862_io_a = FullAdder_809_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1862_io_b = FullAdder_810_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1862_io_ci = FullAdder_811_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1863_io_a = FullAdder_812_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1863_io_b = FullAdder_813_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1863_io_ci = FullAdder_814_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1864_io_a = FullAdder_815_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1864_io_b = FullAdder_816_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1864_io_ci = FullAdder_817_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1865_io_a = FullAdder_818_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1865_io_b = FullAdder_819_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1865_io_ci = FullAdder_820_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1866_io_a = FullAdder_821_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1866_io_b = FullAdder_822_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1866_io_ci = FullAdder_823_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1867_io_a = FullAdder_824_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1867_io_b = FullAdder_825_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1867_io_ci = FullAdder_826_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1868_io_a = io_pp_54[1]; // @[wallace.scala 69:18]
  assign FullAdder_1868_io_b = io_pp_55[0]; // @[wallace.scala 70:18]
  assign FullAdder_1868_io_ci = FullAdder_810_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1869_io_a = FullAdder_811_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1869_io_b = FullAdder_812_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1869_io_ci = FullAdder_813_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1870_io_a = FullAdder_814_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1870_io_b = FullAdder_815_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1870_io_ci = FullAdder_816_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1871_io_a = FullAdder_817_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1871_io_b = FullAdder_818_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1871_io_ci = FullAdder_819_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1872_io_a = FullAdder_820_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1872_io_b = FullAdder_821_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1872_io_ci = FullAdder_822_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1873_io_a = FullAdder_823_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1873_io_b = FullAdder_824_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1873_io_ci = FullAdder_825_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1874_io_a = FullAdder_826_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1874_io_b = FullAdder_827_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1874_io_ci = FullAdder_828_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1875_io_a = FullAdder_829_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1875_io_b = FullAdder_830_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1875_io_ci = FullAdder_831_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1876_io_a = FullAdder_832_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1876_io_b = FullAdder_833_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1876_io_ci = FullAdder_834_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1877_io_a = FullAdder_835_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1877_io_b = FullAdder_836_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1877_io_ci = FullAdder_837_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1878_io_a = FullAdder_838_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1878_io_b = FullAdder_839_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1878_io_ci = FullAdder_840_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1879_io_a = FullAdder_841_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1879_io_b = FullAdder_842_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1879_io_ci = FullAdder_843_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1880_io_a = io_pp_54[0]; // @[wallace.scala 69:18]
  assign FullAdder_1880_io_b = FullAdder_828_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1880_io_ci = FullAdder_829_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1881_io_a = FullAdder_830_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1881_io_b = FullAdder_831_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1881_io_ci = FullAdder_832_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1882_io_a = FullAdder_833_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1882_io_b = FullAdder_834_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1882_io_ci = FullAdder_835_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1883_io_a = FullAdder_836_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1883_io_b = FullAdder_837_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1883_io_ci = FullAdder_838_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1884_io_a = FullAdder_839_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1884_io_b = FullAdder_840_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1884_io_ci = FullAdder_841_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1885_io_a = FullAdder_842_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1885_io_b = FullAdder_843_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1885_io_ci = FullAdder_844_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1886_io_a = FullAdder_845_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1886_io_b = FullAdder_846_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1886_io_ci = FullAdder_847_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1887_io_a = FullAdder_848_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1887_io_b = FullAdder_849_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1887_io_ci = FullAdder_850_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1888_io_a = FullAdder_851_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1888_io_b = FullAdder_852_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1888_io_ci = FullAdder_853_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1889_io_a = FullAdder_854_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1889_io_b = FullAdder_855_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1889_io_ci = FullAdder_856_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1890_io_a = FullAdder_857_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1890_io_b = FullAdder_858_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1890_io_ci = FullAdder_859_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1891_io_a = FullAdder_860_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1891_io_b = FullAdder_861_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1891_io_ci = FullAdder_862_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1892_io_a = FullAdder_846_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1892_io_b = FullAdder_847_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1892_io_ci = FullAdder_848_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1893_io_a = FullAdder_849_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1893_io_b = FullAdder_850_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1893_io_ci = FullAdder_851_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1894_io_a = FullAdder_852_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1894_io_b = FullAdder_853_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1894_io_ci = FullAdder_854_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1895_io_a = FullAdder_855_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1895_io_b = FullAdder_856_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1895_io_ci = FullAdder_857_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1896_io_a = FullAdder_858_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1896_io_b = FullAdder_859_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1896_io_ci = FullAdder_860_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1897_io_a = FullAdder_861_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1897_io_b = FullAdder_862_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1897_io_ci = FullAdder_863_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1898_io_a = FullAdder_864_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1898_io_b = FullAdder_865_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1898_io_ci = FullAdder_866_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1899_io_a = FullAdder_867_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1899_io_b = FullAdder_868_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1899_io_ci = FullAdder_869_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1900_io_a = FullAdder_870_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1900_io_b = FullAdder_871_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1900_io_ci = FullAdder_872_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1901_io_a = FullAdder_873_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1901_io_b = FullAdder_874_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1901_io_ci = FullAdder_875_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1902_io_a = FullAdder_876_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1902_io_b = FullAdder_877_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1902_io_ci = FullAdder_878_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1903_io_a = FullAdder_879_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1903_io_b = FullAdder_880_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1903_io_ci = HalfAdder_20_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1904_io_a = FullAdder_864_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1904_io_b = FullAdder_865_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1904_io_ci = FullAdder_866_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1905_io_a = FullAdder_867_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1905_io_b = FullAdder_868_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1905_io_ci = FullAdder_869_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1906_io_a = FullAdder_870_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1906_io_b = FullAdder_871_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1906_io_ci = FullAdder_872_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1907_io_a = FullAdder_873_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1907_io_b = FullAdder_874_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1907_io_ci = FullAdder_875_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1908_io_a = FullAdder_876_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1908_io_b = FullAdder_877_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1908_io_ci = FullAdder_878_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1909_io_a = FullAdder_879_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1909_io_b = FullAdder_880_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1909_io_ci = HalfAdder_20_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1910_io_a = FullAdder_881_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1910_io_b = FullAdder_882_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1910_io_ci = FullAdder_883_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1911_io_a = FullAdder_884_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1911_io_b = FullAdder_885_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1911_io_ci = FullAdder_886_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1912_io_a = FullAdder_887_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1912_io_b = FullAdder_888_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1912_io_ci = FullAdder_889_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1913_io_a = FullAdder_890_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1913_io_b = FullAdder_891_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1913_io_ci = FullAdder_892_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1914_io_a = FullAdder_893_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1914_io_b = FullAdder_894_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1914_io_ci = FullAdder_895_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1915_io_a = io_pp_51[0]; // @[wallace.scala 69:18]
  assign FullAdder_1915_io_b = FullAdder_881_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1915_io_ci = FullAdder_882_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1916_io_a = FullAdder_883_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1916_io_b = FullAdder_884_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1916_io_ci = FullAdder_885_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1917_io_a = FullAdder_886_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1917_io_b = FullAdder_887_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1917_io_ci = FullAdder_888_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1918_io_a = FullAdder_889_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1918_io_b = FullAdder_890_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1918_io_ci = FullAdder_891_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1919_io_a = FullAdder_892_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1919_io_b = FullAdder_893_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1919_io_ci = FullAdder_894_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1920_io_a = FullAdder_895_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1920_io_b = FullAdder_896_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1920_io_ci = FullAdder_897_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1921_io_a = FullAdder_898_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1921_io_b = FullAdder_899_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1921_io_ci = FullAdder_900_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1922_io_a = FullAdder_901_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1922_io_b = FullAdder_902_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1922_io_ci = FullAdder_903_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1923_io_a = FullAdder_904_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1923_io_b = FullAdder_905_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1923_io_ci = FullAdder_906_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1924_io_a = FullAdder_907_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1924_io_b = FullAdder_908_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1924_io_ci = FullAdder_909_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1925_io_a = FullAdder_910_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1925_io_b = FullAdder_911_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1925_io_ci = FullAdder_912_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_50_io_a = FullAdder_913_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_50_io_b = FullAdder_914_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1926_io_a = FullAdder_898_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1926_io_b = FullAdder_899_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1926_io_ci = FullAdder_900_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1927_io_a = FullAdder_901_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1927_io_b = FullAdder_902_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1927_io_ci = FullAdder_903_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1928_io_a = FullAdder_904_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1928_io_b = FullAdder_905_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1928_io_ci = FullAdder_906_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1929_io_a = FullAdder_907_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1929_io_b = FullAdder_908_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1929_io_ci = FullAdder_909_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1930_io_a = FullAdder_910_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1930_io_b = FullAdder_911_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1930_io_ci = FullAdder_912_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1931_io_a = FullAdder_913_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1931_io_b = FullAdder_914_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1931_io_ci = FullAdder_915_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1932_io_a = FullAdder_916_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1932_io_b = FullAdder_917_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1932_io_ci = FullAdder_918_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1933_io_a = FullAdder_919_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1933_io_b = FullAdder_920_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1933_io_ci = FullAdder_921_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1934_io_a = FullAdder_922_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1934_io_b = FullAdder_923_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1934_io_ci = FullAdder_924_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1935_io_a = FullAdder_925_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1935_io_b = FullAdder_926_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1935_io_ci = FullAdder_927_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1936_io_a = FullAdder_928_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1936_io_b = FullAdder_929_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1936_io_ci = FullAdder_930_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1937_io_a = io_pp_48[1]; // @[wallace.scala 69:18]
  assign FullAdder_1937_io_b = io_pp_49[0]; // @[wallace.scala 70:18]
  assign FullAdder_1937_io_ci = FullAdder_915_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1938_io_a = FullAdder_916_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1938_io_b = FullAdder_917_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1938_io_ci = FullAdder_918_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1939_io_a = FullAdder_919_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1939_io_b = FullAdder_920_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1939_io_ci = FullAdder_921_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1940_io_a = FullAdder_922_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1940_io_b = FullAdder_923_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1940_io_ci = FullAdder_924_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1941_io_a = FullAdder_925_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1941_io_b = FullAdder_926_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1941_io_ci = FullAdder_927_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1942_io_a = FullAdder_928_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1942_io_b = FullAdder_929_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1942_io_ci = FullAdder_930_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1943_io_a = FullAdder_931_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1943_io_b = FullAdder_932_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1943_io_ci = FullAdder_933_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1944_io_a = FullAdder_934_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1944_io_b = FullAdder_935_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1944_io_ci = FullAdder_936_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1945_io_a = FullAdder_937_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1945_io_b = FullAdder_938_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1945_io_ci = FullAdder_939_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1946_io_a = FullAdder_940_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1946_io_b = FullAdder_941_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1946_io_ci = FullAdder_942_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1947_io_a = FullAdder_943_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1947_io_b = FullAdder_944_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1947_io_ci = FullAdder_945_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1948_io_a = io_pp_48[0]; // @[wallace.scala 69:18]
  assign FullAdder_1948_io_b = FullAdder_931_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1948_io_ci = FullAdder_932_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1949_io_a = FullAdder_933_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1949_io_b = FullAdder_934_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1949_io_ci = FullAdder_935_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1950_io_a = FullAdder_936_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1950_io_b = FullAdder_937_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1950_io_ci = FullAdder_938_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1951_io_a = FullAdder_939_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1951_io_b = FullAdder_940_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1951_io_ci = FullAdder_941_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1952_io_a = FullAdder_942_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1952_io_b = FullAdder_943_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1952_io_ci = FullAdder_944_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1953_io_a = FullAdder_945_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1953_io_b = FullAdder_946_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1953_io_ci = FullAdder_947_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1954_io_a = FullAdder_948_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1954_io_b = FullAdder_949_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1954_io_ci = FullAdder_950_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1955_io_a = FullAdder_951_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1955_io_b = FullAdder_952_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1955_io_ci = FullAdder_953_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1956_io_a = FullAdder_954_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1956_io_b = FullAdder_955_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1956_io_ci = FullAdder_956_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1957_io_a = FullAdder_957_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1957_io_b = FullAdder_958_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1957_io_ci = FullAdder_959_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1958_io_a = FullAdder_960_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1958_io_b = FullAdder_961_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1958_io_ci = FullAdder_962_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1959_io_a = FullAdder_947_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1959_io_b = FullAdder_948_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1959_io_ci = FullAdder_949_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1960_io_a = FullAdder_950_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1960_io_b = FullAdder_951_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1960_io_ci = FullAdder_952_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1961_io_a = FullAdder_953_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1961_io_b = FullAdder_954_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1961_io_ci = FullAdder_955_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1962_io_a = FullAdder_956_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1962_io_b = FullAdder_957_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1962_io_ci = FullAdder_958_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1963_io_a = FullAdder_959_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1963_io_b = FullAdder_960_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1963_io_ci = FullAdder_961_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1964_io_a = FullAdder_962_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1964_io_b = FullAdder_963_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1964_io_ci = FullAdder_964_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1965_io_a = FullAdder_965_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1965_io_b = FullAdder_966_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1965_io_ci = FullAdder_967_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1966_io_a = FullAdder_968_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1966_io_b = FullAdder_969_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1966_io_ci = FullAdder_970_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1967_io_a = FullAdder_971_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1967_io_b = FullAdder_972_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1967_io_ci = FullAdder_973_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1968_io_a = FullAdder_974_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1968_io_b = FullAdder_975_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1968_io_ci = FullAdder_976_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_51_io_a = FullAdder_977_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_51_io_b = HalfAdder_21_io_co; // @[wallace.scala 60:18]
  assign FullAdder_1969_io_a = FullAdder_963_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1969_io_b = FullAdder_964_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1969_io_ci = FullAdder_965_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1970_io_a = FullAdder_966_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1970_io_b = FullAdder_967_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1970_io_ci = FullAdder_968_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1971_io_a = FullAdder_969_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1971_io_b = FullAdder_970_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1971_io_ci = FullAdder_971_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1972_io_a = FullAdder_972_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1972_io_b = FullAdder_973_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1972_io_ci = FullAdder_974_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1973_io_a = FullAdder_975_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1973_io_b = FullAdder_976_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1973_io_ci = FullAdder_977_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1974_io_a = HalfAdder_21_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1974_io_b = FullAdder_978_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1974_io_ci = FullAdder_979_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1975_io_a = FullAdder_980_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1975_io_b = FullAdder_981_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1975_io_ci = FullAdder_982_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1976_io_a = FullAdder_983_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1976_io_b = FullAdder_984_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1976_io_ci = FullAdder_985_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1977_io_a = FullAdder_986_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1977_io_b = FullAdder_987_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1977_io_ci = FullAdder_988_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1978_io_a = FullAdder_989_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1978_io_b = FullAdder_990_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1978_io_ci = FullAdder_991_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1979_io_a = io_pp_45[0]; // @[wallace.scala 69:18]
  assign FullAdder_1979_io_b = FullAdder_978_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1979_io_ci = FullAdder_979_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1980_io_a = FullAdder_980_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1980_io_b = FullAdder_981_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1980_io_ci = FullAdder_982_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1981_io_a = FullAdder_983_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1981_io_b = FullAdder_984_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1981_io_ci = FullAdder_985_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1982_io_a = FullAdder_986_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1982_io_b = FullAdder_987_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1982_io_ci = FullAdder_988_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1983_io_a = FullAdder_989_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1983_io_b = FullAdder_990_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1983_io_ci = FullAdder_991_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1984_io_a = FullAdder_992_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1984_io_b = FullAdder_993_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1984_io_ci = FullAdder_994_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1985_io_a = FullAdder_995_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1985_io_b = FullAdder_996_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1985_io_ci = FullAdder_997_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1986_io_a = FullAdder_998_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1986_io_b = FullAdder_999_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1986_io_ci = FullAdder_1000_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1987_io_a = FullAdder_1001_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1987_io_b = FullAdder_1002_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1987_io_ci = FullAdder_1003_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1988_io_a = FullAdder_1004_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1988_io_b = FullAdder_1005_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1988_io_ci = FullAdder_1006_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1989_io_a = FullAdder_993_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1989_io_b = FullAdder_994_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1989_io_ci = FullAdder_995_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1990_io_a = FullAdder_996_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1990_io_b = FullAdder_997_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1990_io_ci = FullAdder_998_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1991_io_a = FullAdder_999_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1991_io_b = FullAdder_1000_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1991_io_ci = FullAdder_1001_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1992_io_a = FullAdder_1002_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1992_io_b = FullAdder_1003_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1992_io_ci = FullAdder_1004_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1993_io_a = FullAdder_1005_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1993_io_b = FullAdder_1006_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1993_io_ci = FullAdder_1007_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1994_io_a = FullAdder_1008_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1994_io_b = FullAdder_1009_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1994_io_ci = FullAdder_1010_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1995_io_a = FullAdder_1011_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1995_io_b = FullAdder_1012_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1995_io_ci = FullAdder_1013_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1996_io_a = FullAdder_1014_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1996_io_b = FullAdder_1015_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1996_io_ci = FullAdder_1016_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1997_io_a = FullAdder_1017_io_co; // @[wallace.scala 69:18]
  assign FullAdder_1997_io_b = FullAdder_1018_io_co; // @[wallace.scala 70:18]
  assign FullAdder_1997_io_ci = FullAdder_1019_io_co; // @[wallace.scala 71:19]
  assign FullAdder_1998_io_a = io_pp_42[1]; // @[wallace.scala 69:18]
  assign FullAdder_1998_io_b = io_pp_43[0]; // @[wallace.scala 70:18]
  assign FullAdder_1998_io_ci = FullAdder_1008_io_s; // @[wallace.scala 71:19]
  assign FullAdder_1999_io_a = FullAdder_1009_io_s; // @[wallace.scala 69:18]
  assign FullAdder_1999_io_b = FullAdder_1010_io_s; // @[wallace.scala 70:18]
  assign FullAdder_1999_io_ci = FullAdder_1011_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2000_io_a = FullAdder_1012_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2000_io_b = FullAdder_1013_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2000_io_ci = FullAdder_1014_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2001_io_a = FullAdder_1015_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2001_io_b = FullAdder_1016_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2001_io_ci = FullAdder_1017_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2002_io_a = FullAdder_1018_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2002_io_b = FullAdder_1019_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2002_io_ci = FullAdder_1020_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2003_io_a = FullAdder_1021_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2003_io_b = FullAdder_1022_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2003_io_ci = FullAdder_1023_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2004_io_a = FullAdder_1024_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2004_io_b = FullAdder_1025_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2004_io_ci = FullAdder_1026_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2005_io_a = FullAdder_1027_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2005_io_b = FullAdder_1028_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2005_io_ci = FullAdder_1029_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2006_io_a = FullAdder_1030_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2006_io_b = FullAdder_1031_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2006_io_ci = FullAdder_1032_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2007_io_a = FullAdder_1033_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2007_io_b = FullAdder_1034_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2007_io_ci = FullAdder_1035_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2008_io_a = io_pp_42[0]; // @[wallace.scala 69:18]
  assign FullAdder_2008_io_b = FullAdder_1022_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2008_io_ci = FullAdder_1023_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2009_io_a = FullAdder_1024_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2009_io_b = FullAdder_1025_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2009_io_ci = FullAdder_1026_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2010_io_a = FullAdder_1027_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2010_io_b = FullAdder_1028_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2010_io_ci = FullAdder_1029_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2011_io_a = FullAdder_1030_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2011_io_b = FullAdder_1031_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2011_io_ci = FullAdder_1032_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2012_io_a = FullAdder_1033_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2012_io_b = FullAdder_1034_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2012_io_ci = FullAdder_1035_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2013_io_a = FullAdder_1036_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2013_io_b = FullAdder_1037_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2013_io_ci = FullAdder_1038_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2014_io_a = FullAdder_1039_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2014_io_b = FullAdder_1040_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2014_io_ci = FullAdder_1041_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2015_io_a = FullAdder_1042_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2015_io_b = FullAdder_1043_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2015_io_ci = FullAdder_1044_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2016_io_a = FullAdder_1045_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2016_io_b = FullAdder_1046_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2016_io_ci = FullAdder_1047_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_52_io_a = FullAdder_1048_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_52_io_b = FullAdder_1049_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2017_io_a = FullAdder_1036_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2017_io_b = FullAdder_1037_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2017_io_ci = FullAdder_1038_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2018_io_a = FullAdder_1039_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2018_io_b = FullAdder_1040_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2018_io_ci = FullAdder_1041_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2019_io_a = FullAdder_1042_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2019_io_b = FullAdder_1043_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2019_io_ci = FullAdder_1044_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2020_io_a = FullAdder_1045_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2020_io_b = FullAdder_1046_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2020_io_ci = FullAdder_1047_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2021_io_a = FullAdder_1048_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2021_io_b = FullAdder_1049_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2021_io_ci = FullAdder_1050_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2022_io_a = FullAdder_1051_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2022_io_b = FullAdder_1052_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2022_io_ci = FullAdder_1053_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2023_io_a = FullAdder_1054_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2023_io_b = FullAdder_1055_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2023_io_ci = FullAdder_1056_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2024_io_a = FullAdder_1057_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2024_io_b = FullAdder_1058_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2024_io_ci = FullAdder_1059_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2025_io_a = FullAdder_1060_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2025_io_b = FullAdder_1061_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2025_io_ci = FullAdder_1062_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2026_io_a = io_pp_39[1]; // @[wallace.scala 69:18]
  assign FullAdder_2026_io_b = io_pp_40[0]; // @[wallace.scala 70:18]
  assign FullAdder_2026_io_ci = FullAdder_1050_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2027_io_a = FullAdder_1051_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2027_io_b = FullAdder_1052_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2027_io_ci = FullAdder_1053_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2028_io_a = FullAdder_1054_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2028_io_b = FullAdder_1055_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2028_io_ci = FullAdder_1056_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2029_io_a = FullAdder_1057_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2029_io_b = FullAdder_1058_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2029_io_ci = FullAdder_1059_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2030_io_a = FullAdder_1060_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2030_io_b = FullAdder_1061_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2030_io_ci = FullAdder_1062_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2031_io_a = FullAdder_1063_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2031_io_b = FullAdder_1064_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2031_io_ci = FullAdder_1065_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2032_io_a = FullAdder_1066_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2032_io_b = FullAdder_1067_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2032_io_ci = FullAdder_1068_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2033_io_a = FullAdder_1069_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2033_io_b = FullAdder_1070_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2033_io_ci = FullAdder_1071_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2034_io_a = FullAdder_1072_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2034_io_b = FullAdder_1073_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2034_io_ci = FullAdder_1074_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2035_io_a = io_pp_39[0]; // @[wallace.scala 69:18]
  assign FullAdder_2035_io_b = FullAdder_1063_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2035_io_ci = FullAdder_1064_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2036_io_a = FullAdder_1065_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2036_io_b = FullAdder_1066_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2036_io_ci = FullAdder_1067_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2037_io_a = FullAdder_1068_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2037_io_b = FullAdder_1069_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2037_io_ci = FullAdder_1070_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2038_io_a = FullAdder_1071_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2038_io_b = FullAdder_1072_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2038_io_ci = FullAdder_1073_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2039_io_a = FullAdder_1074_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2039_io_b = FullAdder_1075_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2039_io_ci = FullAdder_1076_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2040_io_a = FullAdder_1077_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2040_io_b = FullAdder_1078_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2040_io_ci = FullAdder_1079_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2041_io_a = FullAdder_1080_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2041_io_b = FullAdder_1081_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2041_io_ci = FullAdder_1082_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2042_io_a = FullAdder_1083_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2042_io_b = FullAdder_1084_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2042_io_ci = FullAdder_1085_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2043_io_a = FullAdder_1086_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2043_io_b = FullAdder_1087_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2043_io_ci = FullAdder_1088_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2044_io_a = FullAdder_1076_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2044_io_b = FullAdder_1077_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2044_io_ci = FullAdder_1078_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2045_io_a = FullAdder_1079_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2045_io_b = FullAdder_1080_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2045_io_ci = FullAdder_1081_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2046_io_a = FullAdder_1082_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2046_io_b = FullAdder_1083_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2046_io_ci = FullAdder_1084_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2047_io_a = FullAdder_1085_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2047_io_b = FullAdder_1086_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2047_io_ci = FullAdder_1087_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2048_io_a = FullAdder_1088_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2048_io_b = FullAdder_1089_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2048_io_ci = FullAdder_1090_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2049_io_a = FullAdder_1091_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2049_io_b = FullAdder_1092_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2049_io_ci = FullAdder_1093_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2050_io_a = FullAdder_1094_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2050_io_b = FullAdder_1095_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2050_io_ci = FullAdder_1096_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2051_io_a = FullAdder_1097_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2051_io_b = FullAdder_1098_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2051_io_ci = FullAdder_1099_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_53_io_a = FullAdder_1100_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_53_io_b = HalfAdder_22_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2052_io_a = FullAdder_1089_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2052_io_b = FullAdder_1090_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2052_io_ci = FullAdder_1091_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2053_io_a = FullAdder_1092_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2053_io_b = FullAdder_1093_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2053_io_ci = FullAdder_1094_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2054_io_a = FullAdder_1095_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2054_io_b = FullAdder_1096_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2054_io_ci = FullAdder_1097_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2055_io_a = FullAdder_1098_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2055_io_b = FullAdder_1099_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2055_io_ci = FullAdder_1100_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2056_io_a = HalfAdder_22_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2056_io_b = FullAdder_1101_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2056_io_ci = FullAdder_1102_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2057_io_a = FullAdder_1103_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2057_io_b = FullAdder_1104_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2057_io_ci = FullAdder_1105_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2058_io_a = FullAdder_1106_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2058_io_b = FullAdder_1107_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2058_io_ci = FullAdder_1108_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2059_io_a = FullAdder_1109_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2059_io_b = FullAdder_1110_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2059_io_ci = FullAdder_1111_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2060_io_a = io_pp_36[0]; // @[wallace.scala 69:18]
  assign FullAdder_2060_io_b = FullAdder_1101_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2060_io_ci = FullAdder_1102_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2061_io_a = FullAdder_1103_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2061_io_b = FullAdder_1104_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2061_io_ci = FullAdder_1105_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2062_io_a = FullAdder_1106_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2062_io_b = FullAdder_1107_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2062_io_ci = FullAdder_1108_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2063_io_a = FullAdder_1109_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2063_io_b = FullAdder_1110_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2063_io_ci = FullAdder_1111_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2064_io_a = FullAdder_1112_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2064_io_b = FullAdder_1113_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2064_io_ci = FullAdder_1114_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2065_io_a = FullAdder_1115_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2065_io_b = FullAdder_1116_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2065_io_ci = FullAdder_1117_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2066_io_a = FullAdder_1118_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2066_io_b = FullAdder_1119_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2066_io_ci = FullAdder_1120_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2067_io_a = FullAdder_1121_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2067_io_b = FullAdder_1122_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2067_io_ci = FullAdder_1123_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2068_io_a = FullAdder_1113_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2068_io_b = FullAdder_1114_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2068_io_ci = FullAdder_1115_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2069_io_a = FullAdder_1116_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2069_io_b = FullAdder_1117_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2069_io_ci = FullAdder_1118_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2070_io_a = FullAdder_1119_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2070_io_b = FullAdder_1120_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2070_io_ci = FullAdder_1121_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2071_io_a = FullAdder_1122_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2071_io_b = FullAdder_1123_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2071_io_ci = FullAdder_1124_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2072_io_a = FullAdder_1125_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2072_io_b = FullAdder_1126_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2072_io_ci = FullAdder_1127_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2073_io_a = FullAdder_1128_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2073_io_b = FullAdder_1129_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2073_io_ci = FullAdder_1130_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2074_io_a = FullAdder_1131_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2074_io_b = FullAdder_1132_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2074_io_ci = FullAdder_1133_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2075_io_a = FullAdder_1134_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2075_io_b = FullAdder_1135_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2075_io_ci = HalfAdder_23_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2076_io_a = FullAdder_1125_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2076_io_b = FullAdder_1126_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2076_io_ci = FullAdder_1127_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2077_io_a = FullAdder_1128_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2077_io_b = FullAdder_1129_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2077_io_ci = FullAdder_1130_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2078_io_a = FullAdder_1131_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2078_io_b = FullAdder_1132_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2078_io_ci = FullAdder_1133_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2079_io_a = FullAdder_1134_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2079_io_b = FullAdder_1135_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2079_io_ci = HalfAdder_23_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2080_io_a = FullAdder_1136_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2080_io_b = FullAdder_1137_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2080_io_ci = FullAdder_1138_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2081_io_a = FullAdder_1139_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2081_io_b = FullAdder_1140_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2081_io_ci = FullAdder_1141_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2082_io_a = FullAdder_1142_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2082_io_b = FullAdder_1143_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2082_io_ci = FullAdder_1144_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2083_io_a = io_pp_33[0]; // @[wallace.scala 69:18]
  assign FullAdder_2083_io_b = FullAdder_1136_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2083_io_ci = FullAdder_1137_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2084_io_a = FullAdder_1138_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2084_io_b = FullAdder_1139_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2084_io_ci = FullAdder_1140_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2085_io_a = FullAdder_1141_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2085_io_b = FullAdder_1142_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2085_io_ci = FullAdder_1143_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2086_io_a = FullAdder_1144_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2086_io_b = FullAdder_1145_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2086_io_ci = FullAdder_1146_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2087_io_a = FullAdder_1147_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2087_io_b = FullAdder_1148_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2087_io_ci = FullAdder_1149_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2088_io_a = FullAdder_1150_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2088_io_b = FullAdder_1151_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2088_io_ci = FullAdder_1152_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2089_io_a = FullAdder_1153_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2089_io_b = FullAdder_1154_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2089_io_ci = FullAdder_1155_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_54_io_a = FullAdder_1156_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_54_io_b = FullAdder_1157_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2090_io_a = FullAdder_1147_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2090_io_b = FullAdder_1148_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2090_io_ci = FullAdder_1149_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2091_io_a = FullAdder_1150_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2091_io_b = FullAdder_1151_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2091_io_ci = FullAdder_1152_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2092_io_a = FullAdder_1153_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2092_io_b = FullAdder_1154_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2092_io_ci = FullAdder_1155_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2093_io_a = FullAdder_1156_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2093_io_b = FullAdder_1157_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2093_io_ci = FullAdder_1158_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2094_io_a = FullAdder_1159_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2094_io_b = FullAdder_1160_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2094_io_ci = FullAdder_1161_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2095_io_a = FullAdder_1162_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2095_io_b = FullAdder_1163_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2095_io_ci = FullAdder_1164_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2096_io_a = FullAdder_1165_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2096_io_b = FullAdder_1166_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2096_io_ci = FullAdder_1167_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2097_io_a = FullAdder_1158_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2097_io_b = FullAdder_1159_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2097_io_ci = FullAdder_1160_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2098_io_a = FullAdder_1161_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2098_io_b = FullAdder_1162_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2098_io_ci = FullAdder_1163_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2099_io_a = FullAdder_1164_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2099_io_b = FullAdder_1165_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2099_io_ci = FullAdder_1166_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2100_io_a = FullAdder_1167_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2100_io_b = HalfAdder_24_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2100_io_ci = FullAdder_1168_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2101_io_a = FullAdder_1169_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2101_io_b = FullAdder_1170_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2101_io_ci = FullAdder_1171_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2102_io_a = FullAdder_1172_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2102_io_b = FullAdder_1173_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2102_io_ci = FullAdder_1174_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2103_io_a = FullAdder_1175_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2103_io_b = FullAdder_1176_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2103_io_ci = FullAdder_1177_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2104_io_a = io_pp_30[0]; // @[wallace.scala 69:18]
  assign FullAdder_2104_io_b = FullAdder_1168_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2104_io_ci = FullAdder_1169_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2105_io_a = FullAdder_1170_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2105_io_b = FullAdder_1171_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2105_io_ci = FullAdder_1172_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2106_io_a = FullAdder_1173_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2106_io_b = FullAdder_1174_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2106_io_ci = FullAdder_1175_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2107_io_a = FullAdder_1176_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2107_io_b = FullAdder_1177_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2107_io_ci = FullAdder_1178_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2108_io_a = FullAdder_1179_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2108_io_b = FullAdder_1180_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2108_io_ci = FullAdder_1181_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2109_io_a = FullAdder_1182_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2109_io_b = FullAdder_1183_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2109_io_ci = FullAdder_1184_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2110_io_a = FullAdder_1185_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2110_io_b = FullAdder_1186_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2110_io_ci = FullAdder_1187_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2111_io_a = FullAdder_1178_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2111_io_b = FullAdder_1179_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2111_io_ci = FullAdder_1180_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2112_io_a = FullAdder_1181_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2112_io_b = FullAdder_1182_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2112_io_ci = FullAdder_1183_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2113_io_a = FullAdder_1184_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2113_io_b = FullAdder_1185_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2113_io_ci = FullAdder_1186_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2114_io_a = FullAdder_1187_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2114_io_b = FullAdder_1188_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2114_io_ci = FullAdder_1189_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2115_io_a = FullAdder_1190_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2115_io_b = FullAdder_1191_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2115_io_ci = FullAdder_1192_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2116_io_a = FullAdder_1193_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2116_io_b = FullAdder_1194_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2116_io_ci = FullAdder_1195_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_55_io_a = FullAdder_1196_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_55_io_b = HalfAdder_25_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2117_io_a = FullAdder_1188_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2117_io_b = FullAdder_1189_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2117_io_ci = FullAdder_1190_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2118_io_a = FullAdder_1191_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2118_io_b = FullAdder_1192_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2118_io_ci = FullAdder_1193_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2119_io_a = FullAdder_1194_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2119_io_b = FullAdder_1195_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2119_io_ci = FullAdder_1196_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2120_io_a = HalfAdder_25_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2120_io_b = FullAdder_1197_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2120_io_ci = FullAdder_1198_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2121_io_a = FullAdder_1199_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2121_io_b = FullAdder_1200_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2121_io_ci = FullAdder_1201_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2122_io_a = FullAdder_1202_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2122_io_b = FullAdder_1203_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2122_io_ci = FullAdder_1204_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2123_io_a = io_pp_27[0]; // @[wallace.scala 69:18]
  assign FullAdder_2123_io_b = FullAdder_1197_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2123_io_ci = FullAdder_1198_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2124_io_a = FullAdder_1199_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2124_io_b = FullAdder_1200_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2124_io_ci = FullAdder_1201_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2125_io_a = FullAdder_1202_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2125_io_b = FullAdder_1203_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2125_io_ci = FullAdder_1204_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2126_io_a = FullAdder_1205_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2126_io_b = FullAdder_1206_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2126_io_ci = FullAdder_1207_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2127_io_a = FullAdder_1208_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2127_io_b = FullAdder_1209_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2127_io_ci = FullAdder_1210_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2128_io_a = FullAdder_1211_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2128_io_b = FullAdder_1212_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2128_io_ci = FullAdder_1213_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2129_io_a = FullAdder_1206_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2129_io_b = FullAdder_1207_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2129_io_ci = FullAdder_1208_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2130_io_a = FullAdder_1209_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2130_io_b = FullAdder_1210_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2130_io_ci = FullAdder_1211_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2131_io_a = FullAdder_1212_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2131_io_b = FullAdder_1213_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2131_io_ci = FullAdder_1214_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2132_io_a = FullAdder_1215_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2132_io_b = FullAdder_1216_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2132_io_ci = FullAdder_1217_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2133_io_a = FullAdder_1218_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2133_io_b = FullAdder_1219_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2133_io_ci = FullAdder_1220_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_56_io_a = FullAdder_1221_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_56_io_b = FullAdder_1222_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2134_io_a = io_pp_24[1]; // @[wallace.scala 69:18]
  assign FullAdder_2134_io_b = io_pp_25[0]; // @[wallace.scala 70:18]
  assign FullAdder_2134_io_ci = FullAdder_1215_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2135_io_a = FullAdder_1216_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2135_io_b = FullAdder_1217_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2135_io_ci = FullAdder_1218_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2136_io_a = FullAdder_1219_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2136_io_b = FullAdder_1220_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2136_io_ci = FullAdder_1221_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2137_io_a = FullAdder_1222_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2137_io_b = FullAdder_1223_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2137_io_ci = FullAdder_1224_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2138_io_a = FullAdder_1225_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2138_io_b = FullAdder_1226_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2138_io_ci = FullAdder_1227_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2139_io_a = FullAdder_1228_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2139_io_b = FullAdder_1229_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2139_io_ci = FullAdder_1230_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2140_io_a = io_pp_24[0]; // @[wallace.scala 69:18]
  assign FullAdder_2140_io_b = FullAdder_1223_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2140_io_ci = FullAdder_1224_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2141_io_a = FullAdder_1225_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2141_io_b = FullAdder_1226_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2141_io_ci = FullAdder_1227_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2142_io_a = FullAdder_1228_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2142_io_b = FullAdder_1229_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2142_io_ci = FullAdder_1230_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2143_io_a = FullAdder_1231_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2143_io_b = FullAdder_1232_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2143_io_ci = FullAdder_1233_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2144_io_a = FullAdder_1234_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2144_io_b = FullAdder_1235_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2144_io_ci = FullAdder_1236_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2145_io_a = FullAdder_1231_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2145_io_b = FullAdder_1232_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2145_io_ci = FullAdder_1233_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2146_io_a = FullAdder_1234_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2146_io_b = FullAdder_1235_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2146_io_ci = FullAdder_1236_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2147_io_a = FullAdder_1237_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2147_io_b = FullAdder_1238_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2147_io_ci = FullAdder_1239_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2148_io_a = FullAdder_1240_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2148_io_b = FullAdder_1241_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2148_io_ci = FullAdder_1242_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2149_io_a = FullAdder_1243_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2149_io_b = FullAdder_1244_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2149_io_ci = FullAdder_1245_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2150_io_a = FullAdder_1239_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2150_io_b = FullAdder_1240_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2150_io_ci = FullAdder_1241_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2151_io_a = FullAdder_1242_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2151_io_b = FullAdder_1243_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2151_io_ci = FullAdder_1244_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2152_io_a = FullAdder_1245_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2152_io_b = HalfAdder_26_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2152_io_ci = FullAdder_1246_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2153_io_a = FullAdder_1247_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2153_io_b = FullAdder_1248_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2153_io_ci = FullAdder_1249_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2154_io_a = FullAdder_1250_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2154_io_b = FullAdder_1251_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2154_io_ci = FullAdder_1252_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2155_io_a = io_pp_21[0]; // @[wallace.scala 69:18]
  assign FullAdder_2155_io_b = FullAdder_1246_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2155_io_ci = FullAdder_1247_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2156_io_a = FullAdder_1248_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2156_io_b = FullAdder_1249_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2156_io_ci = FullAdder_1250_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2157_io_a = FullAdder_1251_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2157_io_b = FullAdder_1252_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2157_io_ci = FullAdder_1253_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2158_io_a = FullAdder_1254_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2158_io_b = FullAdder_1255_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2158_io_ci = FullAdder_1256_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2159_io_a = FullAdder_1257_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2159_io_b = FullAdder_1258_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2159_io_ci = FullAdder_1259_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2160_io_a = FullAdder_1253_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2160_io_b = FullAdder_1254_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2160_io_ci = FullAdder_1255_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2161_io_a = FullAdder_1256_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2161_io_b = FullAdder_1257_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2161_io_ci = FullAdder_1258_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2162_io_a = FullAdder_1259_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2162_io_b = FullAdder_1260_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2162_io_ci = FullAdder_1261_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2163_io_a = FullAdder_1262_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2163_io_b = FullAdder_1263_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2163_io_ci = FullAdder_1264_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_57_io_a = FullAdder_1265_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_57_io_b = HalfAdder_27_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2164_io_a = FullAdder_1260_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2164_io_b = FullAdder_1261_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2164_io_ci = FullAdder_1262_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2165_io_a = FullAdder_1263_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2165_io_b = FullAdder_1264_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2165_io_ci = FullAdder_1265_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2166_io_a = HalfAdder_27_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2166_io_b = FullAdder_1266_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2166_io_ci = FullAdder_1267_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2167_io_a = FullAdder_1268_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2167_io_b = FullAdder_1269_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2167_io_ci = FullAdder_1270_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2168_io_a = io_pp_18[0]; // @[wallace.scala 69:18]
  assign FullAdder_2168_io_b = FullAdder_1266_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2168_io_ci = FullAdder_1267_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2169_io_a = FullAdder_1268_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2169_io_b = FullAdder_1269_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2169_io_ci = FullAdder_1270_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2170_io_a = FullAdder_1271_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2170_io_b = FullAdder_1272_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2170_io_ci = FullAdder_1273_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2171_io_a = FullAdder_1274_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2171_io_b = FullAdder_1275_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2171_io_ci = FullAdder_1276_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2172_io_a = FullAdder_1272_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2172_io_b = FullAdder_1273_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2172_io_ci = FullAdder_1274_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2173_io_a = FullAdder_1275_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2173_io_b = FullAdder_1276_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2173_io_ci = FullAdder_1277_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2174_io_a = FullAdder_1278_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2174_io_b = FullAdder_1279_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2174_io_ci = FullAdder_1280_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2175_io_a = FullAdder_1281_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2175_io_b = FullAdder_1282_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2175_io_ci = HalfAdder_28_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2176_io_a = FullAdder_1278_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2176_io_b = FullAdder_1279_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2176_io_ci = FullAdder_1280_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2177_io_a = FullAdder_1281_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2177_io_b = FullAdder_1282_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2177_io_ci = HalfAdder_28_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2178_io_a = FullAdder_1283_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2178_io_b = FullAdder_1284_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2178_io_ci = FullAdder_1285_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_58_io_a = FullAdder_1286_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_58_io_b = FullAdder_1287_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2179_io_a = io_pp_15[0]; // @[wallace.scala 69:18]
  assign FullAdder_2179_io_b = FullAdder_1283_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2179_io_ci = FullAdder_1284_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2180_io_a = FullAdder_1285_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2180_io_b = FullAdder_1286_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2180_io_ci = FullAdder_1287_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2181_io_a = FullAdder_1288_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2181_io_b = FullAdder_1289_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2181_io_ci = FullAdder_1290_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_59_io_a = FullAdder_1291_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_59_io_b = FullAdder_1292_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2182_io_a = FullAdder_1288_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2182_io_b = FullAdder_1289_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2182_io_ci = FullAdder_1290_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2183_io_a = FullAdder_1291_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2183_io_b = FullAdder_1292_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2183_io_ci = FullAdder_1293_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2184_io_a = FullAdder_1294_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2184_io_b = FullAdder_1295_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2184_io_ci = FullAdder_1296_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2185_io_a = FullAdder_1293_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2185_io_b = FullAdder_1294_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2185_io_ci = FullAdder_1295_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2186_io_a = FullAdder_1296_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2186_io_b = HalfAdder_29_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2186_io_ci = FullAdder_1297_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2187_io_a = FullAdder_1298_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2187_io_b = FullAdder_1299_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2187_io_ci = FullAdder_1300_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2188_io_a = io_pp_12[0]; // @[wallace.scala 69:18]
  assign FullAdder_2188_io_b = FullAdder_1297_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2188_io_ci = FullAdder_1298_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2189_io_a = FullAdder_1299_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2189_io_b = FullAdder_1300_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2189_io_ci = FullAdder_1301_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2190_io_a = FullAdder_1302_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2190_io_b = FullAdder_1303_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2190_io_ci = FullAdder_1304_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2191_io_a = FullAdder_1301_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2191_io_b = FullAdder_1302_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2191_io_ci = FullAdder_1303_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2192_io_a = FullAdder_1304_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2192_io_b = FullAdder_1305_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2192_io_ci = FullAdder_1306_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2193_io_a = FullAdder_1305_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2193_io_b = FullAdder_1306_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2193_io_ci = FullAdder_1307_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_60_io_a = HalfAdder_30_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_60_io_b = FullAdder_1308_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_61_io_a = FullAdder_1309_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_61_io_b = FullAdder_1310_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2194_io_a = io_pp_9[0]; // @[wallace.scala 69:18]
  assign FullAdder_2194_io_b = FullAdder_1308_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2194_io_ci = FullAdder_1309_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2195_io_a = FullAdder_1310_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2195_io_b = FullAdder_1311_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2195_io_ci = FullAdder_1312_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2196_io_a = FullAdder_1311_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2196_io_b = FullAdder_1312_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2196_io_ci = FullAdder_1313_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2197_io_a = FullAdder_1314_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2197_io_b = FullAdder_1315_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2197_io_ci = HalfAdder_31_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2198_io_a = FullAdder_1314_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2198_io_b = FullAdder_1315_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2198_io_ci = HalfAdder_31_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_62_io_a = FullAdder_1316_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_62_io_b = FullAdder_1317_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2199_io_a = io_pp_6[0]; // @[wallace.scala 69:18]
  assign FullAdder_2199_io_b = FullAdder_1316_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2199_io_ci = FullAdder_1317_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_63_io_a = FullAdder_1318_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_63_io_b = FullAdder_1319_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2200_io_a = FullAdder_1318_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2200_io_b = FullAdder_1319_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2200_io_ci = FullAdder_1320_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_64_io_a = FullAdder_1320_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_64_io_b = HalfAdder_32_io_s; // @[wallace.scala 60:18]
  assign FullAdder_2201_io_a = io_pp_3[0]; // @[wallace.scala 69:18]
  assign FullAdder_2201_io_b = FullAdder_1321_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2201_io_ci = HalfAdder_33_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_65_io_a = io_pp_2[0]; // @[wallace.scala 59:18]
  assign HalfAdder_65_io_b = HalfAdder_33_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_66_io_a = HalfAdder_34_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_66_io_b = HalfAdder_35_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_67_io_a = HalfAdder_35_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_67_io_b = HalfAdder_36_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_68_io_a = HalfAdder_36_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_68_io_b = FullAdder_1322_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_69_io_a = HalfAdder_1_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_69_io_b = FullAdder_1322_io_s; // @[wallace.scala 60:18]
  assign FullAdder_2202_io_a = FullAdder_4_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2202_io_b = FullAdder_1323_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2202_io_ci = FullAdder_1324_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2203_io_a = FullAdder_6_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2203_io_b = FullAdder_1324_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2203_io_ci = FullAdder_1325_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_70_io_a = FullAdder_1325_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_70_io_b = FullAdder_1326_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_71_io_a = FullAdder_1327_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_71_io_b = FullAdder_1328_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2204_io_a = FullAdder_1327_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2204_io_b = FullAdder_1328_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2204_io_ci = FullAdder_1329_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2205_io_a = FullAdder_1329_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2205_io_b = FullAdder_1330_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2205_io_ci = FullAdder_1331_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2206_io_a = FullAdder_17_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2206_io_b = HalfAdder_3_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2206_io_ci = FullAdder_1331_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2207_io_a = FullAdder_1332_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2207_io_b = FullAdder_1333_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2207_io_ci = FullAdder_1334_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2208_io_a = FullAdder_1333_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2208_io_b = FullAdder_1334_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2208_io_ci = HalfAdder_37_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2209_io_a = FullAdder_1335_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2209_io_b = FullAdder_1336_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2209_io_ci = HalfAdder_38_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2210_io_a = FullAdder_1335_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2210_io_b = FullAdder_1336_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2210_io_ci = HalfAdder_38_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2211_io_a = FullAdder_1337_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2211_io_b = FullAdder_1338_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2211_io_ci = FullAdder_1339_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2212_io_a = FullAdder_1337_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2212_io_b = FullAdder_1338_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2212_io_ci = FullAdder_1339_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2213_io_a = FullAdder_1340_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2213_io_b = FullAdder_1341_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2213_io_ci = FullAdder_1342_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2214_io_a = FullAdder_33_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2214_io_b = FullAdder_34_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2214_io_ci = FullAdder_1340_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2215_io_a = FullAdder_1341_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2215_io_b = FullAdder_1342_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2215_io_ci = FullAdder_1343_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2216_io_a = FullAdder_39_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2216_io_b = FullAdder_1343_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2216_io_ci = FullAdder_1344_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2217_io_a = FullAdder_1345_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2217_io_b = FullAdder_1346_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2217_io_ci = FullAdder_1347_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_72_io_a = FullAdder_1348_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_72_io_b = FullAdder_1349_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2218_io_a = FullAdder_1346_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2218_io_b = FullAdder_1347_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2218_io_ci = FullAdder_1348_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2219_io_a = FullAdder_1349_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2219_io_b = FullAdder_1350_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2219_io_ci = FullAdder_1351_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2220_io_a = FullAdder_1350_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2220_io_b = FullAdder_1351_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2220_io_ci = FullAdder_1352_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2221_io_a = FullAdder_1353_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2221_io_b = FullAdder_1354_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2221_io_ci = FullAdder_1355_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_73_io_a = FullAdder_1356_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_73_io_b = FullAdder_1357_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2222_io_a = FullAdder_1354_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2222_io_b = FullAdder_1355_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2222_io_ci = FullAdder_1356_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2223_io_a = FullAdder_1357_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2223_io_b = FullAdder_1358_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2223_io_ci = FullAdder_1359_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2224_io_a = FullAdder_1360_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2224_io_b = FullAdder_1361_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2224_io_ci = HalfAdder_39_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2225_io_a = FullAdder_1358_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2225_io_b = FullAdder_1359_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2225_io_ci = FullAdder_1360_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2226_io_a = FullAdder_1361_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2226_io_b = HalfAdder_39_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2226_io_ci = FullAdder_1362_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2227_io_a = FullAdder_1363_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2227_io_b = FullAdder_1364_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2227_io_ci = FullAdder_1365_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2228_io_a = FullAdder_1362_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2228_io_b = FullAdder_1363_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2228_io_ci = FullAdder_1364_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2229_io_a = FullAdder_1365_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2229_io_b = HalfAdder_40_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2229_io_ci = FullAdder_1366_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2230_io_a = FullAdder_1367_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2230_io_b = FullAdder_1368_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2230_io_ci = FullAdder_1369_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2231_io_a = FullAdder_1366_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2231_io_b = FullAdder_1367_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2231_io_ci = FullAdder_1368_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2232_io_a = FullAdder_1369_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2232_io_b = HalfAdder_41_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2232_io_ci = FullAdder_1370_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2233_io_a = FullAdder_1371_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2233_io_b = FullAdder_1372_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2233_io_ci = FullAdder_1373_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2234_io_a = HalfAdder_6_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2234_io_b = FullAdder_1370_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2234_io_ci = FullAdder_1371_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2235_io_a = FullAdder_1372_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2235_io_b = FullAdder_1373_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2235_io_ci = FullAdder_1374_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2236_io_a = FullAdder_1375_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2236_io_b = FullAdder_1376_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2236_io_ci = FullAdder_1377_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2237_io_a = FullAdder_91_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2237_io_b = FullAdder_1375_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2237_io_ci = FullAdder_1376_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2238_io_a = FullAdder_1377_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2238_io_b = FullAdder_1378_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2238_io_ci = FullAdder_1379_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2239_io_a = FullAdder_1380_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2239_io_b = FullAdder_1381_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2239_io_ci = FullAdder_1382_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_74_io_a = FullAdder_1383_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_74_io_b = FullAdder_1384_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2240_io_a = FullAdder_99_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2240_io_b = FullAdder_1380_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2240_io_ci = FullAdder_1381_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2241_io_a = FullAdder_1382_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2241_io_b = FullAdder_1383_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2241_io_ci = FullAdder_1384_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2242_io_a = FullAdder_1385_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2242_io_b = FullAdder_1386_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2242_io_ci = FullAdder_1387_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2243_io_a = FullAdder_106_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2243_io_b = FullAdder_107_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2243_io_ci = FullAdder_1385_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2244_io_a = FullAdder_1386_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2244_io_b = FullAdder_1387_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2244_io_ci = FullAdder_1388_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2245_io_a = FullAdder_1389_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2245_io_b = FullAdder_1390_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2245_io_ci = FullAdder_1391_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2246_io_a = FullAdder_1392_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2246_io_b = FullAdder_1393_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2246_io_ci = FullAdder_1394_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2247_io_a = FullAdder_116_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2247_io_b = FullAdder_1390_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2247_io_ci = FullAdder_1391_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2248_io_a = FullAdder_1392_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2248_io_b = FullAdder_1393_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2248_io_ci = FullAdder_1394_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2249_io_a = FullAdder_1395_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2249_io_b = FullAdder_1396_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2249_io_ci = FullAdder_1397_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2250_io_a = FullAdder_1398_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2250_io_b = FullAdder_1399_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2250_io_ci = FullAdder_1400_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2251_io_a = FullAdder_1396_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2251_io_b = FullAdder_1397_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2251_io_ci = FullAdder_1398_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2252_io_a = FullAdder_1399_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2252_io_b = FullAdder_1400_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2252_io_ci = FullAdder_1401_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2253_io_a = FullAdder_1402_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2253_io_b = FullAdder_1403_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2253_io_ci = FullAdder_1404_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2254_io_a = FullAdder_1405_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2254_io_b = FullAdder_1406_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2254_io_ci = FullAdder_1407_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2255_io_a = FullAdder_134_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2255_io_b = FullAdder_1402_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2255_io_ci = FullAdder_1403_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2256_io_a = FullAdder_1404_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2256_io_b = FullAdder_1405_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2256_io_ci = FullAdder_1406_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2257_io_a = FullAdder_1407_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2257_io_b = FullAdder_1408_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2257_io_ci = FullAdder_1409_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2258_io_a = FullAdder_1410_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2258_io_b = FullAdder_1411_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2258_io_ci = FullAdder_1412_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2259_io_a = FullAdder_1408_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2259_io_b = FullAdder_1409_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2259_io_ci = FullAdder_1410_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2260_io_a = FullAdder_1411_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2260_io_b = FullAdder_1412_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2260_io_ci = FullAdder_1413_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2261_io_a = FullAdder_1414_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2261_io_b = FullAdder_1415_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2261_io_ci = FullAdder_1416_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2262_io_a = FullAdder_1417_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2262_io_b = FullAdder_1418_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2262_io_ci = FullAdder_1419_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2263_io_a = FullAdder_1415_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2263_io_b = FullAdder_1416_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2263_io_ci = FullAdder_1417_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2264_io_a = FullAdder_1418_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2264_io_b = FullAdder_1419_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2264_io_ci = FullAdder_1420_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2265_io_a = HalfAdder_42_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2265_io_b = FullAdder_1421_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2265_io_ci = FullAdder_1422_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2266_io_a = FullAdder_1423_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2266_io_b = FullAdder_1424_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2266_io_ci = FullAdder_1425_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2267_io_a = HalfAdder_7_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2267_io_b = FullAdder_1421_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2267_io_ci = FullAdder_1422_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2268_io_a = FullAdder_1423_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2268_io_b = FullAdder_1424_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2268_io_ci = FullAdder_1425_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2269_io_a = FullAdder_1426_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2269_io_b = FullAdder_1427_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2269_io_ci = FullAdder_1428_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2270_io_a = FullAdder_1429_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2270_io_b = FullAdder_1430_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2270_io_ci = FullAdder_1431_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2271_io_a = FullAdder_1432_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2271_io_b = FullAdder_1433_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2271_io_ci = FullAdder_1434_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2272_io_a = FullAdder_175_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2272_io_b = FullAdder_1428_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2272_io_ci = FullAdder_1429_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2273_io_a = FullAdder_1430_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2273_io_b = FullAdder_1431_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2273_io_ci = FullAdder_1432_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2274_io_a = FullAdder_1433_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2274_io_b = FullAdder_1434_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2274_io_ci = FullAdder_1435_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2275_io_a = FullAdder_1436_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2275_io_b = FullAdder_1437_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2275_io_ci = FullAdder_1438_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2276_io_a = FullAdder_1439_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2276_io_b = FullAdder_1440_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2276_io_ci = FullAdder_1441_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2277_io_a = FullAdder_186_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2277_io_b = FullAdder_1435_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2277_io_ci = FullAdder_1436_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2278_io_a = FullAdder_1437_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2278_io_b = FullAdder_1438_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2278_io_ci = FullAdder_1439_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2279_io_a = FullAdder_1440_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2279_io_b = FullAdder_1441_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2279_io_ci = FullAdder_1442_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2280_io_a = FullAdder_1443_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2280_io_b = FullAdder_1444_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2280_io_ci = FullAdder_1445_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2281_io_a = FullAdder_1446_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2281_io_b = FullAdder_1447_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2281_io_ci = FullAdder_1448_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2282_io_a = FullAdder_1442_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2282_io_b = FullAdder_1443_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2282_io_ci = FullAdder_1444_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2283_io_a = FullAdder_1445_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2283_io_b = FullAdder_1446_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2283_io_ci = FullAdder_1447_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2284_io_a = FullAdder_1448_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2284_io_b = FullAdder_1449_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2284_io_ci = FullAdder_1450_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2285_io_a = FullAdder_1451_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2285_io_b = FullAdder_1452_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2285_io_ci = FullAdder_1453_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2286_io_a = FullAdder_1454_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2286_io_b = FullAdder_1455_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2286_io_ci = FullAdder_1456_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2287_io_a = FullAdder_1450_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2287_io_b = FullAdder_1451_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2287_io_ci = FullAdder_1452_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2288_io_a = FullAdder_1453_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2288_io_b = FullAdder_1454_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2288_io_ci = FullAdder_1455_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2289_io_a = FullAdder_1456_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2289_io_b = FullAdder_1457_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2289_io_ci = FullAdder_1458_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2290_io_a = FullAdder_1459_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2290_io_b = FullAdder_1460_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2290_io_ci = FullAdder_1461_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2291_io_a = FullAdder_1462_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2291_io_b = FullAdder_1463_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2291_io_ci = FullAdder_1464_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2292_io_a = FullAdder_1458_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2292_io_b = FullAdder_1459_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2292_io_ci = FullAdder_1460_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2293_io_a = FullAdder_1461_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2293_io_b = FullAdder_1462_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2293_io_ci = FullAdder_1463_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2294_io_a = FullAdder_1464_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2294_io_b = FullAdder_1465_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2294_io_ci = FullAdder_1466_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2295_io_a = FullAdder_1467_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2295_io_b = FullAdder_1468_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2295_io_ci = FullAdder_1469_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2296_io_a = FullAdder_1470_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2296_io_b = FullAdder_1471_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2296_io_ci = FullAdder_1472_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2297_io_a = FullAdder_1466_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2297_io_b = FullAdder_1467_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2297_io_ci = FullAdder_1468_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2298_io_a = FullAdder_1469_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2298_io_b = FullAdder_1470_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2298_io_ci = FullAdder_1471_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2299_io_a = FullAdder_1472_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2299_io_b = FullAdder_1473_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2299_io_ci = HalfAdder_43_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2300_io_a = FullAdder_1474_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2300_io_b = FullAdder_1475_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2300_io_ci = FullAdder_1476_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2301_io_a = FullAdder_1477_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2301_io_b = FullAdder_1478_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2301_io_ci = FullAdder_1479_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2302_io_a = FullAdder_1480_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2302_io_b = FullAdder_1481_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2302_io_ci = HalfAdder_44_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2303_io_a = FullAdder_1474_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2303_io_b = FullAdder_1475_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2303_io_ci = FullAdder_1476_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2304_io_a = FullAdder_1477_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2304_io_b = FullAdder_1478_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2304_io_ci = FullAdder_1479_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2305_io_a = FullAdder_1480_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2305_io_b = FullAdder_1481_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2305_io_ci = HalfAdder_44_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2306_io_a = FullAdder_1482_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2306_io_b = FullAdder_1483_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2306_io_ci = FullAdder_1484_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2307_io_a = FullAdder_1485_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2307_io_b = FullAdder_1486_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2307_io_ci = FullAdder_1487_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2308_io_a = FullAdder_1488_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2308_io_b = FullAdder_1489_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2308_io_ci = HalfAdder_45_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2309_io_a = FullAdder_1482_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2309_io_b = FullAdder_1483_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2309_io_ci = FullAdder_1484_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2310_io_a = FullAdder_1485_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2310_io_b = FullAdder_1486_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2310_io_ci = FullAdder_1487_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2311_io_a = FullAdder_1488_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2311_io_b = FullAdder_1489_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2311_io_ci = HalfAdder_45_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2312_io_a = FullAdder_1490_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2312_io_b = FullAdder_1491_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2312_io_ci = FullAdder_1492_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2313_io_a = FullAdder_1493_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2313_io_b = FullAdder_1494_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2313_io_ci = FullAdder_1495_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2314_io_a = FullAdder_1496_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2314_io_b = FullAdder_1497_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2314_io_ci = FullAdder_1498_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2315_io_a = HalfAdder_10_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2315_io_b = FullAdder_1490_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2315_io_ci = FullAdder_1491_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2316_io_a = FullAdder_1492_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2316_io_b = FullAdder_1493_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2316_io_ci = FullAdder_1494_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2317_io_a = FullAdder_1495_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2317_io_b = FullAdder_1496_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2317_io_ci = FullAdder_1497_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2318_io_a = FullAdder_1498_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2318_io_b = FullAdder_1499_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2318_io_ci = FullAdder_1500_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2319_io_a = FullAdder_1501_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2319_io_b = FullAdder_1502_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2319_io_ci = FullAdder_1503_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2320_io_a = FullAdder_1504_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2320_io_b = FullAdder_1505_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2320_io_ci = FullAdder_1506_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2321_io_a = FullAdder_286_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2321_io_b = FullAdder_1499_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2321_io_ci = FullAdder_1500_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2322_io_a = FullAdder_1501_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2322_io_b = FullAdder_1502_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2322_io_ci = FullAdder_1503_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2323_io_a = FullAdder_1504_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2323_io_b = FullAdder_1505_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2323_io_ci = FullAdder_1506_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2324_io_a = FullAdder_1507_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2324_io_b = FullAdder_1508_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2324_io_ci = FullAdder_1509_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2325_io_a = FullAdder_1510_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2325_io_b = FullAdder_1511_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2325_io_ci = FullAdder_1512_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2326_io_a = FullAdder_1513_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2326_io_b = FullAdder_1514_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2326_io_ci = FullAdder_1515_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2327_io_a = FullAdder_300_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2327_io_b = FullAdder_1508_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2327_io_ci = FullAdder_1509_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2328_io_a = FullAdder_1510_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2328_io_b = FullAdder_1511_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2328_io_ci = FullAdder_1512_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2329_io_a = FullAdder_1513_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2329_io_b = FullAdder_1514_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2329_io_ci = FullAdder_1515_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2330_io_a = FullAdder_1516_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2330_io_b = FullAdder_1517_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2330_io_ci = FullAdder_1518_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2331_io_a = FullAdder_1519_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2331_io_b = FullAdder_1520_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2331_io_ci = FullAdder_1521_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2332_io_a = FullAdder_1522_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2332_io_b = FullAdder_1523_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2332_io_ci = FullAdder_1524_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2333_io_a = FullAdder_1517_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2333_io_b = FullAdder_1518_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2333_io_ci = FullAdder_1519_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2334_io_a = FullAdder_1520_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2334_io_b = FullAdder_1521_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2334_io_ci = FullAdder_1522_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2335_io_a = FullAdder_1523_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2335_io_b = FullAdder_1524_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2335_io_ci = FullAdder_1525_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2336_io_a = FullAdder_1526_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2336_io_b = FullAdder_1527_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2336_io_ci = FullAdder_1528_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2337_io_a = FullAdder_1529_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2337_io_b = FullAdder_1530_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2337_io_ci = FullAdder_1531_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2338_io_a = FullAdder_1532_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2338_io_b = FullAdder_1533_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2338_io_ci = FullAdder_1534_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_75_io_a = FullAdder_1535_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_75_io_b = FullAdder_1536_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2339_io_a = FullAdder_1527_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2339_io_b = FullAdder_1528_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2339_io_ci = FullAdder_1529_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2340_io_a = FullAdder_1530_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2340_io_b = FullAdder_1531_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2340_io_ci = FullAdder_1532_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2341_io_a = FullAdder_1533_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2341_io_b = FullAdder_1534_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2341_io_ci = FullAdder_1535_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2342_io_a = FullAdder_1536_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2342_io_b = FullAdder_1537_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2342_io_ci = FullAdder_1538_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2343_io_a = FullAdder_1539_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2343_io_b = FullAdder_1540_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2343_io_ci = FullAdder_1541_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2344_io_a = FullAdder_1542_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2344_io_b = FullAdder_1543_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2344_io_ci = FullAdder_1544_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_76_io_a = FullAdder_1545_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_76_io_b = FullAdder_1546_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2345_io_a = FullAdder_1537_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2345_io_b = FullAdder_1538_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2345_io_ci = FullAdder_1539_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2346_io_a = FullAdder_1540_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2346_io_b = FullAdder_1541_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2346_io_ci = FullAdder_1542_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2347_io_a = FullAdder_1543_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2347_io_b = FullAdder_1544_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2347_io_ci = FullAdder_1545_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2348_io_a = FullAdder_1546_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2348_io_b = FullAdder_1547_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2348_io_ci = FullAdder_1548_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2349_io_a = FullAdder_1549_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2349_io_b = FullAdder_1550_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2349_io_ci = FullAdder_1551_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2350_io_a = FullAdder_1552_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2350_io_b = FullAdder_1553_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2350_io_ci = FullAdder_1554_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2351_io_a = FullAdder_359_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2351_io_b = HalfAdder_12_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2351_io_ci = FullAdder_1547_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2352_io_a = FullAdder_1548_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2352_io_b = FullAdder_1549_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2352_io_ci = FullAdder_1550_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2353_io_a = FullAdder_1551_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2353_io_b = FullAdder_1552_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2353_io_ci = FullAdder_1553_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2354_io_a = FullAdder_1554_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2354_io_b = FullAdder_1555_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2354_io_ci = FullAdder_1556_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2355_io_a = FullAdder_1557_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2355_io_b = FullAdder_1558_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2355_io_ci = FullAdder_1559_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2356_io_a = FullAdder_1560_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2356_io_b = FullAdder_1561_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2356_io_ci = FullAdder_1562_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2357_io_a = FullAdder_1563_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2357_io_b = FullAdder_1564_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2357_io_ci = FullAdder_1565_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2358_io_a = FullAdder_374_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2358_io_b = FullAdder_375_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2358_io_ci = FullAdder_1557_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2359_io_a = FullAdder_1558_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2359_io_b = FullAdder_1559_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2359_io_ci = FullAdder_1560_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2360_io_a = FullAdder_1561_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2360_io_b = FullAdder_1562_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2360_io_ci = FullAdder_1563_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2361_io_a = FullAdder_1564_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2361_io_b = FullAdder_1565_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2361_io_ci = FullAdder_1566_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2362_io_a = FullAdder_1567_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2362_io_b = FullAdder_1568_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2362_io_ci = FullAdder_1569_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2363_io_a = FullAdder_1570_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2363_io_b = FullAdder_1571_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2363_io_ci = FullAdder_1572_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2364_io_a = FullAdder_1573_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2364_io_b = FullAdder_1574_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2364_io_ci = FullAdder_1575_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2365_io_a = FullAdder_1567_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2365_io_b = FullAdder_1568_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2365_io_ci = FullAdder_1569_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2366_io_a = FullAdder_1570_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2366_io_b = FullAdder_1571_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2366_io_ci = FullAdder_1572_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2367_io_a = FullAdder_1573_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2367_io_b = FullAdder_1574_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2367_io_ci = FullAdder_1575_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2368_io_a = FullAdder_1576_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2368_io_b = HalfAdder_46_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2368_io_ci = FullAdder_1577_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2369_io_a = FullAdder_1578_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2369_io_b = FullAdder_1579_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2369_io_ci = FullAdder_1580_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2370_io_a = FullAdder_1581_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2370_io_b = FullAdder_1582_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2370_io_ci = FullAdder_1583_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2371_io_a = FullAdder_1584_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2371_io_b = FullAdder_1585_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2371_io_ci = FullAdder_1586_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2372_io_a = HalfAdder_13_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2372_io_b = FullAdder_1577_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2372_io_ci = FullAdder_1578_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2373_io_a = FullAdder_1579_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2373_io_b = FullAdder_1580_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2373_io_ci = FullAdder_1581_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2374_io_a = FullAdder_1582_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2374_io_b = FullAdder_1583_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2374_io_ci = FullAdder_1584_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2375_io_a = FullAdder_1585_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2375_io_b = FullAdder_1586_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2375_io_ci = FullAdder_1587_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2376_io_a = FullAdder_1588_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2376_io_b = FullAdder_1589_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2376_io_ci = FullAdder_1590_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2377_io_a = FullAdder_1591_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2377_io_b = FullAdder_1592_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2377_io_ci = FullAdder_1593_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2378_io_a = FullAdder_1594_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2378_io_b = FullAdder_1595_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2378_io_ci = FullAdder_1596_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2379_io_a = FullAdder_424_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2379_io_b = FullAdder_1588_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2379_io_ci = FullAdder_1589_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2380_io_a = FullAdder_1590_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2380_io_b = FullAdder_1591_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2380_io_ci = FullAdder_1592_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2381_io_a = FullAdder_1593_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2381_io_b = FullAdder_1594_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2381_io_ci = FullAdder_1595_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2382_io_a = FullAdder_1596_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2382_io_b = FullAdder_1597_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2382_io_ci = FullAdder_1598_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2383_io_a = FullAdder_1599_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2383_io_b = FullAdder_1600_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2383_io_ci = FullAdder_1601_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2384_io_a = FullAdder_1602_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2384_io_b = FullAdder_1603_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2384_io_ci = FullAdder_1604_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2385_io_a = FullAdder_1605_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2385_io_b = FullAdder_1606_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2385_io_ci = FullAdder_1607_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_77_io_a = FullAdder_1608_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_77_io_b = FullAdder_1609_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2386_io_a = FullAdder_441_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2386_io_b = FullAdder_1599_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2386_io_ci = FullAdder_1600_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2387_io_a = FullAdder_1601_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2387_io_b = FullAdder_1602_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2387_io_ci = FullAdder_1603_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2388_io_a = FullAdder_1604_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2388_io_b = FullAdder_1605_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2388_io_ci = FullAdder_1606_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2389_io_a = FullAdder_1607_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2389_io_b = FullAdder_1608_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2389_io_ci = FullAdder_1609_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2390_io_a = FullAdder_1610_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2390_io_b = FullAdder_1611_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2390_io_ci = FullAdder_1612_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2391_io_a = FullAdder_1613_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2391_io_b = FullAdder_1614_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2391_io_ci = FullAdder_1615_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2392_io_a = FullAdder_1616_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2392_io_b = FullAdder_1617_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2392_io_ci = FullAdder_1618_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2393_io_a = FullAdder_1619_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2393_io_b = FullAdder_1620_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2393_io_ci = FullAdder_1621_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2394_io_a = FullAdder_1610_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2394_io_b = FullAdder_1611_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2394_io_ci = FullAdder_1612_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2395_io_a = FullAdder_1613_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2395_io_b = FullAdder_1614_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2395_io_ci = FullAdder_1615_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2396_io_a = FullAdder_1616_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2396_io_b = FullAdder_1617_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2396_io_ci = FullAdder_1618_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2397_io_a = FullAdder_1619_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2397_io_b = FullAdder_1620_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2397_io_ci = FullAdder_1621_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2398_io_a = FullAdder_1622_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2398_io_b = FullAdder_1623_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2398_io_ci = FullAdder_1624_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2399_io_a = FullAdder_1625_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2399_io_b = FullAdder_1626_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2399_io_ci = FullAdder_1627_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2400_io_a = FullAdder_1628_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2400_io_b = FullAdder_1629_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2400_io_ci = FullAdder_1630_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2401_io_a = FullAdder_1631_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2401_io_b = FullAdder_1632_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2401_io_ci = FullAdder_1633_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2402_io_a = FullAdder_1622_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2402_io_b = FullAdder_1623_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2402_io_ci = FullAdder_1624_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2403_io_a = FullAdder_1625_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2403_io_b = FullAdder_1626_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2403_io_ci = FullAdder_1627_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2404_io_a = FullAdder_1628_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2404_io_b = FullAdder_1629_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2404_io_ci = FullAdder_1630_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2405_io_a = FullAdder_1631_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2405_io_b = FullAdder_1632_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2405_io_ci = FullAdder_1633_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2406_io_a = FullAdder_1634_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2406_io_b = FullAdder_1635_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2406_io_ci = FullAdder_1636_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2407_io_a = FullAdder_1637_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2407_io_b = FullAdder_1638_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2407_io_ci = FullAdder_1639_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2408_io_a = FullAdder_1640_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2408_io_b = FullAdder_1641_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2408_io_ci = FullAdder_1642_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2409_io_a = FullAdder_1643_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2409_io_b = FullAdder_1644_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2409_io_ci = FullAdder_1645_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2410_io_a = FullAdder_1634_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2410_io_b = FullAdder_1635_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2410_io_ci = FullAdder_1636_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2411_io_a = FullAdder_1637_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2411_io_b = FullAdder_1638_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2411_io_ci = FullAdder_1639_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2412_io_a = FullAdder_1640_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2412_io_b = FullAdder_1641_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2412_io_ci = FullAdder_1642_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2413_io_a = FullAdder_1643_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2413_io_b = FullAdder_1644_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2413_io_ci = FullAdder_1645_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2414_io_a = FullAdder_1646_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2414_io_b = FullAdder_1647_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2414_io_ci = FullAdder_1648_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2415_io_a = FullAdder_1649_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2415_io_b = FullAdder_1650_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2415_io_ci = FullAdder_1651_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2416_io_a = FullAdder_1652_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2416_io_b = FullAdder_1653_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2416_io_ci = FullAdder_1654_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2417_io_a = FullAdder_1655_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2417_io_b = FullAdder_1656_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2417_io_ci = FullAdder_1657_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2418_io_a = FullAdder_1646_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2418_io_b = FullAdder_1647_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2418_io_ci = FullAdder_1648_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2419_io_a = FullAdder_1649_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2419_io_b = FullAdder_1650_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2419_io_ci = FullAdder_1651_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2420_io_a = FullAdder_1652_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2420_io_b = FullAdder_1653_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2420_io_ci = FullAdder_1654_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2421_io_a = FullAdder_1655_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2421_io_b = FullAdder_1656_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2421_io_ci = FullAdder_1657_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2422_io_a = HalfAdder_47_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2422_io_b = FullAdder_1658_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2422_io_ci = FullAdder_1659_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2423_io_a = FullAdder_1660_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2423_io_b = FullAdder_1661_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2423_io_ci = FullAdder_1662_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2424_io_a = FullAdder_1663_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2424_io_b = FullAdder_1664_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2424_io_ci = FullAdder_1665_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2425_io_a = FullAdder_1666_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2425_io_b = FullAdder_1667_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2425_io_ci = FullAdder_1668_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2426_io_a = FullAdder_1658_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2426_io_b = FullAdder_1659_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2426_io_ci = FullAdder_1660_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2427_io_a = FullAdder_1661_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2427_io_b = FullAdder_1662_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2427_io_ci = FullAdder_1663_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2428_io_a = FullAdder_1664_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2428_io_b = FullAdder_1665_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2428_io_ci = FullAdder_1666_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2429_io_a = FullAdder_1667_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2429_io_b = FullAdder_1668_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2429_io_ci = FullAdder_1669_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2430_io_a = HalfAdder_48_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2430_io_b = FullAdder_1670_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2430_io_ci = FullAdder_1671_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2431_io_a = FullAdder_1672_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2431_io_b = FullAdder_1673_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2431_io_ci = FullAdder_1674_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2432_io_a = FullAdder_1675_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2432_io_b = FullAdder_1676_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2432_io_ci = FullAdder_1677_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2433_io_a = FullAdder_1678_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2433_io_b = FullAdder_1679_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2433_io_ci = FullAdder_1680_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2434_io_a = FullAdder_549_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2434_io_b = FullAdder_550_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2434_io_ci = FullAdder_1670_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2435_io_a = FullAdder_1671_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2435_io_b = FullAdder_1672_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2435_io_ci = FullAdder_1673_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2436_io_a = FullAdder_1674_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2436_io_b = FullAdder_1675_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2436_io_ci = FullAdder_1676_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2437_io_a = FullAdder_1677_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2437_io_b = FullAdder_1678_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2437_io_ci = FullAdder_1679_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2438_io_a = FullAdder_1680_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2438_io_b = FullAdder_1681_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2438_io_ci = FullAdder_1682_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2439_io_a = FullAdder_1683_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2439_io_b = FullAdder_1684_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2439_io_ci = FullAdder_1685_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2440_io_a = FullAdder_1686_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2440_io_b = FullAdder_1687_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2440_io_ci = FullAdder_1688_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2441_io_a = FullAdder_1689_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2441_io_b = FullAdder_1690_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2441_io_ci = FullAdder_1691_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2442_io_a = FullAdder_1692_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2442_io_b = FullAdder_1693_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2442_io_ci = FullAdder_1694_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2443_io_a = HalfAdder_16_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2443_io_b = FullAdder_1682_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2443_io_ci = FullAdder_1683_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2444_io_a = FullAdder_1684_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2444_io_b = FullAdder_1685_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2444_io_ci = FullAdder_1686_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2445_io_a = FullAdder_1687_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2445_io_b = FullAdder_1688_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2445_io_ci = FullAdder_1689_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2446_io_a = FullAdder_1690_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2446_io_b = FullAdder_1691_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2446_io_ci = FullAdder_1692_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2447_io_a = FullAdder_1693_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2447_io_b = FullAdder_1694_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2447_io_ci = FullAdder_1695_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2448_io_a = FullAdder_1696_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2448_io_b = FullAdder_1697_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2448_io_ci = FullAdder_1698_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2449_io_a = FullAdder_1699_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2449_io_b = FullAdder_1700_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2449_io_ci = FullAdder_1701_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2450_io_a = FullAdder_1702_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2450_io_b = FullAdder_1703_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2450_io_ci = FullAdder_1704_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2451_io_a = FullAdder_1705_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2451_io_b = FullAdder_1706_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2451_io_ci = FullAdder_1707_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2452_io_a = FullAdder_589_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2452_io_b = FullAdder_1695_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2452_io_ci = FullAdder_1696_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2453_io_a = FullAdder_1697_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2453_io_b = FullAdder_1698_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2453_io_ci = FullAdder_1699_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2454_io_a = FullAdder_1700_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2454_io_b = FullAdder_1701_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2454_io_ci = FullAdder_1702_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2455_io_a = FullAdder_1703_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2455_io_b = FullAdder_1704_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2455_io_ci = FullAdder_1705_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2456_io_a = FullAdder_1706_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2456_io_b = FullAdder_1707_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2456_io_ci = FullAdder_1708_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2457_io_a = FullAdder_1709_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2457_io_b = FullAdder_1710_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2457_io_ci = FullAdder_1711_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2458_io_a = FullAdder_1712_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2458_io_b = FullAdder_1713_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2458_io_ci = FullAdder_1714_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2459_io_a = FullAdder_1715_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2459_io_b = FullAdder_1716_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2459_io_ci = FullAdder_1717_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2460_io_a = FullAdder_1718_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2460_io_b = FullAdder_1719_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2460_io_ci = FullAdder_1720_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2461_io_a = FullAdder_609_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2461_io_b = FullAdder_1708_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2461_io_ci = FullAdder_1709_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2462_io_a = FullAdder_1710_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2462_io_b = FullAdder_1711_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2462_io_ci = FullAdder_1712_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2463_io_a = FullAdder_1713_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2463_io_b = FullAdder_1714_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2463_io_ci = FullAdder_1715_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2464_io_a = FullAdder_1716_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2464_io_b = FullAdder_1717_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2464_io_ci = FullAdder_1718_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2465_io_a = FullAdder_1719_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2465_io_b = FullAdder_1720_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2465_io_ci = FullAdder_1721_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2466_io_a = FullAdder_1722_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2466_io_b = FullAdder_1723_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2466_io_ci = FullAdder_1724_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2467_io_a = FullAdder_1725_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2467_io_b = FullAdder_1726_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2467_io_ci = FullAdder_1727_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2468_io_a = FullAdder_1728_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2468_io_b = FullAdder_1729_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2468_io_ci = FullAdder_1730_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2469_io_a = FullAdder_1731_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2469_io_b = FullAdder_1732_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2469_io_ci = FullAdder_1733_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2470_io_a = FullAdder_1721_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2470_io_b = FullAdder_1722_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2470_io_ci = FullAdder_1723_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2471_io_a = FullAdder_1724_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2471_io_b = FullAdder_1725_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2471_io_ci = FullAdder_1726_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2472_io_a = FullAdder_1727_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2472_io_b = FullAdder_1728_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2472_io_ci = FullAdder_1729_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2473_io_a = FullAdder_1730_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2473_io_b = FullAdder_1731_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2473_io_ci = FullAdder_1732_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2474_io_a = FullAdder_1733_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2474_io_b = FullAdder_1734_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2474_io_ci = FullAdder_1735_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2475_io_a = FullAdder_1736_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2475_io_b = FullAdder_1737_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2475_io_ci = FullAdder_1738_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2476_io_a = FullAdder_1739_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2476_io_b = FullAdder_1740_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2476_io_ci = FullAdder_1741_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2477_io_a = FullAdder_1742_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2477_io_b = FullAdder_1743_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2477_io_ci = FullAdder_1744_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2478_io_a = FullAdder_1745_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2478_io_b = FullAdder_1746_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2478_io_ci = FullAdder_1747_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2479_io_a = FullAdder_1735_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2479_io_b = FullAdder_1736_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2479_io_ci = FullAdder_1737_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2480_io_a = FullAdder_1738_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2480_io_b = FullAdder_1739_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2480_io_ci = FullAdder_1740_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2481_io_a = FullAdder_1741_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2481_io_b = FullAdder_1742_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2481_io_ci = FullAdder_1743_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2482_io_a = FullAdder_1744_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2482_io_b = FullAdder_1745_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2482_io_ci = FullAdder_1746_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2483_io_a = FullAdder_1747_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2483_io_b = FullAdder_1748_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2483_io_ci = FullAdder_1749_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2484_io_a = FullAdder_1750_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2484_io_b = FullAdder_1751_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2484_io_ci = FullAdder_1752_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2485_io_a = FullAdder_1753_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2485_io_b = FullAdder_1754_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2485_io_ci = FullAdder_1755_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2486_io_a = FullAdder_1756_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2486_io_b = FullAdder_1757_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2486_io_ci = FullAdder_1758_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2487_io_a = FullAdder_1759_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2487_io_b = FullAdder_1760_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2487_io_ci = FullAdder_1761_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2488_io_a = FullAdder_1749_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2488_io_b = FullAdder_1750_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2488_io_ci = FullAdder_1751_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2489_io_a = FullAdder_1752_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2489_io_b = FullAdder_1753_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2489_io_ci = FullAdder_1754_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2490_io_a = FullAdder_1755_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2490_io_b = FullAdder_1756_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2490_io_ci = FullAdder_1757_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2491_io_a = FullAdder_1758_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2491_io_b = FullAdder_1759_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2491_io_ci = FullAdder_1760_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2492_io_a = FullAdder_1761_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2492_io_b = FullAdder_1762_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2492_io_ci = FullAdder_1763_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2493_io_a = FullAdder_1764_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2493_io_b = FullAdder_1765_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2493_io_ci = FullAdder_1766_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2494_io_a = FullAdder_1767_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2494_io_b = FullAdder_1768_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2494_io_ci = FullAdder_1769_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2495_io_a = FullAdder_1770_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2495_io_b = FullAdder_1771_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2495_io_ci = FullAdder_1772_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2496_io_a = FullAdder_1773_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2496_io_b = FullAdder_1774_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2496_io_ci = FullAdder_1775_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2497_io_a = FullAdder_692_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2497_io_b = FullAdder_1763_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2497_io_ci = FullAdder_1764_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2498_io_a = FullAdder_1765_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2498_io_b = FullAdder_1766_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2498_io_ci = FullAdder_1767_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2499_io_a = FullAdder_1768_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2499_io_b = FullAdder_1769_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2499_io_ci = FullAdder_1770_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2500_io_a = FullAdder_1771_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2500_io_b = FullAdder_1772_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2500_io_ci = FullAdder_1773_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2501_io_a = FullAdder_1774_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2501_io_b = FullAdder_1775_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2501_io_ci = FullAdder_1776_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2502_io_a = FullAdder_1777_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2502_io_b = FullAdder_1778_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2502_io_ci = FullAdder_1779_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2503_io_a = FullAdder_1780_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2503_io_b = FullAdder_1781_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2503_io_ci = FullAdder_1782_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2504_io_a = FullAdder_1783_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2504_io_b = FullAdder_1784_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2504_io_ci = FullAdder_1785_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2505_io_a = FullAdder_1786_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2505_io_b = FullAdder_1787_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2505_io_ci = FullAdder_1788_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_78_io_a = FullAdder_1789_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_78_io_b = FullAdder_1790_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2506_io_a = FullAdder_1777_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2506_io_b = FullAdder_1778_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2506_io_ci = FullAdder_1779_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2507_io_a = FullAdder_1780_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2507_io_b = FullAdder_1781_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2507_io_ci = FullAdder_1782_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2508_io_a = FullAdder_1783_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2508_io_b = FullAdder_1784_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2508_io_ci = FullAdder_1785_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2509_io_a = FullAdder_1786_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2509_io_b = FullAdder_1787_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2509_io_ci = FullAdder_1788_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2510_io_a = FullAdder_1789_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2510_io_b = FullAdder_1790_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2510_io_ci = FullAdder_1791_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2511_io_a = FullAdder_1792_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2511_io_b = FullAdder_1793_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2511_io_ci = FullAdder_1794_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2512_io_a = FullAdder_1795_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2512_io_b = FullAdder_1796_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2512_io_ci = FullAdder_1797_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2513_io_a = FullAdder_1798_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2513_io_b = FullAdder_1799_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2513_io_ci = FullAdder_1800_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2514_io_a = FullAdder_1801_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2514_io_b = FullAdder_1802_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2514_io_ci = FullAdder_1803_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2515_io_a = FullAdder_1791_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2515_io_b = FullAdder_1792_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2515_io_ci = FullAdder_1793_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2516_io_a = FullAdder_1794_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2516_io_b = FullAdder_1795_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2516_io_ci = FullAdder_1796_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2517_io_a = FullAdder_1797_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2517_io_b = FullAdder_1798_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2517_io_ci = FullAdder_1799_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2518_io_a = FullAdder_1800_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2518_io_b = FullAdder_1801_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2518_io_ci = FullAdder_1802_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2519_io_a = FullAdder_1803_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2519_io_b = HalfAdder_49_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2519_io_ci = FullAdder_1804_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2520_io_a = FullAdder_1805_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2520_io_b = FullAdder_1806_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2520_io_ci = FullAdder_1807_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2521_io_a = FullAdder_1808_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2521_io_b = FullAdder_1809_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2521_io_ci = FullAdder_1810_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2522_io_a = FullAdder_1811_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2522_io_b = FullAdder_1812_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2522_io_ci = FullAdder_1813_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2523_io_a = FullAdder_1814_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2523_io_b = FullAdder_1815_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2523_io_ci = FullAdder_1816_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2524_io_a = FullAdder_751_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2524_io_b = FullAdder_752_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2524_io_ci = FullAdder_1804_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2525_io_a = FullAdder_1805_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2525_io_b = FullAdder_1806_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2525_io_ci = FullAdder_1807_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2526_io_a = FullAdder_1808_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2526_io_b = FullAdder_1809_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2526_io_ci = FullAdder_1810_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2527_io_a = FullAdder_1811_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2527_io_b = FullAdder_1812_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2527_io_ci = FullAdder_1813_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2528_io_a = FullAdder_1814_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2528_io_b = FullAdder_1815_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2528_io_ci = FullAdder_1816_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2529_io_a = FullAdder_1817_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2529_io_b = FullAdder_1818_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2529_io_ci = FullAdder_1819_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2530_io_a = FullAdder_1820_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2530_io_b = FullAdder_1821_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2530_io_ci = FullAdder_1822_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2531_io_a = FullAdder_1823_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2531_io_b = FullAdder_1824_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2531_io_ci = FullAdder_1825_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2532_io_a = FullAdder_1826_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2532_io_b = FullAdder_1827_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2532_io_ci = FullAdder_1828_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2533_io_a = HalfAdder_19_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2533_io_b = FullAdder_1817_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2533_io_ci = FullAdder_1818_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2534_io_a = FullAdder_1819_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2534_io_b = FullAdder_1820_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2534_io_ci = FullAdder_1821_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2535_io_a = FullAdder_1822_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2535_io_b = FullAdder_1823_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2535_io_ci = FullAdder_1824_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2536_io_a = FullAdder_1825_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2536_io_b = FullAdder_1826_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2536_io_ci = FullAdder_1827_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2537_io_a = FullAdder_1828_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2537_io_b = FullAdder_1829_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2537_io_ci = FullAdder_1830_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2538_io_a = FullAdder_1831_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2538_io_b = FullAdder_1832_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2538_io_ci = FullAdder_1833_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2539_io_a = FullAdder_1834_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2539_io_b = FullAdder_1835_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2539_io_ci = FullAdder_1836_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2540_io_a = FullAdder_1837_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2540_io_b = FullAdder_1838_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2540_io_ci = FullAdder_1839_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2541_io_a = FullAdder_1840_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2541_io_b = FullAdder_1841_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2541_io_ci = FullAdder_1842_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2542_io_a = FullAdder_1830_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2542_io_b = FullAdder_1831_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2542_io_ci = FullAdder_1832_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2543_io_a = FullAdder_1833_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2543_io_b = FullAdder_1834_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2543_io_ci = FullAdder_1835_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2544_io_a = FullAdder_1836_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2544_io_b = FullAdder_1837_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2544_io_ci = FullAdder_1838_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2545_io_a = FullAdder_1839_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2545_io_b = FullAdder_1840_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2545_io_ci = FullAdder_1841_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2546_io_a = FullAdder_1842_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2546_io_b = FullAdder_1843_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2546_io_ci = FullAdder_1844_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2547_io_a = FullAdder_1845_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2547_io_b = FullAdder_1846_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2547_io_ci = FullAdder_1847_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2548_io_a = FullAdder_1848_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2548_io_b = FullAdder_1849_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2548_io_ci = FullAdder_1850_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2549_io_a = FullAdder_1851_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2549_io_b = FullAdder_1852_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2549_io_ci = FullAdder_1853_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_79_io_a = FullAdder_1854_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_79_io_b = FullAdder_1855_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2550_io_a = FullAdder_1843_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2550_io_b = FullAdder_1844_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2550_io_ci = FullAdder_1845_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2551_io_a = FullAdder_1846_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2551_io_b = FullAdder_1847_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2551_io_ci = FullAdder_1848_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2552_io_a = FullAdder_1849_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2552_io_b = FullAdder_1850_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2552_io_ci = FullAdder_1851_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2553_io_a = FullAdder_1852_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2553_io_b = FullAdder_1853_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2553_io_ci = FullAdder_1854_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2554_io_a = FullAdder_1855_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2554_io_b = FullAdder_1856_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2554_io_ci = FullAdder_1857_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2555_io_a = FullAdder_1858_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2555_io_b = FullAdder_1859_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2555_io_ci = FullAdder_1860_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2556_io_a = FullAdder_1861_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2556_io_b = FullAdder_1862_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2556_io_ci = FullAdder_1863_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2557_io_a = FullAdder_1864_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2557_io_b = FullAdder_1865_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2557_io_ci = FullAdder_1866_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2558_io_a = FullAdder_827_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2558_io_b = FullAdder_1856_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2558_io_ci = FullAdder_1857_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2559_io_a = FullAdder_1858_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2559_io_b = FullAdder_1859_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2559_io_ci = FullAdder_1860_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2560_io_a = FullAdder_1861_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2560_io_b = FullAdder_1862_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2560_io_ci = FullAdder_1863_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2561_io_a = FullAdder_1864_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2561_io_b = FullAdder_1865_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2561_io_ci = FullAdder_1866_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2562_io_a = FullAdder_1867_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2562_io_b = FullAdder_1868_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2562_io_ci = FullAdder_1869_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2563_io_a = FullAdder_1870_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2563_io_b = FullAdder_1871_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2563_io_ci = FullAdder_1872_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2564_io_a = FullAdder_1873_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2564_io_b = FullAdder_1874_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2564_io_ci = FullAdder_1875_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2565_io_a = FullAdder_1876_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2565_io_b = FullAdder_1877_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2565_io_ci = FullAdder_1878_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2566_io_a = FullAdder_844_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2566_io_b = FullAdder_845_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2566_io_ci = FullAdder_1868_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2567_io_a = FullAdder_1869_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2567_io_b = FullAdder_1870_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2567_io_ci = FullAdder_1871_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2568_io_a = FullAdder_1872_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2568_io_b = FullAdder_1873_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2568_io_ci = FullAdder_1874_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2569_io_a = FullAdder_1875_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2569_io_b = FullAdder_1876_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2569_io_ci = FullAdder_1877_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2570_io_a = FullAdder_1878_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2570_io_b = FullAdder_1879_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2570_io_ci = FullAdder_1880_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2571_io_a = FullAdder_1881_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2571_io_b = FullAdder_1882_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2571_io_ci = FullAdder_1883_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2572_io_a = FullAdder_1884_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2572_io_b = FullAdder_1885_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2572_io_ci = FullAdder_1886_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2573_io_a = FullAdder_1887_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2573_io_b = FullAdder_1888_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2573_io_ci = FullAdder_1889_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2574_io_a = FullAdder_863_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2574_io_b = FullAdder_1880_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2574_io_ci = FullAdder_1881_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2575_io_a = FullAdder_1882_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2575_io_b = FullAdder_1883_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2575_io_ci = FullAdder_1884_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2576_io_a = FullAdder_1885_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2576_io_b = FullAdder_1886_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2576_io_ci = FullAdder_1887_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2577_io_a = FullAdder_1888_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2577_io_b = FullAdder_1889_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2577_io_ci = FullAdder_1890_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2578_io_a = FullAdder_1891_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2578_io_b = FullAdder_1892_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2578_io_ci = FullAdder_1893_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2579_io_a = FullAdder_1894_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2579_io_b = FullAdder_1895_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2579_io_ci = FullAdder_1896_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2580_io_a = FullAdder_1897_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2580_io_b = FullAdder_1898_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2580_io_ci = FullAdder_1899_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2581_io_a = FullAdder_1900_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2581_io_b = FullAdder_1901_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2581_io_ci = FullAdder_1902_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2582_io_a = FullAdder_1892_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2582_io_b = FullAdder_1893_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2582_io_ci = FullAdder_1894_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2583_io_a = FullAdder_1895_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2583_io_b = FullAdder_1896_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2583_io_ci = FullAdder_1897_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2584_io_a = FullAdder_1898_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2584_io_b = FullAdder_1899_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2584_io_ci = FullAdder_1900_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2585_io_a = FullAdder_1901_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2585_io_b = FullAdder_1902_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2585_io_ci = FullAdder_1903_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2586_io_a = FullAdder_1904_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2586_io_b = FullAdder_1905_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2586_io_ci = FullAdder_1906_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2587_io_a = FullAdder_1907_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2587_io_b = FullAdder_1908_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2587_io_ci = FullAdder_1909_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2588_io_a = FullAdder_1910_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2588_io_b = FullAdder_1911_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2588_io_ci = FullAdder_1912_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2589_io_a = FullAdder_896_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2589_io_b = FullAdder_897_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2589_io_ci = FullAdder_1904_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2590_io_a = FullAdder_1905_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2590_io_b = FullAdder_1906_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2590_io_ci = FullAdder_1907_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2591_io_a = FullAdder_1908_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2591_io_b = FullAdder_1909_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2591_io_ci = FullAdder_1910_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2592_io_a = FullAdder_1911_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2592_io_b = FullAdder_1912_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2592_io_ci = FullAdder_1913_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2593_io_a = FullAdder_1914_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2593_io_b = FullAdder_1915_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2593_io_ci = FullAdder_1916_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2594_io_a = FullAdder_1917_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2594_io_b = FullAdder_1918_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2594_io_ci = FullAdder_1919_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2595_io_a = FullAdder_1920_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2595_io_b = FullAdder_1921_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2595_io_ci = FullAdder_1922_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2596_io_a = FullAdder_1923_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2596_io_b = FullAdder_1924_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2596_io_ci = FullAdder_1925_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2597_io_a = FullAdder_1915_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2597_io_b = FullAdder_1916_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2597_io_ci = FullAdder_1917_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2598_io_a = FullAdder_1918_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2598_io_b = FullAdder_1919_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2598_io_ci = FullAdder_1920_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2599_io_a = FullAdder_1921_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2599_io_b = FullAdder_1922_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2599_io_ci = FullAdder_1923_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2600_io_a = FullAdder_1924_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2600_io_b = FullAdder_1925_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2600_io_ci = HalfAdder_50_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2601_io_a = FullAdder_1926_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2601_io_b = FullAdder_1927_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2601_io_ci = FullAdder_1928_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2602_io_a = FullAdder_1929_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2602_io_b = FullAdder_1930_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2602_io_ci = FullAdder_1931_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2603_io_a = FullAdder_1932_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2603_io_b = FullAdder_1933_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2603_io_ci = FullAdder_1934_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_80_io_a = FullAdder_1935_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_80_io_b = FullAdder_1936_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2604_io_a = FullAdder_1926_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2604_io_b = FullAdder_1927_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2604_io_ci = FullAdder_1928_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2605_io_a = FullAdder_1929_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2605_io_b = FullAdder_1930_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2605_io_ci = FullAdder_1931_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2606_io_a = FullAdder_1932_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2606_io_b = FullAdder_1933_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2606_io_ci = FullAdder_1934_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2607_io_a = FullAdder_1935_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2607_io_b = FullAdder_1936_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2607_io_ci = FullAdder_1937_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2608_io_a = FullAdder_1938_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2608_io_b = FullAdder_1939_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2608_io_ci = FullAdder_1940_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2609_io_a = FullAdder_1941_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2609_io_b = FullAdder_1942_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2609_io_ci = FullAdder_1943_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2610_io_a = FullAdder_1944_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2610_io_b = FullAdder_1945_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2610_io_ci = FullAdder_1946_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2611_io_a = FullAdder_946_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2611_io_b = FullAdder_1937_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2611_io_ci = FullAdder_1938_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2612_io_a = FullAdder_1939_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2612_io_b = FullAdder_1940_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2612_io_ci = FullAdder_1941_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2613_io_a = FullAdder_1942_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2613_io_b = FullAdder_1943_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2613_io_ci = FullAdder_1944_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2614_io_a = FullAdder_1945_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2614_io_b = FullAdder_1946_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2614_io_ci = FullAdder_1947_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2615_io_a = FullAdder_1948_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2615_io_b = FullAdder_1949_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2615_io_ci = FullAdder_1950_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2616_io_a = FullAdder_1951_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2616_io_b = FullAdder_1952_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2616_io_ci = FullAdder_1953_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2617_io_a = FullAdder_1954_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2617_io_b = FullAdder_1955_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2617_io_ci = FullAdder_1956_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2618_io_a = FullAdder_1948_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2618_io_b = FullAdder_1949_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2618_io_ci = FullAdder_1950_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2619_io_a = FullAdder_1951_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2619_io_b = FullAdder_1952_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2619_io_ci = FullAdder_1953_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2620_io_a = FullAdder_1954_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2620_io_b = FullAdder_1955_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2620_io_ci = FullAdder_1956_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2621_io_a = FullAdder_1957_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2621_io_b = FullAdder_1958_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2621_io_ci = FullAdder_1959_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2622_io_a = FullAdder_1960_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2622_io_b = FullAdder_1961_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2622_io_ci = FullAdder_1962_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2623_io_a = FullAdder_1963_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2623_io_b = FullAdder_1964_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2623_io_ci = FullAdder_1965_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2624_io_a = FullAdder_1966_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2624_io_b = FullAdder_1967_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2624_io_ci = FullAdder_1968_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2625_io_a = FullAdder_1959_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2625_io_b = FullAdder_1960_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2625_io_ci = FullAdder_1961_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2626_io_a = FullAdder_1962_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2626_io_b = FullAdder_1963_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2626_io_ci = FullAdder_1964_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2627_io_a = FullAdder_1965_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2627_io_b = FullAdder_1966_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2627_io_ci = FullAdder_1967_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2628_io_a = FullAdder_1968_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2628_io_b = HalfAdder_51_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2628_io_ci = FullAdder_1969_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2629_io_a = FullAdder_1970_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2629_io_b = FullAdder_1971_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2629_io_ci = FullAdder_1972_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2630_io_a = FullAdder_1973_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2630_io_b = FullAdder_1974_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2630_io_ci = FullAdder_1975_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2631_io_a = FullAdder_1976_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2631_io_b = FullAdder_1977_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2631_io_ci = FullAdder_1978_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2632_io_a = FullAdder_992_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2632_io_b = FullAdder_1969_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2632_io_ci = FullAdder_1970_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2633_io_a = FullAdder_1971_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2633_io_b = FullAdder_1972_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2633_io_ci = FullAdder_1973_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2634_io_a = FullAdder_1974_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2634_io_b = FullAdder_1975_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2634_io_ci = FullAdder_1976_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2635_io_a = FullAdder_1977_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2635_io_b = FullAdder_1978_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2635_io_ci = FullAdder_1979_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2636_io_a = FullAdder_1980_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2636_io_b = FullAdder_1981_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2636_io_ci = FullAdder_1982_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2637_io_a = FullAdder_1983_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2637_io_b = FullAdder_1984_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2637_io_ci = FullAdder_1985_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2638_io_a = FullAdder_1986_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2638_io_b = FullAdder_1987_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2638_io_ci = FullAdder_1988_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2639_io_a = FullAdder_1007_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2639_io_b = FullAdder_1979_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2639_io_ci = FullAdder_1980_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2640_io_a = FullAdder_1981_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2640_io_b = FullAdder_1982_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2640_io_ci = FullAdder_1983_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2641_io_a = FullAdder_1984_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2641_io_b = FullAdder_1985_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2641_io_ci = FullAdder_1986_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2642_io_a = FullAdder_1987_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2642_io_b = FullAdder_1988_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2642_io_ci = FullAdder_1989_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2643_io_a = FullAdder_1990_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2643_io_b = FullAdder_1991_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2643_io_ci = FullAdder_1992_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2644_io_a = FullAdder_1993_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2644_io_b = FullAdder_1994_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2644_io_ci = FullAdder_1995_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_81_io_a = FullAdder_1996_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_81_io_b = FullAdder_1997_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2645_io_a = FullAdder_1020_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2645_io_b = FullAdder_1021_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2645_io_ci = FullAdder_1989_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2646_io_a = FullAdder_1990_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2646_io_b = FullAdder_1991_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2646_io_ci = FullAdder_1992_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2647_io_a = FullAdder_1993_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2647_io_b = FullAdder_1994_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2647_io_ci = FullAdder_1995_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2648_io_a = FullAdder_1996_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2648_io_b = FullAdder_1997_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2648_io_ci = FullAdder_1998_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2649_io_a = FullAdder_1999_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2649_io_b = FullAdder_2000_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2649_io_ci = FullAdder_2001_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2650_io_a = FullAdder_2002_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2650_io_b = FullAdder_2003_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2650_io_ci = FullAdder_2004_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2651_io_a = FullAdder_2005_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2651_io_b = FullAdder_2006_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2651_io_ci = FullAdder_2007_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2652_io_a = FullAdder_1998_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2652_io_b = FullAdder_1999_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2652_io_ci = FullAdder_2000_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2653_io_a = FullAdder_2001_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2653_io_b = FullAdder_2002_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2653_io_ci = FullAdder_2003_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2654_io_a = FullAdder_2004_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2654_io_b = FullAdder_2005_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2654_io_ci = FullAdder_2006_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2655_io_a = FullAdder_2007_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2655_io_b = FullAdder_2008_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2655_io_ci = FullAdder_2009_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2656_io_a = FullAdder_2010_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2656_io_b = FullAdder_2011_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2656_io_ci = FullAdder_2012_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2657_io_a = FullAdder_2013_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2657_io_b = FullAdder_2014_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2657_io_ci = FullAdder_2015_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2658_io_a = FullAdder_2008_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2658_io_b = FullAdder_2009_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2658_io_ci = FullAdder_2010_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2659_io_a = FullAdder_2011_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2659_io_b = FullAdder_2012_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2659_io_ci = FullAdder_2013_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2660_io_a = FullAdder_2014_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2660_io_b = FullAdder_2015_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2660_io_ci = FullAdder_2016_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2661_io_a = HalfAdder_52_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2661_io_b = FullAdder_2017_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2661_io_ci = FullAdder_2018_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2662_io_a = FullAdder_2019_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2662_io_b = FullAdder_2020_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2662_io_ci = FullAdder_2021_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2663_io_a = FullAdder_2022_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2663_io_b = FullAdder_2023_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2663_io_ci = FullAdder_2024_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2664_io_a = FullAdder_2017_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2664_io_b = FullAdder_2018_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2664_io_ci = FullAdder_2019_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2665_io_a = FullAdder_2020_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2665_io_b = FullAdder_2021_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2665_io_ci = FullAdder_2022_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2666_io_a = FullAdder_2023_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2666_io_b = FullAdder_2024_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2666_io_ci = FullAdder_2025_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2667_io_a = FullAdder_2026_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2667_io_b = FullAdder_2027_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2667_io_ci = FullAdder_2028_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2668_io_a = FullAdder_2029_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2668_io_b = FullAdder_2030_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2668_io_ci = FullAdder_2031_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2669_io_a = FullAdder_2032_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2669_io_b = FullAdder_2033_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2669_io_ci = FullAdder_2034_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2670_io_a = FullAdder_1075_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2670_io_b = FullAdder_2026_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2670_io_ci = FullAdder_2027_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2671_io_a = FullAdder_2028_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2671_io_b = FullAdder_2029_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2671_io_ci = FullAdder_2030_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2672_io_a = FullAdder_2031_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2672_io_b = FullAdder_2032_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2672_io_ci = FullAdder_2033_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2673_io_a = FullAdder_2034_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2673_io_b = FullAdder_2035_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2673_io_ci = FullAdder_2036_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2674_io_a = FullAdder_2037_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2674_io_b = FullAdder_2038_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2674_io_ci = FullAdder_2039_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2675_io_a = FullAdder_2040_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2675_io_b = FullAdder_2041_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2675_io_ci = FullAdder_2042_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2676_io_a = FullAdder_2035_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2676_io_b = FullAdder_2036_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2676_io_ci = FullAdder_2037_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2677_io_a = FullAdder_2038_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2677_io_b = FullAdder_2039_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2677_io_ci = FullAdder_2040_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2678_io_a = FullAdder_2041_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2678_io_b = FullAdder_2042_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2678_io_ci = FullAdder_2043_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2679_io_a = FullAdder_2044_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2679_io_b = FullAdder_2045_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2679_io_ci = FullAdder_2046_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2680_io_a = FullAdder_2047_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2680_io_b = FullAdder_2048_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2680_io_ci = FullAdder_2049_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2681_io_a = FullAdder_2050_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2681_io_b = FullAdder_2051_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2681_io_ci = HalfAdder_53_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2682_io_a = FullAdder_2044_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2682_io_b = FullAdder_2045_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2682_io_ci = FullAdder_2046_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2683_io_a = FullAdder_2047_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2683_io_b = FullAdder_2048_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2683_io_ci = FullAdder_2049_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2684_io_a = FullAdder_2050_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2684_io_b = FullAdder_2051_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2684_io_ci = HalfAdder_53_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2685_io_a = FullAdder_2052_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2685_io_b = FullAdder_2053_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2685_io_ci = FullAdder_2054_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2686_io_a = FullAdder_2055_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2686_io_b = FullAdder_2056_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2686_io_ci = FullAdder_2057_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2687_io_a = FullAdder_1112_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2687_io_b = FullAdder_2052_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2687_io_ci = FullAdder_2053_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2688_io_a = FullAdder_2054_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2688_io_b = FullAdder_2055_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2688_io_ci = FullAdder_2056_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2689_io_a = FullAdder_2057_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2689_io_b = FullAdder_2058_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2689_io_ci = FullAdder_2059_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2690_io_a = FullAdder_2060_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2690_io_b = FullAdder_2061_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2690_io_ci = FullAdder_2062_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2691_io_a = FullAdder_2063_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2691_io_b = FullAdder_2064_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2691_io_ci = FullAdder_2065_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_82_io_a = FullAdder_2066_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_82_io_b = FullAdder_2067_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2692_io_a = FullAdder_1124_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2692_io_b = FullAdder_2060_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2692_io_ci = FullAdder_2061_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2693_io_a = FullAdder_2062_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2693_io_b = FullAdder_2063_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2693_io_ci = FullAdder_2064_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2694_io_a = FullAdder_2065_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2694_io_b = FullAdder_2066_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2694_io_ci = FullAdder_2067_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2695_io_a = FullAdder_2068_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2695_io_b = FullAdder_2069_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2695_io_ci = FullAdder_2070_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2696_io_a = FullAdder_2071_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2696_io_b = FullAdder_2072_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2696_io_ci = FullAdder_2073_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_83_io_a = FullAdder_2074_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_83_io_b = FullAdder_2075_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2697_io_a = FullAdder_2068_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2697_io_b = FullAdder_2069_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2697_io_ci = FullAdder_2070_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2698_io_a = FullAdder_2071_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2698_io_b = FullAdder_2072_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2698_io_ci = FullAdder_2073_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2699_io_a = FullAdder_2074_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2699_io_b = FullAdder_2075_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2699_io_ci = FullAdder_2076_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2700_io_a = FullAdder_2077_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2700_io_b = FullAdder_2078_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2700_io_ci = FullAdder_2079_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2701_io_a = FullAdder_2080_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2701_io_b = FullAdder_2081_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2701_io_ci = FullAdder_2082_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2702_io_a = FullAdder_1145_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2702_io_b = FullAdder_1146_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2702_io_ci = FullAdder_2076_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2703_io_a = FullAdder_2077_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2703_io_b = FullAdder_2078_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2703_io_ci = FullAdder_2079_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2704_io_a = FullAdder_2080_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2704_io_b = FullAdder_2081_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2704_io_ci = FullAdder_2082_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2705_io_a = FullAdder_2083_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2705_io_b = FullAdder_2084_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2705_io_ci = FullAdder_2085_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2706_io_a = FullAdder_2086_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2706_io_b = FullAdder_2087_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2706_io_ci = FullAdder_2088_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2707_io_a = FullAdder_2083_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2707_io_b = FullAdder_2084_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2707_io_ci = FullAdder_2085_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2708_io_a = FullAdder_2086_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2708_io_b = FullAdder_2087_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2708_io_ci = FullAdder_2088_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2709_io_a = FullAdder_2089_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2709_io_b = HalfAdder_54_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2709_io_ci = FullAdder_2090_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2710_io_a = FullAdder_2091_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2710_io_b = FullAdder_2092_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2710_io_ci = FullAdder_2093_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2711_io_a = FullAdder_2094_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2711_io_b = FullAdder_2095_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2711_io_ci = FullAdder_2096_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2712_io_a = HalfAdder_24_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2712_io_b = FullAdder_2090_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2712_io_ci = FullAdder_2091_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2713_io_a = FullAdder_2092_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2713_io_b = FullAdder_2093_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2713_io_ci = FullAdder_2094_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2714_io_a = FullAdder_2095_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2714_io_b = FullAdder_2096_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2714_io_ci = FullAdder_2097_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2715_io_a = FullAdder_2098_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2715_io_b = FullAdder_2099_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2715_io_ci = FullAdder_2100_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2716_io_a = FullAdder_2101_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2716_io_b = FullAdder_2102_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2716_io_ci = FullAdder_2103_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2717_io_a = FullAdder_2097_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2717_io_b = FullAdder_2098_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2717_io_ci = FullAdder_2099_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2718_io_a = FullAdder_2100_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2718_io_b = FullAdder_2101_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2718_io_ci = FullAdder_2102_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2719_io_a = FullAdder_2103_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2719_io_b = FullAdder_2104_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2719_io_ci = FullAdder_2105_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2720_io_a = FullAdder_2106_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2720_io_b = FullAdder_2107_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2720_io_ci = FullAdder_2108_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2721_io_a = FullAdder_2104_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2721_io_b = FullAdder_2105_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2721_io_ci = FullAdder_2106_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2722_io_a = FullAdder_2107_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2722_io_b = FullAdder_2108_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2722_io_ci = FullAdder_2109_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2723_io_a = FullAdder_2110_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2723_io_b = FullAdder_2111_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2723_io_ci = FullAdder_2112_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2724_io_a = FullAdder_2113_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2724_io_b = FullAdder_2114_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2724_io_ci = FullAdder_2115_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_84_io_a = FullAdder_2116_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_84_io_b = HalfAdder_55_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2725_io_a = FullAdder_2111_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2725_io_b = FullAdder_2112_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2725_io_ci = FullAdder_2113_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2726_io_a = FullAdder_2114_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2726_io_b = FullAdder_2115_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2726_io_ci = FullAdder_2116_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2727_io_a = HalfAdder_55_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2727_io_b = FullAdder_2117_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2727_io_ci = FullAdder_2118_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2728_io_a = FullAdder_2119_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2728_io_b = FullAdder_2120_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2728_io_ci = FullAdder_2121_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2729_io_a = FullAdder_1205_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2729_io_b = FullAdder_2117_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2729_io_ci = FullAdder_2118_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2730_io_a = FullAdder_2119_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2730_io_b = FullAdder_2120_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2730_io_ci = FullAdder_2121_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2731_io_a = FullAdder_2122_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2731_io_b = FullAdder_2123_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2731_io_ci = FullAdder_2124_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2732_io_a = FullAdder_2125_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2732_io_b = FullAdder_2126_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2732_io_ci = FullAdder_2127_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2733_io_a = FullAdder_1214_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2733_io_b = FullAdder_2123_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2733_io_ci = FullAdder_2124_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2734_io_a = FullAdder_2125_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2734_io_b = FullAdder_2126_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2734_io_ci = FullAdder_2127_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2735_io_a = FullAdder_2128_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2735_io_b = FullAdder_2129_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2735_io_ci = FullAdder_2130_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2736_io_a = FullAdder_2131_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2736_io_b = FullAdder_2132_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2736_io_ci = FullAdder_2133_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2737_io_a = FullAdder_2129_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2737_io_b = FullAdder_2130_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2737_io_ci = FullAdder_2131_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2738_io_a = FullAdder_2132_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2738_io_b = FullAdder_2133_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2738_io_ci = HalfAdder_56_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2739_io_a = FullAdder_2134_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2739_io_b = FullAdder_2135_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2739_io_ci = FullAdder_2136_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2740_io_a = FullAdder_2137_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2740_io_b = FullAdder_2138_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2740_io_ci = FullAdder_2139_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2741_io_a = FullAdder_2134_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2741_io_b = FullAdder_2135_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2741_io_ci = FullAdder_2136_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2742_io_a = FullAdder_2137_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2742_io_b = FullAdder_2138_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2742_io_ci = FullAdder_2139_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2743_io_a = FullAdder_2140_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2743_io_b = FullAdder_2141_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2743_io_ci = FullAdder_2142_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2744_io_a = FullAdder_1237_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2744_io_b = FullAdder_1238_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2744_io_ci = FullAdder_2140_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2745_io_a = FullAdder_2141_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2745_io_b = FullAdder_2142_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2745_io_ci = FullAdder_2143_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2746_io_a = FullAdder_2144_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2746_io_b = FullAdder_2145_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2746_io_ci = FullAdder_2146_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2747_io_a = FullAdder_2147_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2747_io_b = FullAdder_2148_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2747_io_ci = FullAdder_2149_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2748_io_a = HalfAdder_26_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2748_io_b = FullAdder_2145_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2748_io_ci = FullAdder_2146_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2749_io_a = FullAdder_2147_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2749_io_b = FullAdder_2148_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2749_io_ci = FullAdder_2149_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2750_io_a = FullAdder_2150_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2750_io_b = FullAdder_2151_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2750_io_ci = FullAdder_2152_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_85_io_a = FullAdder_2153_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_85_io_b = FullAdder_2154_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2751_io_a = FullAdder_2150_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2751_io_b = FullAdder_2151_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2751_io_ci = FullAdder_2152_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2752_io_a = FullAdder_2153_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2752_io_b = FullAdder_2154_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2752_io_ci = FullAdder_2155_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2753_io_a = FullAdder_2156_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2753_io_b = FullAdder_2157_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2753_io_ci = FullAdder_2158_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2754_io_a = FullAdder_2155_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2754_io_b = FullAdder_2156_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2754_io_ci = FullAdder_2157_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2755_io_a = FullAdder_2158_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2755_io_b = FullAdder_2159_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2755_io_ci = FullAdder_2160_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2756_io_a = FullAdder_2161_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2756_io_b = FullAdder_2162_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2756_io_ci = FullAdder_2163_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2757_io_a = FullAdder_2160_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2757_io_b = FullAdder_2161_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2757_io_ci = FullAdder_2162_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2758_io_a = FullAdder_2163_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2758_io_b = HalfAdder_57_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2758_io_ci = FullAdder_2164_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2759_io_a = FullAdder_2165_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2759_io_b = FullAdder_2166_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2759_io_ci = FullAdder_2167_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2760_io_a = FullAdder_1271_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2760_io_b = FullAdder_2164_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2760_io_ci = FullAdder_2165_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2761_io_a = FullAdder_2166_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2761_io_b = FullAdder_2167_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2761_io_ci = FullAdder_2168_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2762_io_a = FullAdder_2169_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2762_io_b = FullAdder_2170_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2762_io_ci = FullAdder_2171_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2763_io_a = FullAdder_1277_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2763_io_b = FullAdder_2168_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2763_io_ci = FullAdder_2169_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2764_io_a = FullAdder_2170_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2764_io_b = FullAdder_2171_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2764_io_ci = FullAdder_2172_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2765_io_a = FullAdder_2173_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2765_io_b = FullAdder_2174_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2765_io_ci = FullAdder_2175_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2766_io_a = FullAdder_2172_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2766_io_b = FullAdder_2173_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2766_io_ci = FullAdder_2174_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2767_io_a = FullAdder_2175_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2767_io_b = FullAdder_2176_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2767_io_ci = FullAdder_2177_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2768_io_a = FullAdder_2176_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2768_io_b = FullAdder_2177_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2768_io_ci = FullAdder_2178_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2769_io_a = HalfAdder_58_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2769_io_b = FullAdder_2179_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2769_io_ci = FullAdder_2180_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_86_io_a = FullAdder_2181_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_86_io_b = HalfAdder_59_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2770_io_a = FullAdder_2179_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2770_io_b = FullAdder_2180_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2770_io_ci = FullAdder_2181_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2771_io_a = HalfAdder_59_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2771_io_b = FullAdder_2182_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2771_io_ci = FullAdder_2183_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2772_io_a = HalfAdder_29_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2772_io_b = FullAdder_2182_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2772_io_ci = FullAdder_2183_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2773_io_a = FullAdder_2184_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2773_io_b = FullAdder_2185_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2773_io_ci = FullAdder_2186_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2774_io_a = FullAdder_2185_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2774_io_b = FullAdder_2186_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2774_io_ci = FullAdder_2187_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2775_io_a = FullAdder_2188_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2775_io_b = FullAdder_2189_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2775_io_ci = FullAdder_2190_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2776_io_a = FullAdder_2188_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2776_io_b = FullAdder_2189_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2776_io_ci = FullAdder_2190_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2777_io_a = FullAdder_1307_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2777_io_b = HalfAdder_30_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2777_io_ci = FullAdder_2191_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2778_io_a = FullAdder_2192_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2778_io_b = FullAdder_2193_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2778_io_ci = HalfAdder_60_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_87_io_a = FullAdder_2193_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_87_io_b = HalfAdder_60_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_88_io_a = HalfAdder_61_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_88_io_b = FullAdder_2194_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2779_io_a = FullAdder_1313_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2779_io_b = FullAdder_2194_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2779_io_ci = FullAdder_2195_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_89_io_a = FullAdder_2196_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_89_io_b = FullAdder_2197_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2780_io_a = FullAdder_2196_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2780_io_b = FullAdder_2197_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2780_io_ci = FullAdder_2198_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2781_io_a = FullAdder_2198_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2781_io_b = HalfAdder_62_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2781_io_ci = FullAdder_2199_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2782_io_a = FullAdder_2199_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2782_io_b = HalfAdder_63_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2782_io_ci = FullAdder_2200_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2783_io_a = HalfAdder_32_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2783_io_b = FullAdder_2200_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2783_io_ci = HalfAdder_64_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_90_io_a = FullAdder_1321_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_90_io_b = HalfAdder_64_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_91_io_a = FullAdder_2201_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_91_io_b = HalfAdder_65_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_92_io_a = HalfAdder_66_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_92_io_b = HalfAdder_67_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_93_io_a = HalfAdder_67_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_93_io_b = HalfAdder_68_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_94_io_a = FullAdder_1323_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_94_io_b = HalfAdder_69_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_95_io_a = FullAdder_2202_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_95_io_b = FullAdder_2203_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2784_io_a = FullAdder_1326_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2784_io_b = FullAdder_2203_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2784_io_ci = HalfAdder_70_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_96_io_a = HalfAdder_70_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_96_io_b = HalfAdder_71_io_s; // @[wallace.scala 60:18]
  assign FullAdder_2785_io_a = FullAdder_1330_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2785_io_b = FullAdder_2204_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2785_io_ci = FullAdder_2205_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2786_io_a = FullAdder_1332_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2786_io_b = FullAdder_2205_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2786_io_ci = FullAdder_2206_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2787_io_a = HalfAdder_37_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2787_io_b = FullAdder_2206_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2787_io_ci = FullAdder_2207_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2788_io_a = FullAdder_2208_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2788_io_b = FullAdder_2209_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2788_io_ci = FullAdder_2210_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2789_io_a = FullAdder_2210_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2789_io_b = FullAdder_2211_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2789_io_ci = FullAdder_2212_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2790_io_a = FullAdder_2212_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2790_io_b = FullAdder_2213_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2790_io_ci = FullAdder_2214_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2791_io_a = FullAdder_1344_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2791_io_b = FullAdder_1345_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2791_io_ci = FullAdder_2214_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2792_io_a = FullAdder_2215_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2792_io_b = FullAdder_2216_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2792_io_ci = FullAdder_2217_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2793_io_a = FullAdder_2216_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2793_io_b = FullAdder_2217_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2793_io_ci = HalfAdder_72_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2794_io_a = FullAdder_1352_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2794_io_b = FullAdder_1353_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2794_io_ci = FullAdder_2218_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2795_io_a = FullAdder_2219_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2795_io_b = FullAdder_2220_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2795_io_ci = FullAdder_2221_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2796_io_a = FullAdder_2220_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2796_io_b = FullAdder_2221_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2796_io_ci = HalfAdder_73_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2797_io_a = FullAdder_2222_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2797_io_b = FullAdder_2223_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2797_io_ci = FullAdder_2224_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2798_io_a = FullAdder_2222_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2798_io_b = FullAdder_2223_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2798_io_ci = FullAdder_2224_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2799_io_a = FullAdder_2225_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2799_io_b = FullAdder_2226_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2799_io_ci = FullAdder_2227_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2800_io_a = HalfAdder_40_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2800_io_b = FullAdder_2225_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2800_io_ci = FullAdder_2226_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2801_io_a = FullAdder_2227_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2801_io_b = FullAdder_2228_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2801_io_ci = FullAdder_2229_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2802_io_a = HalfAdder_41_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2802_io_b = FullAdder_2228_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2802_io_ci = FullAdder_2229_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2803_io_a = FullAdder_2230_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2803_io_b = FullAdder_2231_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2803_io_ci = FullAdder_2232_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2804_io_a = FullAdder_1374_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2804_io_b = FullAdder_2231_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2804_io_ci = FullAdder_2232_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2805_io_a = FullAdder_2233_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2805_io_b = FullAdder_2234_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2805_io_ci = FullAdder_2235_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2806_io_a = FullAdder_1378_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2806_io_b = FullAdder_1379_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2806_io_ci = FullAdder_2234_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2807_io_a = FullAdder_2235_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2807_io_b = FullAdder_2236_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2807_io_ci = FullAdder_2237_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2808_io_a = FullAdder_2238_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2808_io_b = FullAdder_2239_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2808_io_ci = HalfAdder_74_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2809_io_a = FullAdder_2237_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2809_io_b = FullAdder_2238_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2809_io_ci = FullAdder_2239_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2810_io_a = HalfAdder_74_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2810_io_b = FullAdder_2240_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2810_io_ci = FullAdder_2241_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2811_io_a = FullAdder_1388_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2811_io_b = FullAdder_1389_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2811_io_ci = FullAdder_2240_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2812_io_a = FullAdder_2241_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2812_io_b = FullAdder_2242_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2812_io_ci = FullAdder_2243_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2813_io_a = FullAdder_2244_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2813_io_b = FullAdder_2245_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2813_io_ci = FullAdder_2246_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2814_io_a = FullAdder_1395_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2814_io_b = FullAdder_2243_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2814_io_ci = FullAdder_2244_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2815_io_a = FullAdder_2245_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2815_io_b = FullAdder_2246_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2815_io_ci = FullAdder_2247_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2816_io_a = FullAdder_2248_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2816_io_b = FullAdder_2249_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2816_io_ci = FullAdder_2250_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2817_io_a = FullAdder_1401_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2817_io_b = FullAdder_2247_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2817_io_ci = FullAdder_2248_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2818_io_a = FullAdder_2249_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2818_io_b = FullAdder_2250_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2818_io_ci = FullAdder_2251_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2819_io_a = FullAdder_2252_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2819_io_b = FullAdder_2253_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2819_io_ci = FullAdder_2254_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2820_io_a = FullAdder_2251_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2820_io_b = FullAdder_2252_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2820_io_ci = FullAdder_2253_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2821_io_a = FullAdder_2254_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2821_io_b = FullAdder_2255_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2821_io_ci = FullAdder_2256_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_97_io_a = FullAdder_2257_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_97_io_b = FullAdder_2258_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2822_io_a = FullAdder_1413_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2822_io_b = FullAdder_1414_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2822_io_ci = FullAdder_2255_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2823_io_a = FullAdder_2256_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2823_io_b = FullAdder_2257_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2823_io_ci = FullAdder_2258_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2824_io_a = FullAdder_2259_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2824_io_b = FullAdder_2260_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2824_io_ci = FullAdder_2261_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2825_io_a = FullAdder_1420_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2825_io_b = HalfAdder_42_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2825_io_ci = FullAdder_2259_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2826_io_a = FullAdder_2260_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2826_io_b = FullAdder_2261_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2826_io_ci = FullAdder_2262_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2827_io_a = FullAdder_2263_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2827_io_b = FullAdder_2264_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2827_io_ci = FullAdder_2265_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2828_io_a = FullAdder_1426_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2828_io_b = FullAdder_1427_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2828_io_ci = FullAdder_2263_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2829_io_a = FullAdder_2264_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2829_io_b = FullAdder_2265_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2829_io_ci = FullAdder_2266_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2830_io_a = FullAdder_2267_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2830_io_b = FullAdder_2268_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2830_io_ci = FullAdder_2269_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2831_io_a = FullAdder_2267_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2831_io_b = FullAdder_2268_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2831_io_ci = FullAdder_2269_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2832_io_a = FullAdder_2270_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2832_io_b = FullAdder_2271_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2832_io_ci = FullAdder_2272_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2833_io_a = FullAdder_2273_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2833_io_b = FullAdder_2274_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2833_io_ci = FullAdder_2275_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2834_io_a = FullAdder_2272_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2834_io_b = FullAdder_2273_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2834_io_ci = FullAdder_2274_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2835_io_a = FullAdder_2275_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2835_io_b = FullAdder_2276_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2835_io_ci = FullAdder_2277_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2836_io_a = FullAdder_2278_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2836_io_b = FullAdder_2279_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2836_io_ci = FullAdder_2280_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2837_io_a = FullAdder_1449_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2837_io_b = FullAdder_2277_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2837_io_ci = FullAdder_2278_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2838_io_a = FullAdder_2279_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2838_io_b = FullAdder_2280_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2838_io_ci = FullAdder_2281_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2839_io_a = FullAdder_2282_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2839_io_b = FullAdder_2283_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2839_io_ci = FullAdder_2284_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_98_io_a = FullAdder_2285_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_98_io_b = FullAdder_2286_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2840_io_a = FullAdder_1457_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2840_io_b = FullAdder_2282_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2840_io_ci = FullAdder_2283_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2841_io_a = FullAdder_2284_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2841_io_b = FullAdder_2285_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2841_io_ci = FullAdder_2286_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2842_io_a = FullAdder_2287_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2842_io_b = FullAdder_2288_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2842_io_ci = FullAdder_2289_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_99_io_a = FullAdder_2290_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_99_io_b = FullAdder_2291_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2843_io_a = FullAdder_1465_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2843_io_b = FullAdder_2287_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2843_io_ci = FullAdder_2288_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2844_io_a = FullAdder_2289_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2844_io_b = FullAdder_2290_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2844_io_ci = FullAdder_2291_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2845_io_a = FullAdder_2292_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2845_io_b = FullAdder_2293_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2845_io_ci = FullAdder_2294_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_100_io_a = FullAdder_2295_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_100_io_b = FullAdder_2296_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2846_io_a = FullAdder_1473_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2846_io_b = HalfAdder_43_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2846_io_ci = FullAdder_2292_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2847_io_a = FullAdder_2293_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2847_io_b = FullAdder_2294_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2847_io_ci = FullAdder_2295_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2848_io_a = FullAdder_2296_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2848_io_b = FullAdder_2297_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2848_io_ci = FullAdder_2298_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2849_io_a = FullAdder_2299_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2849_io_b = FullAdder_2300_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2849_io_ci = FullAdder_2301_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2850_io_a = FullAdder_2297_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2850_io_b = FullAdder_2298_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2850_io_ci = FullAdder_2299_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2851_io_a = FullAdder_2300_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2851_io_b = FullAdder_2301_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2851_io_ci = FullAdder_2302_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2852_io_a = FullAdder_2303_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2852_io_b = FullAdder_2304_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2852_io_ci = FullAdder_2305_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2853_io_a = FullAdder_2306_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2853_io_b = FullAdder_2307_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2853_io_ci = FullAdder_2308_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2854_io_a = FullAdder_2303_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2854_io_b = FullAdder_2304_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2854_io_ci = FullAdder_2305_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2855_io_a = FullAdder_2306_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2855_io_b = FullAdder_2307_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2855_io_ci = FullAdder_2308_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2856_io_a = FullAdder_2309_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2856_io_b = FullAdder_2310_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2856_io_ci = FullAdder_2311_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2857_io_a = FullAdder_2312_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2857_io_b = FullAdder_2313_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2857_io_ci = FullAdder_2314_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2858_io_a = FullAdder_2309_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2858_io_b = FullAdder_2310_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2858_io_ci = FullAdder_2311_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2859_io_a = FullAdder_2312_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2859_io_b = FullAdder_2313_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2859_io_ci = FullAdder_2314_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2860_io_a = FullAdder_2315_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2860_io_b = FullAdder_2316_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2860_io_ci = FullAdder_2317_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2861_io_a = FullAdder_2318_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2861_io_b = FullAdder_2319_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2861_io_ci = FullAdder_2320_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2862_io_a = FullAdder_1507_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2862_io_b = FullAdder_2315_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2862_io_ci = FullAdder_2316_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2863_io_a = FullAdder_2317_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2863_io_b = FullAdder_2318_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2863_io_ci = FullAdder_2319_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2864_io_a = FullAdder_2320_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2864_io_b = FullAdder_2321_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2864_io_ci = FullAdder_2322_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2865_io_a = FullAdder_2323_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2865_io_b = FullAdder_2324_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2865_io_ci = FullAdder_2325_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2866_io_a = FullAdder_1516_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2866_io_b = FullAdder_2321_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2866_io_ci = FullAdder_2322_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2867_io_a = FullAdder_2323_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2867_io_b = FullAdder_2324_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2867_io_ci = FullAdder_2325_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2868_io_a = FullAdder_2326_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2868_io_b = FullAdder_2327_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2868_io_ci = FullAdder_2328_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2869_io_a = FullAdder_2329_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2869_io_b = FullAdder_2330_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2869_io_ci = FullAdder_2331_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2870_io_a = FullAdder_1525_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2870_io_b = FullAdder_1526_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2870_io_ci = FullAdder_2327_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2871_io_a = FullAdder_2328_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2871_io_b = FullAdder_2329_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2871_io_ci = FullAdder_2330_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2872_io_a = FullAdder_2331_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2872_io_b = FullAdder_2332_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2872_io_ci = FullAdder_2333_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2873_io_a = FullAdder_2334_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2873_io_b = FullAdder_2335_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2873_io_ci = FullAdder_2336_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2874_io_a = FullAdder_2337_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2874_io_b = FullAdder_2338_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2874_io_ci = HalfAdder_75_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2875_io_a = FullAdder_2333_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2875_io_b = FullAdder_2334_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2875_io_ci = FullAdder_2335_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2876_io_a = FullAdder_2336_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2876_io_b = FullAdder_2337_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2876_io_ci = FullAdder_2338_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2877_io_a = HalfAdder_75_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2877_io_b = FullAdder_2339_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2877_io_ci = FullAdder_2340_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2878_io_a = FullAdder_2341_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2878_io_b = FullAdder_2342_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2878_io_ci = FullAdder_2343_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_101_io_a = FullAdder_2344_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_101_io_b = HalfAdder_76_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2879_io_a = FullAdder_2339_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2879_io_b = FullAdder_2340_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2879_io_ci = FullAdder_2341_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2880_io_a = FullAdder_2342_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2880_io_b = FullAdder_2343_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2880_io_ci = FullAdder_2344_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2881_io_a = HalfAdder_76_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2881_io_b = FullAdder_2345_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2881_io_ci = FullAdder_2346_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2882_io_a = FullAdder_2347_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2882_io_b = FullAdder_2348_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2882_io_ci = FullAdder_2349_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2883_io_a = FullAdder_1555_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2883_io_b = FullAdder_1556_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2883_io_ci = FullAdder_2345_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2884_io_a = FullAdder_2346_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2884_io_b = FullAdder_2347_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2884_io_ci = FullAdder_2348_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2885_io_a = FullAdder_2349_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2885_io_b = FullAdder_2350_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2885_io_ci = FullAdder_2351_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2886_io_a = FullAdder_2352_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2886_io_b = FullAdder_2353_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2886_io_ci = FullAdder_2354_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2887_io_a = FullAdder_2355_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2887_io_b = FullAdder_2356_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2887_io_ci = FullAdder_2357_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2888_io_a = FullAdder_1566_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2888_io_b = FullAdder_2351_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2888_io_ci = FullAdder_2352_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2889_io_a = FullAdder_2353_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2889_io_b = FullAdder_2354_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2889_io_ci = FullAdder_2355_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2890_io_a = FullAdder_2356_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2890_io_b = FullAdder_2357_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2890_io_ci = FullAdder_2358_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2891_io_a = FullAdder_2359_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2891_io_b = FullAdder_2360_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2891_io_ci = FullAdder_2361_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2892_io_a = FullAdder_2362_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2892_io_b = FullAdder_2363_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2892_io_ci = FullAdder_2364_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2893_io_a = FullAdder_1576_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2893_io_b = HalfAdder_46_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2893_io_ci = FullAdder_2358_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2894_io_a = FullAdder_2359_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2894_io_b = FullAdder_2360_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2894_io_ci = FullAdder_2361_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2895_io_a = FullAdder_2362_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2895_io_b = FullAdder_2363_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2895_io_ci = FullAdder_2364_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2896_io_a = FullAdder_2365_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2896_io_b = FullAdder_2366_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2896_io_ci = FullAdder_2367_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2897_io_a = FullAdder_2368_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2897_io_b = FullAdder_2369_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2897_io_ci = FullAdder_2370_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2898_io_a = FullAdder_1587_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2898_io_b = FullAdder_2365_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2898_io_ci = FullAdder_2366_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2899_io_a = FullAdder_2367_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2899_io_b = FullAdder_2368_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2899_io_ci = FullAdder_2369_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2900_io_a = FullAdder_2370_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2900_io_b = FullAdder_2371_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2900_io_ci = FullAdder_2372_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2901_io_a = FullAdder_2373_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2901_io_b = FullAdder_2374_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2901_io_ci = FullAdder_2375_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2902_io_a = FullAdder_2376_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2902_io_b = FullAdder_2377_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2902_io_ci = FullAdder_2378_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2903_io_a = FullAdder_1597_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2903_io_b = FullAdder_1598_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2903_io_ci = FullAdder_2372_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2904_io_a = FullAdder_2373_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2904_io_b = FullAdder_2374_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2904_io_ci = FullAdder_2375_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2905_io_a = FullAdder_2376_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2905_io_b = FullAdder_2377_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2905_io_ci = FullAdder_2378_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2906_io_a = FullAdder_2379_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2906_io_b = FullAdder_2380_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2906_io_ci = FullAdder_2381_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2907_io_a = FullAdder_2382_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2907_io_b = FullAdder_2383_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2907_io_ci = FullAdder_2384_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2908_io_a = FullAdder_2379_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2908_io_b = FullAdder_2380_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2908_io_ci = FullAdder_2381_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2909_io_a = FullAdder_2382_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2909_io_b = FullAdder_2383_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2909_io_ci = FullAdder_2384_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2910_io_a = FullAdder_2385_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2910_io_b = HalfAdder_77_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2910_io_ci = FullAdder_2386_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2911_io_a = FullAdder_2387_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2911_io_b = FullAdder_2388_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2911_io_ci = FullAdder_2389_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2912_io_a = FullAdder_2390_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2912_io_b = FullAdder_2391_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2912_io_ci = FullAdder_2392_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2913_io_a = FullAdder_2386_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2913_io_b = FullAdder_2387_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2913_io_ci = FullAdder_2388_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2914_io_a = FullAdder_2389_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2914_io_b = FullAdder_2390_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2914_io_ci = FullAdder_2391_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2915_io_a = FullAdder_2392_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2915_io_b = FullAdder_2393_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2915_io_ci = FullAdder_2394_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2916_io_a = FullAdder_2395_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2916_io_b = FullAdder_2396_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2916_io_ci = FullAdder_2397_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2917_io_a = FullAdder_2398_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2917_io_b = FullAdder_2399_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2917_io_ci = FullAdder_2400_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2918_io_a = FullAdder_2394_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2918_io_b = FullAdder_2395_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2918_io_ci = FullAdder_2396_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2919_io_a = FullAdder_2397_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2919_io_b = FullAdder_2398_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2919_io_ci = FullAdder_2399_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2920_io_a = FullAdder_2400_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2920_io_b = FullAdder_2401_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2920_io_ci = FullAdder_2402_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2921_io_a = FullAdder_2403_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2921_io_b = FullAdder_2404_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2921_io_ci = FullAdder_2405_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2922_io_a = FullAdder_2406_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2922_io_b = FullAdder_2407_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2922_io_ci = FullAdder_2408_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2923_io_a = FullAdder_2402_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2923_io_b = FullAdder_2403_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2923_io_ci = FullAdder_2404_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2924_io_a = FullAdder_2405_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2924_io_b = FullAdder_2406_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2924_io_ci = FullAdder_2407_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2925_io_a = FullAdder_2408_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2925_io_b = FullAdder_2409_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2925_io_ci = FullAdder_2410_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2926_io_a = FullAdder_2411_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2926_io_b = FullAdder_2412_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2926_io_ci = FullAdder_2413_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2927_io_a = FullAdder_2414_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2927_io_b = FullAdder_2415_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2927_io_ci = FullAdder_2416_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2928_io_a = HalfAdder_47_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2928_io_b = FullAdder_2410_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2928_io_ci = FullAdder_2411_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2929_io_a = FullAdder_2412_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2929_io_b = FullAdder_2413_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2929_io_ci = FullAdder_2414_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2930_io_a = FullAdder_2415_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2930_io_b = FullAdder_2416_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2930_io_ci = FullAdder_2417_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2931_io_a = FullAdder_2418_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2931_io_b = FullAdder_2419_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2931_io_ci = FullAdder_2420_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2932_io_a = FullAdder_2421_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2932_io_b = FullAdder_2422_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2932_io_ci = FullAdder_2423_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_102_io_a = FullAdder_2424_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_102_io_b = FullAdder_2425_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2933_io_a = FullAdder_1669_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2933_io_b = HalfAdder_48_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2933_io_ci = FullAdder_2418_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2934_io_a = FullAdder_2419_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2934_io_b = FullAdder_2420_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2934_io_ci = FullAdder_2421_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2935_io_a = FullAdder_2422_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2935_io_b = FullAdder_2423_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2935_io_ci = FullAdder_2424_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2936_io_a = FullAdder_2425_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2936_io_b = FullAdder_2426_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2936_io_ci = FullAdder_2427_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2937_io_a = FullAdder_2428_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2937_io_b = FullAdder_2429_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2937_io_ci = FullAdder_2430_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2938_io_a = FullAdder_2431_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2938_io_b = FullAdder_2432_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2938_io_ci = FullAdder_2433_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2939_io_a = FullAdder_1681_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2939_io_b = FullAdder_2426_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2939_io_ci = FullAdder_2427_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2940_io_a = FullAdder_2428_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2940_io_b = FullAdder_2429_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2940_io_ci = FullAdder_2430_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2941_io_a = FullAdder_2431_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2941_io_b = FullAdder_2432_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2941_io_ci = FullAdder_2433_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2942_io_a = FullAdder_2434_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2942_io_b = FullAdder_2435_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2942_io_ci = FullAdder_2436_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2943_io_a = FullAdder_2437_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2943_io_b = FullAdder_2438_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2943_io_ci = FullAdder_2439_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2944_io_a = FullAdder_2440_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2944_io_b = FullAdder_2441_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2944_io_ci = FullAdder_2442_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2945_io_a = FullAdder_2434_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2945_io_b = FullAdder_2435_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2945_io_ci = FullAdder_2436_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2946_io_a = FullAdder_2437_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2946_io_b = FullAdder_2438_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2946_io_ci = FullAdder_2439_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2947_io_a = FullAdder_2440_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2947_io_b = FullAdder_2441_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2947_io_ci = FullAdder_2442_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2948_io_a = FullAdder_2443_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2948_io_b = FullAdder_2444_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2948_io_ci = FullAdder_2445_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2949_io_a = FullAdder_2446_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2949_io_b = FullAdder_2447_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2949_io_ci = FullAdder_2448_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2950_io_a = FullAdder_2449_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2950_io_b = FullAdder_2450_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2950_io_ci = FullAdder_2451_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2951_io_a = FullAdder_2443_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2951_io_b = FullAdder_2444_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2951_io_ci = FullAdder_2445_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2952_io_a = FullAdder_2446_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2952_io_b = FullAdder_2447_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2952_io_ci = FullAdder_2448_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2953_io_a = FullAdder_2449_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2953_io_b = FullAdder_2450_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2953_io_ci = FullAdder_2451_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2954_io_a = FullAdder_2452_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2954_io_b = FullAdder_2453_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2954_io_ci = FullAdder_2454_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2955_io_a = FullAdder_2455_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2955_io_b = FullAdder_2456_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2955_io_ci = FullAdder_2457_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2956_io_a = FullAdder_2458_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2956_io_b = FullAdder_2459_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2956_io_ci = FullAdder_2460_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2957_io_a = FullAdder_2452_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2957_io_b = FullAdder_2453_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2957_io_ci = FullAdder_2454_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2958_io_a = FullAdder_2455_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2958_io_b = FullAdder_2456_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2958_io_ci = FullAdder_2457_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2959_io_a = FullAdder_2458_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2959_io_b = FullAdder_2459_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2959_io_ci = FullAdder_2460_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2960_io_a = FullAdder_2461_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2960_io_b = FullAdder_2462_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2960_io_ci = FullAdder_2463_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2961_io_a = FullAdder_2464_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2961_io_b = FullAdder_2465_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2961_io_ci = FullAdder_2466_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2962_io_a = FullAdder_2467_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2962_io_b = FullAdder_2468_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2962_io_ci = FullAdder_2469_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2963_io_a = FullAdder_1734_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2963_io_b = FullAdder_2461_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2963_io_ci = FullAdder_2462_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2964_io_a = FullAdder_2463_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2964_io_b = FullAdder_2464_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2964_io_ci = FullAdder_2465_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2965_io_a = FullAdder_2466_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2965_io_b = FullAdder_2467_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2965_io_ci = FullAdder_2468_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2966_io_a = FullAdder_2469_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2966_io_b = FullAdder_2470_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2966_io_ci = FullAdder_2471_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2967_io_a = FullAdder_2472_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2967_io_b = FullAdder_2473_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2967_io_ci = FullAdder_2474_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2968_io_a = FullAdder_2475_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2968_io_b = FullAdder_2476_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2968_io_ci = FullAdder_2477_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2969_io_a = FullAdder_1748_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2969_io_b = FullAdder_2470_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2969_io_ci = FullAdder_2471_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2970_io_a = FullAdder_2472_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2970_io_b = FullAdder_2473_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2970_io_ci = FullAdder_2474_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2971_io_a = FullAdder_2475_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2971_io_b = FullAdder_2476_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2971_io_ci = FullAdder_2477_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2972_io_a = FullAdder_2478_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2972_io_b = FullAdder_2479_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2972_io_ci = FullAdder_2480_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2973_io_a = FullAdder_2481_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2973_io_b = FullAdder_2482_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2973_io_ci = FullAdder_2483_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2974_io_a = FullAdder_2484_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2974_io_b = FullAdder_2485_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2974_io_ci = FullAdder_2486_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2975_io_a = FullAdder_1762_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2975_io_b = FullAdder_2479_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2975_io_ci = FullAdder_2480_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2976_io_a = FullAdder_2481_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2976_io_b = FullAdder_2482_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2976_io_ci = FullAdder_2483_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2977_io_a = FullAdder_2484_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2977_io_b = FullAdder_2485_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2977_io_ci = FullAdder_2486_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2978_io_a = FullAdder_2487_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2978_io_b = FullAdder_2488_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2978_io_ci = FullAdder_2489_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2979_io_a = FullAdder_2490_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2979_io_b = FullAdder_2491_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2979_io_ci = FullAdder_2492_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2980_io_a = FullAdder_2493_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2980_io_b = FullAdder_2494_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2980_io_ci = FullAdder_2495_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2981_io_a = FullAdder_1776_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2981_io_b = FullAdder_2488_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2981_io_ci = FullAdder_2489_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2982_io_a = FullAdder_2490_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2982_io_b = FullAdder_2491_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2982_io_ci = FullAdder_2492_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2983_io_a = FullAdder_2493_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2983_io_b = FullAdder_2494_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2983_io_ci = FullAdder_2495_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2984_io_a = FullAdder_2496_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2984_io_b = FullAdder_2497_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2984_io_ci = FullAdder_2498_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2985_io_a = FullAdder_2499_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2985_io_b = FullAdder_2500_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2985_io_ci = FullAdder_2501_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2986_io_a = FullAdder_2502_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2986_io_b = FullAdder_2503_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2986_io_ci = FullAdder_2504_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_103_io_a = FullAdder_2505_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_103_io_b = HalfAdder_78_io_co; // @[wallace.scala 60:18]
  assign FullAdder_2987_io_a = FullAdder_2497_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2987_io_b = FullAdder_2498_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2987_io_ci = FullAdder_2499_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2988_io_a = FullAdder_2500_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2988_io_b = FullAdder_2501_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2988_io_ci = FullAdder_2502_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2989_io_a = FullAdder_2503_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2989_io_b = FullAdder_2504_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2989_io_ci = FullAdder_2505_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2990_io_a = HalfAdder_78_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2990_io_b = FullAdder_2506_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2990_io_ci = FullAdder_2507_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2991_io_a = FullAdder_2508_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2991_io_b = FullAdder_2509_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2991_io_ci = FullAdder_2510_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2992_io_a = FullAdder_2511_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2992_io_b = FullAdder_2512_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2992_io_ci = FullAdder_2513_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2993_io_a = HalfAdder_49_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2993_io_b = FullAdder_2506_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2993_io_ci = FullAdder_2507_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2994_io_a = FullAdder_2508_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2994_io_b = FullAdder_2509_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2994_io_ci = FullAdder_2510_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2995_io_a = FullAdder_2511_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2995_io_b = FullAdder_2512_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2995_io_ci = FullAdder_2513_io_s; // @[wallace.scala 71:19]
  assign FullAdder_2996_io_a = FullAdder_2514_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2996_io_b = FullAdder_2515_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2996_io_ci = FullAdder_2516_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2997_io_a = FullAdder_2517_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2997_io_b = FullAdder_2518_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2997_io_ci = FullAdder_2519_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2998_io_a = FullAdder_2520_io_co; // @[wallace.scala 69:18]
  assign FullAdder_2998_io_b = FullAdder_2521_io_co; // @[wallace.scala 70:18]
  assign FullAdder_2998_io_ci = FullAdder_2522_io_co; // @[wallace.scala 71:19]
  assign FullAdder_2999_io_a = FullAdder_2515_io_s; // @[wallace.scala 69:18]
  assign FullAdder_2999_io_b = FullAdder_2516_io_s; // @[wallace.scala 70:18]
  assign FullAdder_2999_io_ci = FullAdder_2517_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3000_io_a = FullAdder_2518_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3000_io_b = FullAdder_2519_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3000_io_ci = FullAdder_2520_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3001_io_a = FullAdder_2521_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3001_io_b = FullAdder_2522_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3001_io_ci = FullAdder_2523_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3002_io_a = FullAdder_2524_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3002_io_b = FullAdder_2525_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3002_io_ci = FullAdder_2526_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3003_io_a = FullAdder_2527_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3003_io_b = FullAdder_2528_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3003_io_ci = FullAdder_2529_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3004_io_a = FullAdder_2530_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3004_io_b = FullAdder_2531_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3004_io_ci = FullAdder_2532_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3005_io_a = FullAdder_1829_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3005_io_b = FullAdder_2524_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3005_io_ci = FullAdder_2525_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3006_io_a = FullAdder_2526_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3006_io_b = FullAdder_2527_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3006_io_ci = FullAdder_2528_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3007_io_a = FullAdder_2529_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3007_io_b = FullAdder_2530_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3007_io_ci = FullAdder_2531_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3008_io_a = FullAdder_2532_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3008_io_b = FullAdder_2533_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3008_io_ci = FullAdder_2534_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3009_io_a = FullAdder_2535_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3009_io_b = FullAdder_2536_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3009_io_ci = FullAdder_2537_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3010_io_a = FullAdder_2538_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3010_io_b = FullAdder_2539_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3010_io_ci = FullAdder_2540_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3011_io_a = FullAdder_2533_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3011_io_b = FullAdder_2534_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3011_io_ci = FullAdder_2535_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3012_io_a = FullAdder_2536_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3012_io_b = FullAdder_2537_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3012_io_ci = FullAdder_2538_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3013_io_a = FullAdder_2539_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3013_io_b = FullAdder_2540_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3013_io_ci = FullAdder_2541_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3014_io_a = FullAdder_2542_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3014_io_b = FullAdder_2543_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3014_io_ci = FullAdder_2544_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3015_io_a = FullAdder_2545_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3015_io_b = FullAdder_2546_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3015_io_ci = FullAdder_2547_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3016_io_a = FullAdder_2548_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3016_io_b = FullAdder_2549_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3016_io_ci = HalfAdder_79_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3017_io_a = FullAdder_2542_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3017_io_b = FullAdder_2543_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3017_io_ci = FullAdder_2544_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3018_io_a = FullAdder_2545_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3018_io_b = FullAdder_2546_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3018_io_ci = FullAdder_2547_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3019_io_a = FullAdder_2548_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3019_io_b = FullAdder_2549_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3019_io_ci = HalfAdder_79_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3020_io_a = FullAdder_2550_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3020_io_b = FullAdder_2551_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3020_io_ci = FullAdder_2552_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3021_io_a = FullAdder_2553_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3021_io_b = FullAdder_2554_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3021_io_ci = FullAdder_2555_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3022_io_a = FullAdder_1867_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3022_io_b = FullAdder_2550_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3022_io_ci = FullAdder_2551_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3023_io_a = FullAdder_2552_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3023_io_b = FullAdder_2553_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3023_io_ci = FullAdder_2554_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3024_io_a = FullAdder_2555_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3024_io_b = FullAdder_2556_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3024_io_ci = FullAdder_2557_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3025_io_a = FullAdder_2558_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3025_io_b = FullAdder_2559_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3025_io_ci = FullAdder_2560_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3026_io_a = FullAdder_2561_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3026_io_b = FullAdder_2562_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3026_io_ci = FullAdder_2563_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_104_io_a = FullAdder_2564_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_104_io_b = FullAdder_2565_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3027_io_a = FullAdder_1879_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3027_io_b = FullAdder_2558_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3027_io_ci = FullAdder_2559_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3028_io_a = FullAdder_2560_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3028_io_b = FullAdder_2561_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3028_io_ci = FullAdder_2562_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3029_io_a = FullAdder_2563_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3029_io_b = FullAdder_2564_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3029_io_ci = FullAdder_2565_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3030_io_a = FullAdder_2566_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3030_io_b = FullAdder_2567_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3030_io_ci = FullAdder_2568_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3031_io_a = FullAdder_2569_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3031_io_b = FullAdder_2570_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3031_io_ci = FullAdder_2571_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_105_io_a = FullAdder_2572_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_105_io_b = FullAdder_2573_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3032_io_a = FullAdder_1890_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3032_io_b = FullAdder_1891_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3032_io_ci = FullAdder_2566_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3033_io_a = FullAdder_2567_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3033_io_b = FullAdder_2568_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3033_io_ci = FullAdder_2569_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3034_io_a = FullAdder_2570_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3034_io_b = FullAdder_2571_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3034_io_ci = FullAdder_2572_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3035_io_a = FullAdder_2573_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3035_io_b = FullAdder_2574_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3035_io_ci = FullAdder_2575_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3036_io_a = FullAdder_2576_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3036_io_b = FullAdder_2577_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3036_io_ci = FullAdder_2578_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3037_io_a = FullAdder_2579_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3037_io_b = FullAdder_2580_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3037_io_ci = FullAdder_2581_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3038_io_a = FullAdder_1903_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3038_io_b = FullAdder_2574_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3038_io_ci = FullAdder_2575_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3039_io_a = FullAdder_2576_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3039_io_b = FullAdder_2577_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3039_io_ci = FullAdder_2578_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3040_io_a = FullAdder_2579_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3040_io_b = FullAdder_2580_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3040_io_ci = FullAdder_2581_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3041_io_a = FullAdder_2582_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3041_io_b = FullAdder_2583_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3041_io_ci = FullAdder_2584_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3042_io_a = FullAdder_2585_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3042_io_b = FullAdder_2586_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3042_io_ci = FullAdder_2587_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3043_io_a = FullAdder_1913_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3043_io_b = FullAdder_1914_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3043_io_ci = FullAdder_2582_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3044_io_a = FullAdder_2583_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3044_io_b = FullAdder_2584_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3044_io_ci = FullAdder_2585_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3045_io_a = FullAdder_2586_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3045_io_b = FullAdder_2587_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3045_io_ci = FullAdder_2588_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3046_io_a = FullAdder_2589_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3046_io_b = FullAdder_2590_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3046_io_ci = FullAdder_2591_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3047_io_a = FullAdder_2592_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3047_io_b = FullAdder_2593_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3047_io_ci = FullAdder_2594_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3048_io_a = HalfAdder_50_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3048_io_b = FullAdder_2589_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3048_io_ci = FullAdder_2590_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3049_io_a = FullAdder_2591_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3049_io_b = FullAdder_2592_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3049_io_ci = FullAdder_2593_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3050_io_a = FullAdder_2594_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3050_io_b = FullAdder_2595_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3050_io_ci = FullAdder_2596_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3051_io_a = FullAdder_2597_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3051_io_b = FullAdder_2598_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3051_io_ci = FullAdder_2599_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3052_io_a = FullAdder_2600_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3052_io_b = FullAdder_2601_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3052_io_ci = FullAdder_2602_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3053_io_a = FullAdder_2597_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3053_io_b = FullAdder_2598_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3053_io_ci = FullAdder_2599_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3054_io_a = FullAdder_2600_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3054_io_b = FullAdder_2601_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3054_io_ci = FullAdder_2602_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3055_io_a = FullAdder_2603_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3055_io_b = HalfAdder_80_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3055_io_ci = FullAdder_2604_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3056_io_a = FullAdder_2605_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3056_io_b = FullAdder_2606_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3056_io_ci = FullAdder_2607_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3057_io_a = FullAdder_2608_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3057_io_b = FullAdder_2609_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3057_io_ci = FullAdder_2610_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3058_io_a = FullAdder_1947_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3058_io_b = FullAdder_2604_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3058_io_ci = FullAdder_2605_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3059_io_a = FullAdder_2606_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3059_io_b = FullAdder_2607_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3059_io_ci = FullAdder_2608_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3060_io_a = FullAdder_2609_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3060_io_b = FullAdder_2610_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3060_io_ci = FullAdder_2611_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3061_io_a = FullAdder_2612_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3061_io_b = FullAdder_2613_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3061_io_ci = FullAdder_2614_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3062_io_a = FullAdder_2615_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3062_io_b = FullAdder_2616_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3062_io_ci = FullAdder_2617_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3063_io_a = FullAdder_1957_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3063_io_b = FullAdder_1958_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3063_io_ci = FullAdder_2611_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3064_io_a = FullAdder_2612_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3064_io_b = FullAdder_2613_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3064_io_ci = FullAdder_2614_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3065_io_a = FullAdder_2615_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3065_io_b = FullAdder_2616_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3065_io_ci = FullAdder_2617_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3066_io_a = FullAdder_2618_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3066_io_b = FullAdder_2619_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3066_io_ci = FullAdder_2620_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3067_io_a = FullAdder_2621_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3067_io_b = FullAdder_2622_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3067_io_ci = FullAdder_2623_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3068_io_a = HalfAdder_51_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3068_io_b = FullAdder_2618_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3068_io_ci = FullAdder_2619_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3069_io_a = FullAdder_2620_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3069_io_b = FullAdder_2621_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3069_io_ci = FullAdder_2622_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3070_io_a = FullAdder_2623_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3070_io_b = FullAdder_2624_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3070_io_ci = FullAdder_2625_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3071_io_a = FullAdder_2626_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3071_io_b = FullAdder_2627_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3071_io_ci = FullAdder_2628_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3072_io_a = FullAdder_2629_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3072_io_b = FullAdder_2630_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3072_io_ci = FullAdder_2631_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3073_io_a = FullAdder_2625_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3073_io_b = FullAdder_2626_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3073_io_ci = FullAdder_2627_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3074_io_a = FullAdder_2628_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3074_io_b = FullAdder_2629_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3074_io_ci = FullAdder_2630_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3075_io_a = FullAdder_2631_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3075_io_b = FullAdder_2632_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3075_io_ci = FullAdder_2633_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3076_io_a = FullAdder_2634_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3076_io_b = FullAdder_2635_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3076_io_ci = FullAdder_2636_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_106_io_a = FullAdder_2637_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_106_io_b = FullAdder_2638_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3077_io_a = FullAdder_2632_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3077_io_b = FullAdder_2633_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3077_io_ci = FullAdder_2634_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3078_io_a = FullAdder_2635_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3078_io_b = FullAdder_2636_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3078_io_ci = FullAdder_2637_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3079_io_a = FullAdder_2638_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3079_io_b = FullAdder_2639_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3079_io_ci = FullAdder_2640_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3080_io_a = FullAdder_2641_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3080_io_b = FullAdder_2642_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3080_io_ci = FullAdder_2643_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3081_io_a = FullAdder_2639_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3081_io_b = FullAdder_2640_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3081_io_ci = FullAdder_2641_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3082_io_a = FullAdder_2642_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3082_io_b = FullAdder_2643_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3082_io_ci = FullAdder_2644_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3083_io_a = HalfAdder_81_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3083_io_b = FullAdder_2645_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3083_io_ci = FullAdder_2646_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3084_io_a = FullAdder_2647_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3084_io_b = FullAdder_2648_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3084_io_ci = FullAdder_2649_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3085_io_a = FullAdder_2645_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3085_io_b = FullAdder_2646_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3085_io_ci = FullAdder_2647_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3086_io_a = FullAdder_2648_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3086_io_b = FullAdder_2649_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3086_io_ci = FullAdder_2650_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3087_io_a = FullAdder_2651_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3087_io_b = FullAdder_2652_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3087_io_ci = FullAdder_2653_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3088_io_a = FullAdder_2654_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3088_io_b = FullAdder_2655_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3088_io_ci = FullAdder_2656_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3089_io_a = FullAdder_2016_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3089_io_b = HalfAdder_52_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3089_io_ci = FullAdder_2652_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3090_io_a = FullAdder_2653_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3090_io_b = FullAdder_2654_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3090_io_ci = FullAdder_2655_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3091_io_a = FullAdder_2656_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3091_io_b = FullAdder_2657_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3091_io_ci = FullAdder_2658_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3092_io_a = FullAdder_2659_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3092_io_b = FullAdder_2660_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3092_io_ci = FullAdder_2661_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3093_io_a = FullAdder_2025_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3093_io_b = FullAdder_2658_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3093_io_ci = FullAdder_2659_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3094_io_a = FullAdder_2660_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3094_io_b = FullAdder_2661_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3094_io_ci = FullAdder_2662_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3095_io_a = FullAdder_2663_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3095_io_b = FullAdder_2664_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3095_io_ci = FullAdder_2665_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3096_io_a = FullAdder_2666_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3096_io_b = FullAdder_2667_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3096_io_ci = FullAdder_2668_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3097_io_a = FullAdder_2664_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3097_io_b = FullAdder_2665_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3097_io_ci = FullAdder_2666_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3098_io_a = FullAdder_2667_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3098_io_b = FullAdder_2668_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3098_io_ci = FullAdder_2669_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3099_io_a = FullAdder_2670_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3099_io_b = FullAdder_2671_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3099_io_ci = FullAdder_2672_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3100_io_a = FullAdder_2673_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3100_io_b = FullAdder_2674_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3100_io_ci = FullAdder_2675_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3101_io_a = FullAdder_2043_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3101_io_b = FullAdder_2670_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3101_io_ci = FullAdder_2671_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3102_io_a = FullAdder_2672_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3102_io_b = FullAdder_2673_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3102_io_ci = FullAdder_2674_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3103_io_a = FullAdder_2675_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3103_io_b = FullAdder_2676_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3103_io_ci = FullAdder_2677_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3104_io_a = FullAdder_2678_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3104_io_b = FullAdder_2679_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3104_io_ci = FullAdder_2680_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3105_io_a = FullAdder_2676_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3105_io_b = FullAdder_2677_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3105_io_ci = FullAdder_2678_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3106_io_a = FullAdder_2679_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3106_io_b = FullAdder_2680_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3106_io_ci = FullAdder_2681_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3107_io_a = FullAdder_2682_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3107_io_b = FullAdder_2683_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3107_io_ci = FullAdder_2684_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3108_io_a = FullAdder_2058_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3108_io_b = FullAdder_2059_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3108_io_ci = FullAdder_2682_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3109_io_a = FullAdder_2683_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3109_io_b = FullAdder_2684_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3109_io_ci = FullAdder_2685_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3110_io_a = FullAdder_2686_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3110_io_b = FullAdder_2687_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3110_io_ci = FullAdder_2688_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3111_io_a = FullAdder_2689_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3111_io_b = FullAdder_2690_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3111_io_ci = FullAdder_2691_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3112_io_a = FullAdder_2687_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3112_io_b = FullAdder_2688_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3112_io_ci = FullAdder_2689_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3113_io_a = FullAdder_2690_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3113_io_b = FullAdder_2691_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3113_io_ci = HalfAdder_82_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3114_io_a = FullAdder_2692_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3114_io_b = FullAdder_2693_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3114_io_ci = FullAdder_2694_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3115_io_a = FullAdder_2695_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3115_io_b = FullAdder_2696_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3115_io_ci = HalfAdder_83_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3116_io_a = FullAdder_2692_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3116_io_b = FullAdder_2693_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3116_io_ci = FullAdder_2694_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3117_io_a = FullAdder_2695_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3117_io_b = FullAdder_2696_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3117_io_ci = HalfAdder_83_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3118_io_a = FullAdder_2697_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3118_io_b = FullAdder_2698_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3118_io_ci = FullAdder_2699_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_107_io_a = FullAdder_2700_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_107_io_b = FullAdder_2701_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3119_io_a = FullAdder_2697_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3119_io_b = FullAdder_2698_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3119_io_ci = FullAdder_2699_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3120_io_a = FullAdder_2700_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3120_io_b = FullAdder_2701_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3120_io_ci = FullAdder_2702_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3121_io_a = FullAdder_2703_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3121_io_b = FullAdder_2704_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3121_io_ci = FullAdder_2705_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3122_io_a = FullAdder_2089_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3122_io_b = HalfAdder_54_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3122_io_ci = FullAdder_2702_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3123_io_a = FullAdder_2703_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3123_io_b = FullAdder_2704_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3123_io_ci = FullAdder_2705_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3124_io_a = FullAdder_2706_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3124_io_b = FullAdder_2707_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3124_io_ci = FullAdder_2708_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3125_io_a = FullAdder_2709_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3125_io_b = FullAdder_2710_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3125_io_ci = FullAdder_2711_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3126_io_a = FullAdder_2707_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3126_io_b = FullAdder_2708_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3126_io_ci = FullAdder_2709_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3127_io_a = FullAdder_2710_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3127_io_b = FullAdder_2711_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3127_io_ci = FullAdder_2712_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3128_io_a = FullAdder_2713_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3128_io_b = FullAdder_2714_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3128_io_ci = FullAdder_2715_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3129_io_a = FullAdder_2712_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3129_io_b = FullAdder_2713_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3129_io_ci = FullAdder_2714_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3130_io_a = FullAdder_2715_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3130_io_b = FullAdder_2716_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3130_io_ci = FullAdder_2717_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3131_io_a = FullAdder_2718_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3131_io_b = FullAdder_2719_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3131_io_ci = FullAdder_2720_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3132_io_a = FullAdder_2109_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3132_io_b = FullAdder_2110_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3132_io_ci = FullAdder_2717_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3133_io_a = FullAdder_2718_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3133_io_b = FullAdder_2719_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3133_io_ci = FullAdder_2720_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3134_io_a = FullAdder_2721_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3134_io_b = FullAdder_2722_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3134_io_ci = FullAdder_2723_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3135_io_a = FullAdder_2721_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3135_io_b = FullAdder_2722_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3135_io_ci = FullAdder_2723_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3136_io_a = FullAdder_2724_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3136_io_b = HalfAdder_84_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3136_io_ci = FullAdder_2725_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3137_io_a = FullAdder_2726_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3137_io_b = FullAdder_2727_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3137_io_ci = FullAdder_2728_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3138_io_a = FullAdder_2122_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3138_io_b = FullAdder_2725_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3138_io_ci = FullAdder_2726_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3139_io_a = FullAdder_2727_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3139_io_b = FullAdder_2728_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3139_io_ci = FullAdder_2729_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3140_io_a = FullAdder_2730_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3140_io_b = FullAdder_2731_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3140_io_ci = FullAdder_2732_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3141_io_a = FullAdder_2128_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3141_io_b = FullAdder_2729_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3141_io_ci = FullAdder_2730_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3142_io_a = FullAdder_2731_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3142_io_b = FullAdder_2732_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3142_io_ci = FullAdder_2733_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3143_io_a = FullAdder_2734_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3143_io_b = FullAdder_2735_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3143_io_ci = FullAdder_2736_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3144_io_a = HalfAdder_56_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3144_io_b = FullAdder_2733_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3144_io_ci = FullAdder_2734_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3145_io_a = FullAdder_2735_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3145_io_b = FullAdder_2736_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3145_io_ci = FullAdder_2737_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3146_io_a = FullAdder_2738_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3146_io_b = FullAdder_2739_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3146_io_ci = FullAdder_2740_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3147_io_a = FullAdder_2737_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3147_io_b = FullAdder_2738_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3147_io_ci = FullAdder_2739_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3148_io_a = FullAdder_2740_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3148_io_b = FullAdder_2741_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3148_io_ci = FullAdder_2742_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3149_io_a = FullAdder_2143_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3149_io_b = FullAdder_2144_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3149_io_ci = FullAdder_2741_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3150_io_a = FullAdder_2742_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3150_io_b = FullAdder_2743_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3150_io_ci = FullAdder_2744_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3151_io_a = FullAdder_2745_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3151_io_b = FullAdder_2746_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3151_io_ci = FullAdder_2747_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3152_io_a = FullAdder_2744_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3152_io_b = FullAdder_2745_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3152_io_ci = FullAdder_2746_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3153_io_a = FullAdder_2747_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3153_io_b = FullAdder_2748_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3153_io_ci = FullAdder_2749_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3154_io_a = FullAdder_2748_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3154_io_b = FullAdder_2749_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3154_io_ci = FullAdder_2750_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3155_io_a = HalfAdder_85_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3155_io_b = FullAdder_2751_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3155_io_ci = FullAdder_2752_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3156_io_a = FullAdder_2159_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3156_io_b = FullAdder_2751_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3156_io_ci = FullAdder_2752_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3157_io_a = FullAdder_2753_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3157_io_b = FullAdder_2754_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3157_io_ci = FullAdder_2755_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3158_io_a = HalfAdder_57_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3158_io_b = FullAdder_2754_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3158_io_ci = FullAdder_2755_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3159_io_a = FullAdder_2756_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3159_io_b = FullAdder_2757_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3159_io_ci = FullAdder_2758_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3160_io_a = FullAdder_2757_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3160_io_b = FullAdder_2758_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3160_io_ci = FullAdder_2759_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3161_io_a = FullAdder_2760_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3161_io_b = FullAdder_2761_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3161_io_ci = FullAdder_2762_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3162_io_a = FullAdder_2760_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3162_io_b = FullAdder_2761_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3162_io_ci = FullAdder_2762_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3163_io_a = FullAdder_2763_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3163_io_b = FullAdder_2764_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3163_io_ci = FullAdder_2765_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3164_io_a = FullAdder_2763_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3164_io_b = FullAdder_2764_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3164_io_ci = FullAdder_2765_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3165_io_a = FullAdder_2178_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3165_io_b = HalfAdder_58_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3165_io_ci = FullAdder_2766_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3166_io_a = FullAdder_2767_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3166_io_b = FullAdder_2768_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3166_io_ci = FullAdder_2769_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3167_io_a = FullAdder_2768_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3167_io_b = FullAdder_2769_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3167_io_ci = HalfAdder_86_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_108_io_a = FullAdder_2770_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_108_io_b = FullAdder_2771_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3168_io_a = FullAdder_2184_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3168_io_b = FullAdder_2770_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3168_io_ci = FullAdder_2771_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3169_io_a = FullAdder_2187_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3169_io_b = FullAdder_2772_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3169_io_ci = FullAdder_2773_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_109_io_a = FullAdder_2774_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_109_io_b = FullAdder_2775_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3170_io_a = FullAdder_2774_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3170_io_b = FullAdder_2775_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3170_io_ci = FullAdder_2776_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3171_io_a = FullAdder_2191_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3171_io_b = FullAdder_2192_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3171_io_ci = FullAdder_2776_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3172_io_a = HalfAdder_61_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3172_io_b = FullAdder_2777_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3172_io_ci = FullAdder_2778_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_110_io_a = FullAdder_2195_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_110_io_b = HalfAdder_87_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_111_io_a = HalfAdder_88_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_111_io_b = FullAdder_2779_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3173_io_a = FullAdder_2779_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3173_io_b = HalfAdder_89_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3173_io_ci = FullAdder_2780_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3174_io_a = HalfAdder_62_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3174_io_b = FullAdder_2780_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3174_io_ci = FullAdder_2781_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3175_io_a = HalfAdder_63_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3175_io_b = FullAdder_2781_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3175_io_ci = FullAdder_2782_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_112_io_a = FullAdder_2782_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_112_io_b = FullAdder_2783_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_113_io_a = FullAdder_2783_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_113_io_b = HalfAdder_90_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_114_io_a = FullAdder_2201_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_114_io_b = HalfAdder_90_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_115_io_a = HalfAdder_92_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_115_io_b = HalfAdder_93_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3176_io_a = HalfAdder_68_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3176_io_b = HalfAdder_69_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3176_io_ci = HalfAdder_94_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_116_io_a = FullAdder_2202_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_116_io_b = HalfAdder_94_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_117_io_a = HalfAdder_95_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_117_io_b = FullAdder_2784_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3177_io_a = HalfAdder_71_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3177_io_b = FullAdder_2784_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3177_io_ci = HalfAdder_96_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_118_io_a = FullAdder_2204_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_118_io_b = HalfAdder_96_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_119_io_a = FullAdder_2785_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_119_io_b = FullAdder_2786_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3178_io_a = FullAdder_2207_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3178_io_b = FullAdder_2786_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3178_io_ci = FullAdder_2787_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3179_io_a = FullAdder_2208_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3179_io_b = FullAdder_2209_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3179_io_ci = FullAdder_2787_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3180_io_a = FullAdder_2211_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3180_io_b = FullAdder_2788_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3180_io_ci = FullAdder_2789_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3181_io_a = FullAdder_2213_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3181_io_b = FullAdder_2789_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3181_io_ci = FullAdder_2790_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3182_io_a = FullAdder_2215_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3182_io_b = FullAdder_2790_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3182_io_ci = FullAdder_2791_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3183_io_a = HalfAdder_72_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3183_io_b = FullAdder_2791_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3183_io_ci = FullAdder_2792_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3184_io_a = FullAdder_2218_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3184_io_b = FullAdder_2219_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3184_io_ci = FullAdder_2793_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3185_io_a = HalfAdder_73_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3185_io_b = FullAdder_2794_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3185_io_ci = FullAdder_2795_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3186_io_a = FullAdder_2796_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3186_io_b = FullAdder_2797_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3186_io_ci = FullAdder_2798_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3187_io_a = FullAdder_2798_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3187_io_b = FullAdder_2799_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3187_io_ci = FullAdder_2800_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3188_io_a = FullAdder_2230_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3188_io_b = FullAdder_2800_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3188_io_ci = FullAdder_2801_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_120_io_a = FullAdder_2802_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_120_io_b = FullAdder_2803_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3189_io_a = FullAdder_2233_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3189_io_b = FullAdder_2802_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3189_io_ci = FullAdder_2803_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_121_io_a = FullAdder_2804_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_121_io_b = FullAdder_2805_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3190_io_a = FullAdder_2236_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3190_io_b = FullAdder_2804_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3190_io_ci = FullAdder_2805_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3191_io_a = FullAdder_2806_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3191_io_b = FullAdder_2807_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3191_io_ci = FullAdder_2808_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3192_io_a = FullAdder_2806_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3192_io_b = FullAdder_2807_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3192_io_ci = FullAdder_2808_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3193_io_a = FullAdder_2242_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3193_io_b = FullAdder_2809_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3193_io_ci = FullAdder_2810_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3194_io_a = FullAdder_2811_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3194_io_b = FullAdder_2812_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3194_io_ci = FullAdder_2813_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3195_io_a = FullAdder_2811_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3195_io_b = FullAdder_2812_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3195_io_ci = FullAdder_2813_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3196_io_a = FullAdder_2814_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3196_io_b = FullAdder_2815_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3196_io_ci = FullAdder_2816_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3197_io_a = FullAdder_2814_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3197_io_b = FullAdder_2815_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3197_io_ci = FullAdder_2816_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3198_io_a = FullAdder_2817_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3198_io_b = FullAdder_2818_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3198_io_ci = FullAdder_2819_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3199_io_a = FullAdder_2817_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3199_io_b = FullAdder_2818_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3199_io_ci = FullAdder_2819_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3200_io_a = FullAdder_2820_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3200_io_b = FullAdder_2821_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3200_io_ci = HalfAdder_97_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3201_io_a = FullAdder_2820_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3201_io_b = FullAdder_2821_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3201_io_ci = HalfAdder_97_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3202_io_a = FullAdder_2822_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3202_io_b = FullAdder_2823_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3202_io_ci = FullAdder_2824_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3203_io_a = FullAdder_2262_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3203_io_b = FullAdder_2822_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3203_io_ci = FullAdder_2823_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3204_io_a = FullAdder_2824_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3204_io_b = FullAdder_2825_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3204_io_ci = FullAdder_2826_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3205_io_a = FullAdder_2266_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3205_io_b = FullAdder_2825_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3205_io_ci = FullAdder_2826_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3206_io_a = FullAdder_2827_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3206_io_b = FullAdder_2828_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3206_io_ci = FullAdder_2829_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3207_io_a = FullAdder_2270_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3207_io_b = FullAdder_2271_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3207_io_ci = FullAdder_2828_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3208_io_a = FullAdder_2829_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3208_io_b = FullAdder_2830_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3208_io_ci = FullAdder_2831_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3209_io_a = FullAdder_2276_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3209_io_b = FullAdder_2831_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3209_io_ci = FullAdder_2832_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3210_io_a = FullAdder_2833_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3210_io_b = FullAdder_2834_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3210_io_ci = FullAdder_2835_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3211_io_a = FullAdder_2281_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3211_io_b = FullAdder_2834_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3211_io_ci = FullAdder_2835_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3212_io_a = FullAdder_2836_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3212_io_b = FullAdder_2837_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3212_io_ci = FullAdder_2838_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3213_io_a = FullAdder_2837_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3213_io_b = FullAdder_2838_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3213_io_ci = FullAdder_2839_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3214_io_a = HalfAdder_98_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3214_io_b = FullAdder_2840_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3214_io_ci = FullAdder_2841_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_122_io_a = FullAdder_2842_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_122_io_b = HalfAdder_99_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3215_io_a = FullAdder_2840_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3215_io_b = FullAdder_2841_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3215_io_ci = FullAdder_2842_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3216_io_a = HalfAdder_99_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3216_io_b = FullAdder_2843_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3216_io_ci = FullAdder_2844_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_123_io_a = FullAdder_2845_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_123_io_b = HalfAdder_100_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3217_io_a = FullAdder_2843_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3217_io_b = FullAdder_2844_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3217_io_ci = FullAdder_2845_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3218_io_a = HalfAdder_100_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3218_io_b = FullAdder_2846_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3218_io_ci = FullAdder_2847_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_124_io_a = FullAdder_2848_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_124_io_b = FullAdder_2849_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3219_io_a = FullAdder_2302_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3219_io_b = FullAdder_2846_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3219_io_ci = FullAdder_2847_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3220_io_a = FullAdder_2848_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3220_io_b = FullAdder_2849_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3220_io_ci = FullAdder_2850_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3221_io_a = FullAdder_2851_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3221_io_b = FullAdder_2852_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3221_io_ci = FullAdder_2853_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3222_io_a = FullAdder_2850_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3222_io_b = FullAdder_2851_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3222_io_ci = FullAdder_2852_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3223_io_a = FullAdder_2853_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3223_io_b = FullAdder_2854_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3223_io_ci = FullAdder_2855_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3224_io_a = FullAdder_2854_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3224_io_b = FullAdder_2855_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3224_io_ci = FullAdder_2856_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3225_io_a = FullAdder_2857_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3225_io_b = FullAdder_2858_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3225_io_ci = FullAdder_2859_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_125_io_a = FullAdder_2860_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_125_io_b = FullAdder_2861_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3226_io_a = FullAdder_2858_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3226_io_b = FullAdder_2859_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3226_io_ci = FullAdder_2860_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3227_io_a = FullAdder_2861_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3227_io_b = FullAdder_2862_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3227_io_ci = FullAdder_2863_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_126_io_a = FullAdder_2864_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_126_io_b = FullAdder_2865_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3228_io_a = FullAdder_2326_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3228_io_b = FullAdder_2862_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3228_io_ci = FullAdder_2863_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3229_io_a = FullAdder_2864_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3229_io_b = FullAdder_2865_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3229_io_ci = FullAdder_2866_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3230_io_a = FullAdder_2867_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3230_io_b = FullAdder_2868_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3230_io_ci = FullAdder_2869_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3231_io_a = FullAdder_2332_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3231_io_b = FullAdder_2866_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3231_io_ci = FullAdder_2867_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3232_io_a = FullAdder_2868_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3232_io_b = FullAdder_2869_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3232_io_ci = FullAdder_2870_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3233_io_a = FullAdder_2871_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3233_io_b = FullAdder_2872_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3233_io_ci = FullAdder_2873_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3234_io_a = FullAdder_2870_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3234_io_b = FullAdder_2871_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3234_io_ci = FullAdder_2872_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3235_io_a = FullAdder_2873_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3235_io_b = FullAdder_2874_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3235_io_ci = FullAdder_2875_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3236_io_a = FullAdder_2876_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3236_io_b = FullAdder_2877_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3236_io_ci = FullAdder_2878_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3237_io_a = FullAdder_2875_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3237_io_b = FullAdder_2876_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3237_io_ci = FullAdder_2877_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3238_io_a = FullAdder_2878_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3238_io_b = HalfAdder_101_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3238_io_ci = FullAdder_2879_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3239_io_a = FullAdder_2880_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3239_io_b = FullAdder_2881_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3239_io_ci = FullAdder_2882_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3240_io_a = FullAdder_2350_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3240_io_b = FullAdder_2879_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3240_io_ci = FullAdder_2880_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3241_io_a = FullAdder_2881_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3241_io_b = FullAdder_2882_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3241_io_ci = FullAdder_2883_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3242_io_a = FullAdder_2884_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3242_io_b = FullAdder_2885_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3242_io_ci = FullAdder_2886_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3243_io_a = FullAdder_2883_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3243_io_b = FullAdder_2884_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3243_io_ci = FullAdder_2885_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3244_io_a = FullAdder_2886_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3244_io_b = FullAdder_2887_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3244_io_ci = FullAdder_2888_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3245_io_a = FullAdder_2889_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3245_io_b = FullAdder_2890_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3245_io_ci = FullAdder_2891_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3246_io_a = FullAdder_2888_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3246_io_b = FullAdder_2889_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3246_io_ci = FullAdder_2890_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3247_io_a = FullAdder_2891_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3247_io_b = FullAdder_2892_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3247_io_ci = FullAdder_2893_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3248_io_a = FullAdder_2894_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3248_io_b = FullAdder_2895_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3248_io_ci = FullAdder_2896_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3249_io_a = FullAdder_2371_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3249_io_b = FullAdder_2893_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3249_io_ci = FullAdder_2894_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3250_io_a = FullAdder_2895_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3250_io_b = FullAdder_2896_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3250_io_ci = FullAdder_2897_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3251_io_a = FullAdder_2898_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3251_io_b = FullAdder_2899_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3251_io_ci = FullAdder_2900_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3252_io_a = FullAdder_2898_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3252_io_b = FullAdder_2899_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3252_io_ci = FullAdder_2900_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3253_io_a = FullAdder_2901_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3253_io_b = FullAdder_2902_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3253_io_ci = FullAdder_2903_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3254_io_a = FullAdder_2904_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3254_io_b = FullAdder_2905_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3254_io_ci = FullAdder_2906_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3255_io_a = FullAdder_2385_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3255_io_b = HalfAdder_77_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3255_io_ci = FullAdder_2903_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3256_io_a = FullAdder_2904_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3256_io_b = FullAdder_2905_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3256_io_ci = FullAdder_2906_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3257_io_a = FullAdder_2907_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3257_io_b = FullAdder_2908_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3257_io_ci = FullAdder_2909_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3258_io_a = FullAdder_2910_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3258_io_b = FullAdder_2911_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3258_io_ci = FullAdder_2912_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3259_io_a = FullAdder_2393_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3259_io_b = FullAdder_2908_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3259_io_ci = FullAdder_2909_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3260_io_a = FullAdder_2910_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3260_io_b = FullAdder_2911_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3260_io_ci = FullAdder_2912_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3261_io_a = FullAdder_2913_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3261_io_b = FullAdder_2914_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3261_io_ci = FullAdder_2915_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_127_io_a = FullAdder_2916_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_127_io_b = FullAdder_2917_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3262_io_a = FullAdder_2401_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3262_io_b = FullAdder_2913_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3262_io_ci = FullAdder_2914_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3263_io_a = FullAdder_2915_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3263_io_b = FullAdder_2916_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3263_io_ci = FullAdder_2917_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3264_io_a = FullAdder_2918_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3264_io_b = FullAdder_2919_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3264_io_ci = FullAdder_2920_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_128_io_a = FullAdder_2921_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_128_io_b = FullAdder_2922_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3265_io_a = FullAdder_2409_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3265_io_b = FullAdder_2918_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3265_io_ci = FullAdder_2919_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3266_io_a = FullAdder_2920_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3266_io_b = FullAdder_2921_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3266_io_ci = FullAdder_2922_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3267_io_a = FullAdder_2923_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3267_io_b = FullAdder_2924_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3267_io_ci = FullAdder_2925_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_129_io_a = FullAdder_2926_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_129_io_b = FullAdder_2927_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3268_io_a = FullAdder_2417_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3268_io_b = FullAdder_2923_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3268_io_ci = FullAdder_2924_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3269_io_a = FullAdder_2925_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3269_io_b = FullAdder_2926_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3269_io_ci = FullAdder_2927_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3270_io_a = FullAdder_2928_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3270_io_b = FullAdder_2929_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3270_io_ci = FullAdder_2930_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3271_io_a = FullAdder_2931_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3271_io_b = FullAdder_2932_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3271_io_ci = HalfAdder_102_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3272_io_a = FullAdder_2928_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3272_io_b = FullAdder_2929_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3272_io_ci = FullAdder_2930_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3273_io_a = FullAdder_2931_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3273_io_b = FullAdder_2932_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3273_io_ci = HalfAdder_102_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3274_io_a = FullAdder_2933_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3274_io_b = FullAdder_2934_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3274_io_ci = FullAdder_2935_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3275_io_a = FullAdder_2936_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3275_io_b = FullAdder_2937_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3275_io_ci = FullAdder_2938_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3276_io_a = FullAdder_2933_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3276_io_b = FullAdder_2934_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3276_io_ci = FullAdder_2935_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3277_io_a = FullAdder_2936_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3277_io_b = FullAdder_2937_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3277_io_ci = FullAdder_2938_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3278_io_a = FullAdder_2939_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3278_io_b = FullAdder_2940_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3278_io_ci = FullAdder_2941_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3279_io_a = FullAdder_2942_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3279_io_b = FullAdder_2943_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3279_io_ci = FullAdder_2944_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3280_io_a = FullAdder_2939_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3280_io_b = FullAdder_2940_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3280_io_ci = FullAdder_2941_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3281_io_a = FullAdder_2942_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3281_io_b = FullAdder_2943_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3281_io_ci = FullAdder_2944_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3282_io_a = FullAdder_2945_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3282_io_b = FullAdder_2946_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3282_io_ci = FullAdder_2947_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3283_io_a = FullAdder_2948_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3283_io_b = FullAdder_2949_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3283_io_ci = FullAdder_2950_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3284_io_a = FullAdder_2945_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3284_io_b = FullAdder_2946_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3284_io_ci = FullAdder_2947_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3285_io_a = FullAdder_2948_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3285_io_b = FullAdder_2949_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3285_io_ci = FullAdder_2950_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3286_io_a = FullAdder_2951_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3286_io_b = FullAdder_2952_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3286_io_ci = FullAdder_2953_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3287_io_a = FullAdder_2954_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3287_io_b = FullAdder_2955_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3287_io_ci = FullAdder_2956_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3288_io_a = FullAdder_2951_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3288_io_b = FullAdder_2952_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3288_io_ci = FullAdder_2953_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3289_io_a = FullAdder_2954_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3289_io_b = FullAdder_2955_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3289_io_ci = FullAdder_2956_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3290_io_a = FullAdder_2957_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3290_io_b = FullAdder_2958_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3290_io_ci = FullAdder_2959_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3291_io_a = FullAdder_2960_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3291_io_b = FullAdder_2961_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3291_io_ci = FullAdder_2962_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3292_io_a = FullAdder_2957_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3292_io_b = FullAdder_2958_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3292_io_ci = FullAdder_2959_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3293_io_a = FullAdder_2960_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3293_io_b = FullAdder_2961_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3293_io_ci = FullAdder_2962_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3294_io_a = FullAdder_2963_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3294_io_b = FullAdder_2964_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3294_io_ci = FullAdder_2965_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3295_io_a = FullAdder_2966_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3295_io_b = FullAdder_2967_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3295_io_ci = FullAdder_2968_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3296_io_a = FullAdder_2478_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3296_io_b = FullAdder_2963_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3296_io_ci = FullAdder_2964_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3297_io_a = FullAdder_2965_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3297_io_b = FullAdder_2966_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3297_io_ci = FullAdder_2967_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3298_io_a = FullAdder_2968_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3298_io_b = FullAdder_2969_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3298_io_ci = FullAdder_2970_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3299_io_a = FullAdder_2971_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3299_io_b = FullAdder_2972_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3299_io_ci = FullAdder_2973_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3300_io_a = FullAdder_2487_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3300_io_b = FullAdder_2969_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3300_io_ci = FullAdder_2970_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3301_io_a = FullAdder_2971_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3301_io_b = FullAdder_2972_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3301_io_ci = FullAdder_2973_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3302_io_a = FullAdder_2974_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3302_io_b = FullAdder_2975_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3302_io_ci = FullAdder_2976_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3303_io_a = FullAdder_2977_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3303_io_b = FullAdder_2978_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3303_io_ci = FullAdder_2979_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3304_io_a = FullAdder_2496_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3304_io_b = FullAdder_2975_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3304_io_ci = FullAdder_2976_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3305_io_a = FullAdder_2977_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3305_io_b = FullAdder_2978_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3305_io_ci = FullAdder_2979_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3306_io_a = FullAdder_2980_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3306_io_b = FullAdder_2981_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3306_io_ci = FullAdder_2982_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3307_io_a = FullAdder_2983_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3307_io_b = FullAdder_2984_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3307_io_ci = FullAdder_2985_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_130_io_a = FullAdder_2986_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_130_io_b = HalfAdder_103_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3308_io_a = FullAdder_2981_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3308_io_b = FullAdder_2982_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3308_io_ci = FullAdder_2983_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3309_io_a = FullAdder_2984_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3309_io_b = FullAdder_2985_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3309_io_ci = FullAdder_2986_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3310_io_a = HalfAdder_103_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3310_io_b = FullAdder_2987_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3310_io_ci = FullAdder_2988_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3311_io_a = FullAdder_2989_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3311_io_b = FullAdder_2990_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3311_io_ci = FullAdder_2991_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3312_io_a = FullAdder_2514_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3312_io_b = FullAdder_2987_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3312_io_ci = FullAdder_2988_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3313_io_a = FullAdder_2989_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3313_io_b = FullAdder_2990_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3313_io_ci = FullAdder_2991_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3314_io_a = FullAdder_2992_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3314_io_b = FullAdder_2993_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3314_io_ci = FullAdder_2994_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3315_io_a = FullAdder_2995_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3315_io_b = FullAdder_2996_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3315_io_ci = FullAdder_2997_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3316_io_a = FullAdder_2523_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3316_io_b = FullAdder_2993_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3316_io_ci = FullAdder_2994_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3317_io_a = FullAdder_2995_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3317_io_b = FullAdder_2996_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3317_io_ci = FullAdder_2997_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3318_io_a = FullAdder_2998_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3318_io_b = FullAdder_2999_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3318_io_ci = FullAdder_3000_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3319_io_a = FullAdder_3001_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3319_io_b = FullAdder_3002_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3319_io_ci = FullAdder_3003_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3320_io_a = FullAdder_2999_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3320_io_b = FullAdder_3000_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3320_io_ci = FullAdder_3001_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3321_io_a = FullAdder_3002_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3321_io_b = FullAdder_3003_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3321_io_ci = FullAdder_3004_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3322_io_a = FullAdder_3005_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3322_io_b = FullAdder_3006_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3322_io_ci = FullAdder_3007_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3323_io_a = FullAdder_3008_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3323_io_b = FullAdder_3009_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3323_io_ci = FullAdder_3010_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3324_io_a = FullAdder_2541_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3324_io_b = FullAdder_3005_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3324_io_ci = FullAdder_3006_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3325_io_a = FullAdder_3007_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3325_io_b = FullAdder_3008_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3325_io_ci = FullAdder_3009_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3326_io_a = FullAdder_3010_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3326_io_b = FullAdder_3011_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3326_io_ci = FullAdder_3012_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3327_io_a = FullAdder_3013_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3327_io_b = FullAdder_3014_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3327_io_ci = FullAdder_3015_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3328_io_a = FullAdder_3011_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3328_io_b = FullAdder_3012_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3328_io_ci = FullAdder_3013_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3329_io_a = FullAdder_3014_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3329_io_b = FullAdder_3015_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3329_io_ci = FullAdder_3016_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3330_io_a = FullAdder_3017_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3330_io_b = FullAdder_3018_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3330_io_ci = FullAdder_3019_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3331_io_a = FullAdder_2556_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3331_io_b = FullAdder_2557_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3331_io_ci = FullAdder_3017_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3332_io_a = FullAdder_3018_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3332_io_b = FullAdder_3019_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3332_io_ci = FullAdder_3020_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3333_io_a = FullAdder_3021_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3333_io_b = FullAdder_3022_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3333_io_ci = FullAdder_3023_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3334_io_a = FullAdder_3024_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3334_io_b = FullAdder_3025_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3334_io_ci = FullAdder_3026_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3335_io_a = FullAdder_3022_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3335_io_b = FullAdder_3023_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3335_io_ci = FullAdder_3024_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3336_io_a = FullAdder_3025_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3336_io_b = FullAdder_3026_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3336_io_ci = HalfAdder_104_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3337_io_a = FullAdder_3027_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3337_io_b = FullAdder_3028_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3337_io_ci = FullAdder_3029_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3338_io_a = FullAdder_3030_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3338_io_b = FullAdder_3031_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3338_io_ci = HalfAdder_105_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3339_io_a = FullAdder_3027_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3339_io_b = FullAdder_3028_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3339_io_ci = FullAdder_3029_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3340_io_a = FullAdder_3030_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3340_io_b = FullAdder_3031_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3340_io_ci = HalfAdder_105_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3341_io_a = FullAdder_3032_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3341_io_b = FullAdder_3033_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3341_io_ci = FullAdder_3034_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3342_io_a = FullAdder_3035_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3342_io_b = FullAdder_3036_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3342_io_ci = FullAdder_3037_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3343_io_a = FullAdder_3032_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3343_io_b = FullAdder_3033_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3343_io_ci = FullAdder_3034_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3344_io_a = FullAdder_3035_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3344_io_b = FullAdder_3036_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3344_io_ci = FullAdder_3037_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3345_io_a = FullAdder_3038_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3345_io_b = FullAdder_3039_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3345_io_ci = FullAdder_3040_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3346_io_a = FullAdder_2588_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3346_io_b = FullAdder_3038_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3346_io_ci = FullAdder_3039_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3347_io_a = FullAdder_3040_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3347_io_b = FullAdder_3041_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3347_io_ci = FullAdder_3042_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3348_io_a = FullAdder_3043_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3348_io_b = FullAdder_3044_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3348_io_ci = FullAdder_3045_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_131_io_a = FullAdder_3046_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_131_io_b = FullAdder_3047_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3349_io_a = FullAdder_2595_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3349_io_b = FullAdder_2596_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3349_io_ci = FullAdder_3043_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3350_io_a = FullAdder_3044_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3350_io_b = FullAdder_3045_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3350_io_ci = FullAdder_3046_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3351_io_a = FullAdder_3047_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3351_io_b = FullAdder_3048_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3351_io_ci = FullAdder_3049_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3352_io_a = FullAdder_3050_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3352_io_b = FullAdder_3051_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3352_io_ci = FullAdder_3052_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3353_io_a = FullAdder_2603_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3353_io_b = HalfAdder_80_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3353_io_ci = FullAdder_3048_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3354_io_a = FullAdder_3049_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3354_io_b = FullAdder_3050_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3354_io_ci = FullAdder_3051_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3355_io_a = FullAdder_3052_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3355_io_b = FullAdder_3053_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3355_io_ci = FullAdder_3054_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3356_io_a = FullAdder_3055_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3356_io_b = FullAdder_3056_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3356_io_ci = FullAdder_3057_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3357_io_a = FullAdder_3053_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3357_io_b = FullAdder_3054_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3357_io_ci = FullAdder_3055_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3358_io_a = FullAdder_3056_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3358_io_b = FullAdder_3057_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3358_io_ci = FullAdder_3058_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3359_io_a = FullAdder_3059_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3359_io_b = FullAdder_3060_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3359_io_ci = FullAdder_3061_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3360_io_a = FullAdder_3058_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3360_io_b = FullAdder_3059_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3360_io_ci = FullAdder_3060_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3361_io_a = FullAdder_3061_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3361_io_b = FullAdder_3062_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3361_io_ci = FullAdder_3063_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3362_io_a = FullAdder_3064_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3362_io_b = FullAdder_3065_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3362_io_ci = FullAdder_3066_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3363_io_a = FullAdder_2624_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3363_io_b = FullAdder_3063_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3363_io_ci = FullAdder_3064_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3364_io_a = FullAdder_3065_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3364_io_b = FullAdder_3066_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3364_io_ci = FullAdder_3067_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3365_io_a = FullAdder_3068_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3365_io_b = FullAdder_3069_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3365_io_ci = FullAdder_3070_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3366_io_a = FullAdder_3068_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3366_io_b = FullAdder_3069_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3366_io_ci = FullAdder_3070_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3367_io_a = FullAdder_3071_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3367_io_b = FullAdder_3072_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3367_io_ci = FullAdder_3073_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3368_io_a = FullAdder_3074_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3368_io_b = FullAdder_3075_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3368_io_ci = FullAdder_3076_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3369_io_a = FullAdder_3073_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3369_io_b = FullAdder_3074_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3369_io_ci = FullAdder_3075_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3370_io_a = FullAdder_3076_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3370_io_b = HalfAdder_106_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3370_io_ci = FullAdder_3077_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3371_io_a = FullAdder_3078_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3371_io_b = FullAdder_3079_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3371_io_ci = FullAdder_3080_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3372_io_a = FullAdder_2644_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3372_io_b = HalfAdder_81_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3372_io_ci = FullAdder_3077_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3373_io_a = FullAdder_3078_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3373_io_b = FullAdder_3079_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3373_io_ci = FullAdder_3080_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3374_io_a = FullAdder_3081_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3374_io_b = FullAdder_3082_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3374_io_ci = FullAdder_3083_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3375_io_a = FullAdder_2650_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3375_io_b = FullAdder_2651_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3375_io_ci = FullAdder_3081_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3376_io_a = FullAdder_3082_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3376_io_b = FullAdder_3083_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3376_io_ci = FullAdder_3084_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3377_io_a = FullAdder_3085_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3377_io_b = FullAdder_3086_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3377_io_ci = FullAdder_3087_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3378_io_a = FullAdder_2657_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3378_io_b = FullAdder_3085_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3378_io_ci = FullAdder_3086_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3379_io_a = FullAdder_3087_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3379_io_b = FullAdder_3088_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3379_io_ci = FullAdder_3089_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3380_io_a = FullAdder_3090_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3380_io_b = FullAdder_3091_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3380_io_ci = FullAdder_3092_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3381_io_a = FullAdder_2662_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3381_io_b = FullAdder_2663_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3381_io_ci = FullAdder_3089_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3382_io_a = FullAdder_3090_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3382_io_b = FullAdder_3091_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3382_io_ci = FullAdder_3092_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3383_io_a = FullAdder_3093_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3383_io_b = FullAdder_3094_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3383_io_ci = FullAdder_3095_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3384_io_a = FullAdder_2669_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3384_io_b = FullAdder_3093_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3384_io_ci = FullAdder_3094_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3385_io_a = FullAdder_3095_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3385_io_b = FullAdder_3096_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3385_io_ci = FullAdder_3097_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3386_io_a = FullAdder_3098_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3386_io_b = FullAdder_3099_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3386_io_ci = FullAdder_3100_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3387_io_a = FullAdder_3097_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3387_io_b = FullAdder_3098_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3387_io_ci = FullAdder_3099_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3388_io_a = FullAdder_3100_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3388_io_b = FullAdder_3101_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3388_io_ci = FullAdder_3102_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_132_io_a = FullAdder_3103_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_132_io_b = FullAdder_3104_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3389_io_a = FullAdder_2681_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3389_io_b = FullAdder_3101_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3389_io_ci = FullAdder_3102_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3390_io_a = FullAdder_3103_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3390_io_b = FullAdder_3104_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3390_io_ci = FullAdder_3105_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3391_io_a = FullAdder_2685_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3391_io_b = FullAdder_2686_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3391_io_ci = FullAdder_3105_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3392_io_a = FullAdder_3106_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3392_io_b = FullAdder_3107_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3392_io_ci = FullAdder_3108_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3393_io_a = FullAdder_3109_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3393_io_b = FullAdder_3110_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3393_io_ci = FullAdder_3111_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3394_io_a = HalfAdder_82_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3394_io_b = FullAdder_3108_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3394_io_ci = FullAdder_3109_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3395_io_a = FullAdder_3110_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3395_io_b = FullAdder_3111_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3395_io_ci = FullAdder_3112_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3396_io_a = FullAdder_3113_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3396_io_b = FullAdder_3114_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3396_io_ci = FullAdder_3115_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3397_io_a = FullAdder_3112_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3397_io_b = FullAdder_3113_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3397_io_ci = FullAdder_3114_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3398_io_a = FullAdder_3115_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3398_io_b = FullAdder_3116_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3398_io_ci = FullAdder_3117_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3399_io_a = FullAdder_3116_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3399_io_b = FullAdder_3117_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3399_io_ci = FullAdder_3118_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3400_io_a = HalfAdder_107_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3400_io_b = FullAdder_3119_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3400_io_ci = FullAdder_3120_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3401_io_a = FullAdder_2706_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3401_io_b = FullAdder_3119_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3401_io_ci = FullAdder_3120_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3402_io_a = FullAdder_3121_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3402_io_b = FullAdder_3122_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3402_io_ci = FullAdder_3123_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_133_io_a = FullAdder_3124_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_133_io_b = FullAdder_3125_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3403_io_a = FullAdder_3122_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3403_io_b = FullAdder_3123_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3403_io_ci = FullAdder_3124_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3404_io_a = FullAdder_3125_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3404_io_b = FullAdder_3126_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3404_io_ci = FullAdder_3127_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3405_io_a = FullAdder_2716_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3405_io_b = FullAdder_3126_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3405_io_ci = FullAdder_3127_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3406_io_a = FullAdder_3128_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3406_io_b = FullAdder_3129_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3406_io_ci = FullAdder_3130_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3407_io_a = FullAdder_3129_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3407_io_b = FullAdder_3130_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3407_io_ci = FullAdder_3131_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3408_io_a = FullAdder_3132_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3408_io_b = FullAdder_3133_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3408_io_ci = FullAdder_3134_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3409_io_a = FullAdder_2724_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3409_io_b = HalfAdder_84_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3409_io_ci = FullAdder_3132_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3410_io_a = FullAdder_3133_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3410_io_b = FullAdder_3134_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3410_io_ci = FullAdder_3135_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3411_io_a = FullAdder_3135_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3411_io_b = FullAdder_3136_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3411_io_ci = FullAdder_3137_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3412_io_a = FullAdder_3138_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3412_io_b = FullAdder_3139_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3412_io_ci = FullAdder_3140_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3413_io_a = FullAdder_3138_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3413_io_b = FullAdder_3139_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3413_io_ci = FullAdder_3140_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3414_io_a = FullAdder_3141_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3414_io_b = FullAdder_3142_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3414_io_ci = FullAdder_3143_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3415_io_a = FullAdder_3141_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3415_io_b = FullAdder_3142_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3415_io_ci = FullAdder_3143_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3416_io_a = FullAdder_3144_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3416_io_b = FullAdder_3145_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3416_io_ci = FullAdder_3146_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3417_io_a = FullAdder_3144_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3417_io_b = FullAdder_3145_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3417_io_ci = FullAdder_3146_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3418_io_a = FullAdder_2743_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3418_io_b = FullAdder_3147_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3418_io_ci = FullAdder_3148_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3419_io_a = FullAdder_3149_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3419_io_b = FullAdder_3150_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3419_io_ci = FullAdder_3151_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3420_io_a = FullAdder_3149_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3420_io_b = FullAdder_3150_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3420_io_ci = FullAdder_3151_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3421_io_a = FullAdder_2750_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3421_io_b = HalfAdder_85_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3421_io_ci = FullAdder_3152_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3422_io_a = FullAdder_3153_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3422_io_b = FullAdder_3154_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3422_io_ci = FullAdder_3155_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3423_io_a = FullAdder_2753_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3423_io_b = FullAdder_3154_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3423_io_ci = FullAdder_3155_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_134_io_a = FullAdder_3156_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_134_io_b = FullAdder_3157_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3424_io_a = FullAdder_2756_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3424_io_b = FullAdder_3156_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3424_io_ci = FullAdder_3157_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_135_io_a = FullAdder_3158_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_135_io_b = FullAdder_3159_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3425_io_a = FullAdder_2759_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3425_io_b = FullAdder_3158_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3425_io_ci = FullAdder_3159_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_136_io_a = FullAdder_3160_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_136_io_b = FullAdder_3161_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3426_io_a = FullAdder_3160_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3426_io_b = FullAdder_3161_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3426_io_ci = FullAdder_3162_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3427_io_a = FullAdder_3162_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3427_io_b = FullAdder_3163_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3427_io_ci = FullAdder_3164_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3428_io_a = FullAdder_2766_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3428_io_b = FullAdder_2767_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3428_io_ci = FullAdder_3164_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3429_io_a = HalfAdder_86_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3429_io_b = FullAdder_3165_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3429_io_ci = FullAdder_3166_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3430_io_a = FullAdder_3167_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3430_io_b = HalfAdder_108_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3430_io_ci = FullAdder_3168_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3431_io_a = FullAdder_2772_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3431_io_b = FullAdder_2773_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3431_io_ci = FullAdder_3168_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3432_io_a = FullAdder_3169_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3432_io_b = HalfAdder_109_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3432_io_ci = FullAdder_3170_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3433_io_a = FullAdder_2777_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3433_io_b = FullAdder_2778_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3433_io_ci = FullAdder_3171_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3434_io_a = HalfAdder_87_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3434_io_b = HalfAdder_88_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3434_io_ci = FullAdder_3172_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_137_io_a = HalfAdder_89_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_137_io_b = HalfAdder_110_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_138_io_a = HalfAdder_111_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_138_io_b = FullAdder_3173_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_139_io_a = FullAdder_3174_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_139_io_b = FullAdder_3175_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_140_io_a = FullAdder_3175_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_140_io_b = HalfAdder_112_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_141_io_a = HalfAdder_112_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_141_io_b = HalfAdder_113_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_142_io_a = HalfAdder_113_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_142_io_b = HalfAdder_114_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_143_io_a = HalfAdder_91_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_143_io_b = HalfAdder_114_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_144_io_a = HalfAdder_93_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_144_io_b = FullAdder_3176_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_145_io_a = HalfAdder_95_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_145_io_b = HalfAdder_116_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_146_io_a = HalfAdder_117_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_146_io_b = FullAdder_3177_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_147_io_a = FullAdder_3177_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_147_io_b = HalfAdder_118_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_148_io_a = FullAdder_2785_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_148_io_b = HalfAdder_118_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_149_io_a = FullAdder_3178_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_149_io_b = FullAdder_3179_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3435_io_a = FullAdder_2788_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3435_io_b = FullAdder_3179_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3435_io_ci = FullAdder_3180_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_150_io_a = FullAdder_3181_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_150_io_b = FullAdder_3182_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3436_io_a = FullAdder_2792_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3436_io_b = FullAdder_3182_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3436_io_ci = FullAdder_3183_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3437_io_a = FullAdder_2793_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3437_io_b = FullAdder_3183_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3437_io_ci = FullAdder_3184_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3438_io_a = FullAdder_2794_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3438_io_b = FullAdder_2795_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3438_io_ci = FullAdder_3184_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3439_io_a = FullAdder_2796_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3439_io_b = FullAdder_2797_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3439_io_ci = FullAdder_3185_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3440_io_a = FullAdder_2799_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3440_io_b = FullAdder_3186_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3440_io_ci = FullAdder_3187_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3441_io_a = FullAdder_2801_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3441_io_b = FullAdder_3187_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3441_io_ci = FullAdder_3188_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3442_io_a = FullAdder_3188_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3442_io_b = HalfAdder_120_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3442_io_ci = FullAdder_3189_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3443_io_a = FullAdder_3189_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3443_io_b = HalfAdder_121_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3443_io_ci = FullAdder_3190_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3444_io_a = FullAdder_3190_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3444_io_b = FullAdder_3191_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3444_io_ci = FullAdder_3192_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3445_io_a = FullAdder_2809_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3445_io_b = FullAdder_2810_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3445_io_ci = FullAdder_3192_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3446_io_a = FullAdder_3193_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3446_io_b = FullAdder_3194_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3446_io_ci = FullAdder_3195_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3447_io_a = FullAdder_3195_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3447_io_b = FullAdder_3196_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3447_io_ci = FullAdder_3197_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3448_io_a = FullAdder_3197_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3448_io_b = FullAdder_3198_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3448_io_ci = FullAdder_3199_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3449_io_a = FullAdder_3199_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3449_io_b = FullAdder_3200_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3449_io_ci = FullAdder_3201_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_151_io_a = FullAdder_3201_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_151_io_b = FullAdder_3202_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_152_io_a = FullAdder_3203_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_152_io_b = FullAdder_3204_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3450_io_a = FullAdder_2827_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3450_io_b = FullAdder_3203_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3450_io_ci = FullAdder_3204_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3451_io_a = FullAdder_2830_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3451_io_b = FullAdder_3205_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3451_io_ci = FullAdder_3206_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3452_io_a = FullAdder_2832_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3452_io_b = FullAdder_2833_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3452_io_ci = FullAdder_3207_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3453_io_a = FullAdder_3208_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3453_io_b = FullAdder_3209_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3453_io_ci = FullAdder_3210_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3454_io_a = FullAdder_2836_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3454_io_b = FullAdder_3209_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3454_io_ci = FullAdder_3210_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_153_io_a = FullAdder_3211_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_153_io_b = FullAdder_3212_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3455_io_a = FullAdder_2839_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3455_io_b = HalfAdder_98_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3455_io_ci = FullAdder_3211_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3456_io_a = FullAdder_3212_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3456_io_b = FullAdder_3213_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3456_io_ci = FullAdder_3214_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3457_io_a = FullAdder_3213_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3457_io_b = FullAdder_3214_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3457_io_ci = HalfAdder_122_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3458_io_a = FullAdder_3215_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3458_io_b = FullAdder_3216_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3458_io_ci = HalfAdder_123_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3459_io_a = FullAdder_3215_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3459_io_b = FullAdder_3216_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3459_io_ci = HalfAdder_123_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_154_io_a = FullAdder_3217_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_154_io_b = FullAdder_3218_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3460_io_a = FullAdder_3217_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3460_io_b = FullAdder_3218_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3460_io_ci = HalfAdder_124_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3461_io_a = FullAdder_3219_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3461_io_b = FullAdder_3220_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3461_io_ci = FullAdder_3221_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3462_io_a = FullAdder_3219_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3462_io_b = FullAdder_3220_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3462_io_ci = FullAdder_3221_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3463_io_a = FullAdder_2856_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3463_io_b = FullAdder_2857_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3463_io_ci = FullAdder_3222_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3464_io_a = FullAdder_3223_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3464_io_b = FullAdder_3224_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3464_io_ci = FullAdder_3225_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3465_io_a = FullAdder_3224_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3465_io_b = FullAdder_3225_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3465_io_ci = HalfAdder_125_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3466_io_a = FullAdder_3226_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3466_io_b = FullAdder_3227_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3466_io_ci = HalfAdder_126_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_155_io_a = FullAdder_3226_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_155_io_b = FullAdder_3227_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_156_io_a = HalfAdder_126_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_156_io_b = FullAdder_3228_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_157_io_a = FullAdder_3229_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_157_io_b = FullAdder_3230_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3467_io_a = FullAdder_3228_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3467_io_b = FullAdder_3229_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3467_io_ci = FullAdder_3230_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3468_io_a = FullAdder_3231_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3468_io_b = FullAdder_3232_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3468_io_ci = FullAdder_3233_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3469_io_a = FullAdder_2874_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3469_io_b = FullAdder_3231_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3469_io_ci = FullAdder_3232_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3470_io_a = FullAdder_3233_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3470_io_b = FullAdder_3234_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3470_io_ci = FullAdder_3235_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3471_io_a = HalfAdder_101_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3471_io_b = FullAdder_3234_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3471_io_ci = FullAdder_3235_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3472_io_a = FullAdder_3236_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3472_io_b = FullAdder_3237_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3472_io_ci = FullAdder_3238_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3473_io_a = FullAdder_3237_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3473_io_b = FullAdder_3238_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3473_io_ci = FullAdder_3239_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3474_io_a = FullAdder_3240_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3474_io_b = FullAdder_3241_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3474_io_ci = FullAdder_3242_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3475_io_a = FullAdder_2887_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3475_io_b = FullAdder_3240_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3475_io_ci = FullAdder_3241_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3476_io_a = FullAdder_3242_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3476_io_b = FullAdder_3243_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3476_io_ci = FullAdder_3244_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3477_io_a = FullAdder_2892_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3477_io_b = FullAdder_3243_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3477_io_ci = FullAdder_3244_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3478_io_a = FullAdder_3245_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3478_io_b = FullAdder_3246_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3478_io_ci = FullAdder_3247_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3479_io_a = FullAdder_2897_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3479_io_b = FullAdder_3246_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3479_io_ci = FullAdder_3247_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3480_io_a = FullAdder_3248_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3480_io_b = FullAdder_3249_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3480_io_ci = FullAdder_3250_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3481_io_a = FullAdder_2901_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3481_io_b = FullAdder_2902_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3481_io_ci = FullAdder_3249_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3482_io_a = FullAdder_3250_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3482_io_b = FullAdder_3251_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3482_io_ci = FullAdder_3252_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3483_io_a = FullAdder_2907_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3483_io_b = FullAdder_3252_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3483_io_ci = FullAdder_3253_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3484_io_a = FullAdder_3254_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3484_io_b = FullAdder_3255_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3484_io_ci = FullAdder_3256_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_158_io_a = FullAdder_3257_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_158_io_b = FullAdder_3258_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3485_io_a = FullAdder_3255_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3485_io_b = FullAdder_3256_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3485_io_ci = FullAdder_3257_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3486_io_a = FullAdder_3258_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3486_io_b = FullAdder_3259_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3486_io_ci = FullAdder_3260_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3487_io_a = FullAdder_3259_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3487_io_b = FullAdder_3260_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3487_io_ci = FullAdder_3261_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3488_io_a = HalfAdder_127_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3488_io_b = FullAdder_3262_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3488_io_ci = FullAdder_3263_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3489_io_a = FullAdder_3262_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3489_io_b = FullAdder_3263_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3489_io_ci = FullAdder_3264_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3490_io_a = HalfAdder_128_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3490_io_b = FullAdder_3265_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3490_io_ci = FullAdder_3266_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_159_io_a = FullAdder_3267_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_159_io_b = HalfAdder_129_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3491_io_a = FullAdder_3265_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3491_io_b = FullAdder_3266_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3491_io_ci = FullAdder_3267_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3492_io_a = HalfAdder_129_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3492_io_b = FullAdder_3268_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3492_io_ci = FullAdder_3269_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3493_io_a = FullAdder_3268_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3493_io_b = FullAdder_3269_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3493_io_ci = FullAdder_3270_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3494_io_a = FullAdder_3271_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3494_io_b = FullAdder_3272_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3494_io_ci = FullAdder_3273_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_160_io_a = FullAdder_3274_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_160_io_b = FullAdder_3275_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3495_io_a = FullAdder_3272_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3495_io_b = FullAdder_3273_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3495_io_ci = FullAdder_3274_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3496_io_a = FullAdder_3275_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3496_io_b = FullAdder_3276_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3496_io_ci = FullAdder_3277_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_161_io_a = FullAdder_3278_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_161_io_b = FullAdder_3279_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3497_io_a = FullAdder_3276_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3497_io_b = FullAdder_3277_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3497_io_ci = FullAdder_3278_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3498_io_a = FullAdder_3279_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3498_io_b = FullAdder_3280_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3498_io_ci = FullAdder_3281_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3499_io_a = FullAdder_3280_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3499_io_b = FullAdder_3281_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3499_io_ci = FullAdder_3282_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3500_io_a = FullAdder_3283_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3500_io_b = FullAdder_3284_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3500_io_ci = FullAdder_3285_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3501_io_a = FullAdder_3284_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3501_io_b = FullAdder_3285_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3501_io_ci = FullAdder_3286_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3502_io_a = FullAdder_3287_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3502_io_b = FullAdder_3288_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3502_io_ci = FullAdder_3289_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3503_io_a = FullAdder_3288_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3503_io_b = FullAdder_3289_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3503_io_ci = FullAdder_3290_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3504_io_a = FullAdder_3291_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3504_io_b = FullAdder_3292_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3504_io_ci = FullAdder_3293_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_162_io_a = FullAdder_3294_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_162_io_b = FullAdder_3295_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3505_io_a = FullAdder_3292_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3505_io_b = FullAdder_3293_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3505_io_ci = FullAdder_3294_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3506_io_a = FullAdder_3295_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3506_io_b = FullAdder_3296_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3506_io_ci = FullAdder_3297_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_163_io_a = FullAdder_3298_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_163_io_b = FullAdder_3299_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3507_io_a = FullAdder_2974_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3507_io_b = FullAdder_3296_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3507_io_ci = FullAdder_3297_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_164_io_a = FullAdder_3298_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_164_io_b = FullAdder_3299_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_165_io_a = FullAdder_3300_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_165_io_b = FullAdder_3301_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_166_io_a = FullAdder_3302_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_166_io_b = FullAdder_3303_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3508_io_a = FullAdder_2980_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3508_io_b = FullAdder_3300_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3508_io_ci = FullAdder_3301_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3509_io_a = FullAdder_3302_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3509_io_b = FullAdder_3303_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3509_io_ci = FullAdder_3304_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3510_io_a = FullAdder_3305_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3510_io_b = FullAdder_3306_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3510_io_ci = FullAdder_3307_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3511_io_a = FullAdder_3304_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3511_io_b = FullAdder_3305_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3511_io_ci = FullAdder_3306_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3512_io_a = FullAdder_3307_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3512_io_b = HalfAdder_130_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3512_io_ci = FullAdder_3308_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3513_io_a = FullAdder_3309_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3513_io_b = FullAdder_3310_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3513_io_ci = FullAdder_3311_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3514_io_a = FullAdder_2992_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3514_io_b = FullAdder_3308_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3514_io_ci = FullAdder_3309_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3515_io_a = FullAdder_3310_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3515_io_b = FullAdder_3311_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3515_io_ci = FullAdder_3312_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3516_io_a = FullAdder_3313_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3516_io_b = FullAdder_3314_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3516_io_ci = FullAdder_3315_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3517_io_a = FullAdder_2998_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3517_io_b = FullAdder_3312_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3517_io_ci = FullAdder_3313_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3518_io_a = FullAdder_3314_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3518_io_b = FullAdder_3315_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3518_io_ci = FullAdder_3316_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3519_io_a = FullAdder_3317_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3519_io_b = FullAdder_3318_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3519_io_ci = FullAdder_3319_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3520_io_a = FullAdder_3004_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3520_io_b = FullAdder_3316_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3520_io_ci = FullAdder_3317_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3521_io_a = FullAdder_3318_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3521_io_b = FullAdder_3319_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3521_io_ci = FullAdder_3320_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3522_io_a = FullAdder_3321_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3522_io_b = FullAdder_3322_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3522_io_ci = FullAdder_3323_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3523_io_a = FullAdder_3320_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3523_io_b = FullAdder_3321_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3523_io_ci = FullAdder_3322_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3524_io_a = FullAdder_3323_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3524_io_b = FullAdder_3324_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3524_io_ci = FullAdder_3325_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3525_io_a = FullAdder_3016_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3525_io_b = FullAdder_3324_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3525_io_ci = FullAdder_3325_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3526_io_a = FullAdder_3326_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3526_io_b = FullAdder_3327_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3526_io_ci = FullAdder_3328_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3527_io_a = FullAdder_3020_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3527_io_b = FullAdder_3021_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3527_io_ci = FullAdder_3328_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3528_io_a = FullAdder_3329_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3528_io_b = FullAdder_3330_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3528_io_ci = FullAdder_3331_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3529_io_a = FullAdder_3332_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3529_io_b = FullAdder_3333_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3529_io_ci = FullAdder_3334_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3530_io_a = HalfAdder_104_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3530_io_b = FullAdder_3331_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3530_io_ci = FullAdder_3332_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3531_io_a = FullAdder_3333_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3531_io_b = FullAdder_3334_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3531_io_ci = FullAdder_3335_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3532_io_a = FullAdder_3336_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3532_io_b = FullAdder_3337_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3532_io_ci = FullAdder_3338_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3533_io_a = FullAdder_3335_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3533_io_b = FullAdder_3336_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3533_io_ci = FullAdder_3337_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3534_io_a = FullAdder_3338_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3534_io_b = FullAdder_3339_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3534_io_ci = FullAdder_3340_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_167_io_a = FullAdder_3341_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_167_io_b = FullAdder_3342_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3535_io_a = FullAdder_3339_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3535_io_b = FullAdder_3340_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3535_io_ci = FullAdder_3341_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3536_io_a = FullAdder_3342_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3536_io_b = FullAdder_3343_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3536_io_ci = FullAdder_3344_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3537_io_a = FullAdder_3041_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3537_io_b = FullAdder_3042_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3537_io_ci = FullAdder_3343_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3538_io_a = FullAdder_3344_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3538_io_b = FullAdder_3345_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3538_io_ci = FullAdder_3346_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3539_io_a = FullAdder_3347_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3539_io_b = FullAdder_3348_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3539_io_ci = HalfAdder_131_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3540_io_a = FullAdder_3346_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3540_io_b = FullAdder_3347_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3540_io_ci = FullAdder_3348_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3541_io_a = HalfAdder_131_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3541_io_b = FullAdder_3349_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3541_io_ci = FullAdder_3350_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3542_io_a = FullAdder_3349_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3542_io_b = FullAdder_3350_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3542_io_ci = FullAdder_3351_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3543_io_a = FullAdder_3352_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3543_io_b = FullAdder_3353_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3543_io_ci = FullAdder_3354_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3544_io_a = FullAdder_3353_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3544_io_b = FullAdder_3354_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3544_io_ci = FullAdder_3355_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3545_io_a = FullAdder_3356_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3545_io_b = FullAdder_3357_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3545_io_ci = FullAdder_3358_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3546_io_a = FullAdder_3062_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3546_io_b = FullAdder_3357_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3546_io_ci = FullAdder_3358_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3547_io_a = FullAdder_3359_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3547_io_b = FullAdder_3360_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3547_io_ci = FullAdder_3361_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3548_io_a = FullAdder_3067_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3548_io_b = FullAdder_3360_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3548_io_ci = FullAdder_3361_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3549_io_a = FullAdder_3362_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3549_io_b = FullAdder_3363_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3549_io_ci = FullAdder_3364_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3550_io_a = FullAdder_3071_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3550_io_b = FullAdder_3072_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3550_io_ci = FullAdder_3363_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3551_io_a = FullAdder_3364_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3551_io_b = FullAdder_3365_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3551_io_ci = FullAdder_3366_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3552_io_a = HalfAdder_106_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3552_io_b = FullAdder_3366_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3552_io_ci = FullAdder_3367_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3553_io_a = FullAdder_3368_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3553_io_b = FullAdder_3369_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3553_io_ci = FullAdder_3370_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3554_io_a = FullAdder_3369_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3554_io_b = FullAdder_3370_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3554_io_ci = FullAdder_3371_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3555_io_a = FullAdder_3372_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3555_io_b = FullAdder_3373_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3555_io_ci = FullAdder_3374_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3556_io_a = FullAdder_3084_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3556_io_b = FullAdder_3372_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3556_io_ci = FullAdder_3373_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3557_io_a = FullAdder_3374_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3557_io_b = FullAdder_3375_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3557_io_ci = FullAdder_3376_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3558_io_a = FullAdder_3088_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3558_io_b = FullAdder_3375_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3558_io_ci = FullAdder_3376_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3559_io_a = FullAdder_3377_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3559_io_b = FullAdder_3378_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3559_io_ci = FullAdder_3379_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3560_io_a = FullAdder_3378_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3560_io_b = FullAdder_3379_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3560_io_ci = FullAdder_3380_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3561_io_a = FullAdder_3381_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3561_io_b = FullAdder_3382_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3561_io_ci = FullAdder_3383_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3562_io_a = FullAdder_3096_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3562_io_b = FullAdder_3381_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3562_io_ci = FullAdder_3382_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3563_io_a = FullAdder_3383_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3563_io_b = FullAdder_3384_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3563_io_ci = FullAdder_3385_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3564_io_a = FullAdder_3384_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3564_io_b = FullAdder_3385_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3564_io_ci = FullAdder_3386_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3565_io_a = FullAdder_3387_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3565_io_b = FullAdder_3388_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3565_io_ci = HalfAdder_132_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3566_io_a = FullAdder_3387_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3566_io_b = FullAdder_3388_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3566_io_ci = HalfAdder_132_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_168_io_a = FullAdder_3389_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_168_io_b = FullAdder_3390_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3567_io_a = FullAdder_3106_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3567_io_b = FullAdder_3107_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3567_io_ci = FullAdder_3389_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3568_io_a = FullAdder_3390_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3568_io_b = FullAdder_3391_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3568_io_ci = FullAdder_3392_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3569_io_a = FullAdder_3391_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3569_io_b = FullAdder_3392_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3569_io_ci = FullAdder_3393_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3570_io_a = FullAdder_3394_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3570_io_b = FullAdder_3395_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3570_io_ci = FullAdder_3396_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3571_io_a = FullAdder_3394_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3571_io_b = FullAdder_3395_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3571_io_ci = FullAdder_3396_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3572_io_a = FullAdder_3118_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3572_io_b = HalfAdder_107_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3572_io_ci = FullAdder_3397_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3573_io_a = FullAdder_3398_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3573_io_b = FullAdder_3399_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3573_io_ci = FullAdder_3400_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3574_io_a = FullAdder_3121_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3574_io_b = FullAdder_3399_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3574_io_ci = FullAdder_3400_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3575_io_a = FullAdder_3401_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3575_io_b = FullAdder_3402_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3575_io_ci = HalfAdder_133_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3576_io_a = FullAdder_3401_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3576_io_b = FullAdder_3402_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3576_io_ci = HalfAdder_133_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_169_io_a = FullAdder_3403_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_169_io_b = FullAdder_3404_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3577_io_a = FullAdder_3128_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3577_io_b = FullAdder_3403_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3577_io_ci = FullAdder_3404_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3578_io_a = FullAdder_3131_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3578_io_b = FullAdder_3405_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3578_io_ci = FullAdder_3406_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_170_io_a = FullAdder_3407_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_170_io_b = FullAdder_3408_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3579_io_a = FullAdder_3407_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3579_io_b = FullAdder_3408_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3579_io_ci = FullAdder_3409_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3580_io_a = FullAdder_3136_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3580_io_b = FullAdder_3137_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3580_io_ci = FullAdder_3409_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3581_io_a = FullAdder_3410_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3581_io_b = FullAdder_3411_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3581_io_ci = FullAdder_3412_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3582_io_a = FullAdder_3411_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3582_io_b = FullAdder_3412_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3582_io_ci = FullAdder_3413_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3583_io_a = FullAdder_3413_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3583_io_b = FullAdder_3414_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3583_io_ci = FullAdder_3415_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3584_io_a = FullAdder_3415_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3584_io_b = FullAdder_3416_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3584_io_ci = FullAdder_3417_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3585_io_a = FullAdder_3147_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3585_io_b = FullAdder_3148_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3585_io_ci = FullAdder_3417_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3586_io_a = FullAdder_3418_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3586_io_b = FullAdder_3419_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3586_io_ci = FullAdder_3420_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3587_io_a = FullAdder_3152_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3587_io_b = FullAdder_3153_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3587_io_ci = FullAdder_3420_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3588_io_a = FullAdder_3421_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3588_io_b = FullAdder_3422_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3588_io_ci = FullAdder_3423_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3589_io_a = FullAdder_3423_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3589_io_b = HalfAdder_134_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3589_io_ci = FullAdder_3424_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3590_io_a = FullAdder_3424_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3590_io_b = HalfAdder_135_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3590_io_ci = FullAdder_3425_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3591_io_a = FullAdder_3425_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3591_io_b = HalfAdder_136_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3591_io_ci = FullAdder_3426_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3592_io_a = FullAdder_3163_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3592_io_b = FullAdder_3426_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3592_io_ci = FullAdder_3427_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_171_io_a = FullAdder_3427_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_171_io_b = FullAdder_3428_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3593_io_a = FullAdder_3165_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3593_io_b = FullAdder_3166_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3593_io_ci = FullAdder_3428_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3594_io_a = FullAdder_3167_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3594_io_b = HalfAdder_108_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3594_io_ci = FullAdder_3429_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_172_io_a = FullAdder_3430_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_172_io_b = FullAdder_3431_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3595_io_a = FullAdder_3169_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3595_io_b = HalfAdder_109_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3595_io_ci = FullAdder_3431_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3596_io_a = FullAdder_3170_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3596_io_b = FullAdder_3171_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3596_io_ci = FullAdder_3433_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3597_io_a = FullAdder_3172_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3597_io_b = FullAdder_3433_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3597_io_ci = FullAdder_3434_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3598_io_a = HalfAdder_110_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3598_io_b = HalfAdder_111_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3598_io_ci = FullAdder_3434_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_173_io_a = HalfAdder_137_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_173_io_b = HalfAdder_138_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3599_io_a = FullAdder_3173_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3599_io_b = FullAdder_3174_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3599_io_ci = HalfAdder_139_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_174_io_a = HalfAdder_142_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_174_io_b = HalfAdder_143_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_175_io_a = HalfAdder_115_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_175_io_b = HalfAdder_144_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3600_io_a = FullAdder_3176_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3600_io_b = HalfAdder_116_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3600_io_ci = HalfAdder_145_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_176_io_a = HalfAdder_117_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_176_io_b = HalfAdder_145_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_177_io_a = HalfAdder_147_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_177_io_b = HalfAdder_148_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_178_io_a = HalfAdder_119_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_178_io_b = HalfAdder_148_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3601_io_a = HalfAdder_119_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3601_io_b = FullAdder_3178_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3601_io_ci = HalfAdder_149_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3602_io_a = FullAdder_3180_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3602_io_b = FullAdder_3181_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3602_io_ci = HalfAdder_150_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3603_io_a = FullAdder_3185_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3603_io_b = FullAdder_3438_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3603_io_ci = FullAdder_3439_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3604_io_a = FullAdder_3186_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3604_io_b = FullAdder_3439_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3604_io_ci = FullAdder_3440_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_179_io_a = FullAdder_3440_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_179_io_b = FullAdder_3441_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3605_io_a = HalfAdder_120_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3605_io_b = FullAdder_3441_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3605_io_ci = FullAdder_3442_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3606_io_a = HalfAdder_121_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3606_io_b = FullAdder_3442_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3606_io_ci = FullAdder_3443_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3607_io_a = FullAdder_3191_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3607_io_b = FullAdder_3443_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3607_io_ci = FullAdder_3444_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_180_io_a = FullAdder_3444_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_180_io_b = FullAdder_3445_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3608_io_a = FullAdder_3193_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3608_io_b = FullAdder_3194_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3608_io_ci = FullAdder_3445_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3609_io_a = FullAdder_3196_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3609_io_b = FullAdder_3446_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3609_io_ci = FullAdder_3447_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3610_io_a = FullAdder_3198_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3610_io_b = FullAdder_3447_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3610_io_ci = FullAdder_3448_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3611_io_a = FullAdder_3200_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3611_io_b = FullAdder_3448_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3611_io_ci = FullAdder_3449_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3612_io_a = FullAdder_3202_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3612_io_b = FullAdder_3449_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3612_io_ci = HalfAdder_151_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_181_io_a = HalfAdder_151_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_181_io_b = HalfAdder_152_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3613_io_a = FullAdder_3205_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3613_io_b = FullAdder_3206_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3613_io_ci = FullAdder_3450_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3614_io_a = FullAdder_3207_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3614_io_b = FullAdder_3208_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3614_io_ci = FullAdder_3451_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3615_io_a = FullAdder_3452_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3615_io_b = FullAdder_3453_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3615_io_ci = FullAdder_3454_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3616_io_a = FullAdder_3454_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3616_io_b = HalfAdder_153_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3616_io_ci = FullAdder_3455_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3617_io_a = HalfAdder_122_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3617_io_b = FullAdder_3455_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3617_io_ci = FullAdder_3456_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3618_io_a = FullAdder_3457_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3618_io_b = FullAdder_3458_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3618_io_ci = FullAdder_3459_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_182_io_a = HalfAdder_124_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_182_io_b = FullAdder_3459_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_183_io_a = HalfAdder_154_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_183_io_b = FullAdder_3460_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3619_io_a = FullAdder_3460_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3619_io_b = FullAdder_3461_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3619_io_ci = FullAdder_3462_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3620_io_a = FullAdder_3222_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3620_io_b = FullAdder_3223_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3620_io_ci = FullAdder_3462_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3621_io_a = HalfAdder_125_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3621_io_b = FullAdder_3463_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3621_io_ci = FullAdder_3464_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3622_io_a = FullAdder_3465_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3622_io_b = FullAdder_3466_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3622_io_ci = HalfAdder_155_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_184_io_a = HalfAdder_156_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_184_io_b = HalfAdder_157_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_185_io_a = HalfAdder_155_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_185_io_b = HalfAdder_156_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_186_io_a = HalfAdder_157_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_186_io_b = FullAdder_3467_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3623_io_a = FullAdder_3467_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3623_io_b = FullAdder_3468_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3623_io_ci = FullAdder_3469_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3624_io_a = FullAdder_3236_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3624_io_b = FullAdder_3469_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3624_io_ci = FullAdder_3470_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_187_io_a = FullAdder_3471_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_187_io_b = FullAdder_3472_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3625_io_a = FullAdder_3239_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3625_io_b = FullAdder_3471_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3625_io_ci = FullAdder_3472_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3626_io_a = FullAdder_3473_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3626_io_b = FullAdder_3474_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3626_io_ci = FullAdder_3475_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_188_io_a = FullAdder_3245_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_188_io_b = FullAdder_3475_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_189_io_a = FullAdder_3476_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_189_io_b = FullAdder_3477_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3627_io_a = FullAdder_3248_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3627_io_b = FullAdder_3477_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3627_io_ci = FullAdder_3478_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3628_io_a = FullAdder_3251_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3628_io_b = FullAdder_3479_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3628_io_ci = FullAdder_3480_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3629_io_a = FullAdder_3253_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3629_io_b = FullAdder_3254_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3629_io_ci = FullAdder_3481_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3630_io_a = FullAdder_3482_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3630_io_b = FullAdder_3483_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3630_io_ci = FullAdder_3484_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3631_io_a = FullAdder_3483_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3631_io_b = FullAdder_3484_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3631_io_ci = HalfAdder_158_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_190_io_a = FullAdder_3485_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_190_io_b = FullAdder_3486_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3632_io_a = FullAdder_3261_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3632_io_b = HalfAdder_127_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3632_io_ci = FullAdder_3485_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3633_io_a = FullAdder_3486_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3633_io_b = FullAdder_3487_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3633_io_ci = FullAdder_3488_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3634_io_a = FullAdder_3264_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3634_io_b = HalfAdder_128_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3634_io_ci = FullAdder_3487_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3635_io_a = FullAdder_3488_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3635_io_b = FullAdder_3489_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3635_io_ci = FullAdder_3490_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3636_io_a = FullAdder_3489_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3636_io_b = FullAdder_3490_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3636_io_ci = HalfAdder_159_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3637_io_a = FullAdder_3270_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3637_io_b = FullAdder_3271_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3637_io_ci = FullAdder_3491_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3638_io_a = FullAdder_3492_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3638_io_b = FullAdder_3493_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3638_io_ci = FullAdder_3494_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3639_io_a = FullAdder_3493_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3639_io_b = FullAdder_3494_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3639_io_ci = HalfAdder_160_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3640_io_a = FullAdder_3495_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3640_io_b = FullAdder_3496_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3640_io_ci = HalfAdder_161_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3641_io_a = FullAdder_3495_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3641_io_b = FullAdder_3496_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3641_io_ci = HalfAdder_161_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_191_io_a = FullAdder_3497_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_191_io_b = FullAdder_3498_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3642_io_a = FullAdder_3282_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3642_io_b = FullAdder_3283_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3642_io_ci = FullAdder_3497_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3643_io_a = FullAdder_3498_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3643_io_b = FullAdder_3499_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3643_io_ci = FullAdder_3500_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3644_io_a = FullAdder_3286_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3644_io_b = FullAdder_3287_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3644_io_ci = FullAdder_3499_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3645_io_a = FullAdder_3500_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3645_io_b = FullAdder_3501_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3645_io_ci = FullAdder_3502_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3646_io_a = FullAdder_3290_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3646_io_b = FullAdder_3291_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3646_io_ci = FullAdder_3501_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3647_io_a = FullAdder_3502_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3647_io_b = FullAdder_3503_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3647_io_ci = FullAdder_3504_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3648_io_a = FullAdder_3503_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3648_io_b = FullAdder_3504_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3648_io_ci = HalfAdder_162_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3649_io_a = FullAdder_3505_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3649_io_b = FullAdder_3506_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3649_io_ci = HalfAdder_163_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3650_io_a = FullAdder_3505_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3650_io_b = FullAdder_3506_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3650_io_ci = HalfAdder_163_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3651_io_a = FullAdder_3507_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3651_io_b = HalfAdder_164_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3651_io_ci = HalfAdder_165_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_192_io_a = FullAdder_3507_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_192_io_b = HalfAdder_164_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_193_io_a = HalfAdder_165_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_193_io_b = HalfAdder_166_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_194_io_a = FullAdder_3508_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_194_io_b = FullAdder_3509_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3652_io_a = HalfAdder_130_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3652_io_b = FullAdder_3508_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3652_io_ci = FullAdder_3509_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3653_io_a = FullAdder_3510_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3653_io_b = FullAdder_3511_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3653_io_ci = FullAdder_3512_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3654_io_a = FullAdder_3511_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3654_io_b = FullAdder_3512_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3654_io_ci = FullAdder_3513_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3655_io_a = FullAdder_3514_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3655_io_b = FullAdder_3515_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3655_io_ci = FullAdder_3516_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3656_io_a = FullAdder_3514_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3656_io_b = FullAdder_3515_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3656_io_ci = FullAdder_3516_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3657_io_a = FullAdder_3517_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3657_io_b = FullAdder_3518_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3657_io_ci = FullAdder_3519_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3658_io_a = FullAdder_3517_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3658_io_b = FullAdder_3518_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3658_io_ci = FullAdder_3519_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3659_io_a = FullAdder_3520_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3659_io_b = FullAdder_3521_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3659_io_ci = FullAdder_3522_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3660_io_a = FullAdder_3520_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3660_io_b = FullAdder_3521_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3660_io_ci = FullAdder_3522_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_195_io_a = FullAdder_3523_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_195_io_b = FullAdder_3524_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3661_io_a = FullAdder_3326_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3661_io_b = FullAdder_3327_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3661_io_ci = FullAdder_3523_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3662_io_a = FullAdder_3524_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3662_io_b = FullAdder_3525_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3662_io_ci = FullAdder_3526_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3663_io_a = FullAdder_3329_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3663_io_b = FullAdder_3330_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3663_io_ci = FullAdder_3525_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3664_io_a = FullAdder_3526_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3664_io_b = FullAdder_3527_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3664_io_ci = FullAdder_3528_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3665_io_a = FullAdder_3527_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3665_io_b = FullAdder_3528_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3665_io_ci = FullAdder_3529_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3666_io_a = FullAdder_3530_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3666_io_b = FullAdder_3531_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3666_io_ci = FullAdder_3532_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3667_io_a = FullAdder_3530_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3667_io_b = FullAdder_3531_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3667_io_ci = FullAdder_3532_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3668_io_a = FullAdder_3533_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3668_io_b = FullAdder_3534_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3668_io_ci = HalfAdder_167_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3669_io_a = FullAdder_3533_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3669_io_b = FullAdder_3534_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3669_io_ci = HalfAdder_167_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3670_io_a = FullAdder_3345_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3670_io_b = FullAdder_3535_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3670_io_ci = FullAdder_3536_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3671_io_a = FullAdder_3537_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3671_io_b = FullAdder_3538_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3671_io_ci = FullAdder_3539_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3672_io_a = FullAdder_3537_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3672_io_b = FullAdder_3538_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3672_io_ci = FullAdder_3539_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3673_io_a = FullAdder_3351_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3673_io_b = FullAdder_3352_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3673_io_ci = FullAdder_3540_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3674_io_a = FullAdder_3541_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3674_io_b = FullAdder_3542_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3674_io_ci = FullAdder_3543_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3675_io_a = FullAdder_3355_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3675_io_b = FullAdder_3356_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3675_io_ci = FullAdder_3542_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3676_io_a = FullAdder_3543_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3676_io_b = FullAdder_3544_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3676_io_ci = FullAdder_3545_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3677_io_a = FullAdder_3359_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3677_io_b = FullAdder_3544_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3677_io_ci = FullAdder_3545_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3678_io_a = FullAdder_3362_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3678_io_b = FullAdder_3546_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3678_io_ci = FullAdder_3547_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_196_io_a = FullAdder_3548_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_196_io_b = FullAdder_3549_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3679_io_a = FullAdder_3365_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3679_io_b = FullAdder_3548_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3679_io_ci = FullAdder_3549_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3680_io_a = FullAdder_3367_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3680_io_b = FullAdder_3368_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3680_io_ci = FullAdder_3550_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3681_io_a = FullAdder_3551_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3681_io_b = FullAdder_3552_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3681_io_ci = FullAdder_3553_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3682_io_a = FullAdder_3371_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3682_io_b = FullAdder_3552_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3682_io_ci = FullAdder_3553_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_197_io_a = FullAdder_3554_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_197_io_b = FullAdder_3555_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3683_io_a = FullAdder_3554_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3683_io_b = FullAdder_3555_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3683_io_ci = FullAdder_3556_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3684_io_a = FullAdder_3377_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3684_io_b = FullAdder_3556_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3684_io_ci = FullAdder_3557_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3685_io_a = FullAdder_3380_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3685_io_b = FullAdder_3558_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3685_io_ci = FullAdder_3559_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3686_io_a = FullAdder_3560_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3686_io_b = FullAdder_3561_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3686_io_ci = FullAdder_3562_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3687_io_a = FullAdder_3386_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3687_io_b = FullAdder_3562_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3687_io_ci = FullAdder_3563_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3688_io_a = FullAdder_3564_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3688_io_b = FullAdder_3565_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3688_io_ci = FullAdder_3566_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3689_io_a = FullAdder_3566_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3689_io_b = HalfAdder_168_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3689_io_ci = FullAdder_3567_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3690_io_a = FullAdder_3393_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3690_io_b = FullAdder_3567_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3690_io_ci = FullAdder_3568_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3691_io_a = FullAdder_3569_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3691_io_b = FullAdder_3570_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3691_io_ci = FullAdder_3571_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3692_io_a = FullAdder_3397_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3692_io_b = FullAdder_3398_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3692_io_ci = FullAdder_3571_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3693_io_a = FullAdder_3572_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3693_io_b = FullAdder_3573_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3693_io_ci = FullAdder_3574_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3694_io_a = FullAdder_3574_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3694_io_b = FullAdder_3575_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3694_io_ci = FullAdder_3576_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3695_io_a = FullAdder_3576_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3695_io_b = HalfAdder_169_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3695_io_ci = FullAdder_3577_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3696_io_a = FullAdder_3405_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3696_io_b = FullAdder_3406_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3696_io_ci = FullAdder_3577_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3697_io_a = FullAdder_3578_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3697_io_b = HalfAdder_170_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3697_io_ci = FullAdder_3579_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3698_io_a = FullAdder_3410_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3698_io_b = FullAdder_3579_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3698_io_ci = FullAdder_3580_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3699_io_a = FullAdder_3580_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3699_io_b = FullAdder_3581_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3699_io_ci = FullAdder_3582_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3700_io_a = FullAdder_3414_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3700_io_b = FullAdder_3582_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3700_io_ci = FullAdder_3583_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3701_io_a = FullAdder_3416_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3701_io_b = FullAdder_3583_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3701_io_ci = FullAdder_3584_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3702_io_a = FullAdder_3418_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3702_io_b = FullAdder_3419_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3702_io_ci = FullAdder_3585_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_198_io_a = FullAdder_3586_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_198_io_b = FullAdder_3587_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3703_io_a = FullAdder_3421_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3703_io_b = FullAdder_3422_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3703_io_ci = FullAdder_3587_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3704_io_a = HalfAdder_134_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3704_io_b = FullAdder_3588_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3704_io_ci = FullAdder_3589_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3705_io_a = HalfAdder_135_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3705_io_b = FullAdder_3589_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3705_io_ci = FullAdder_3590_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3706_io_a = HalfAdder_136_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3706_io_b = FullAdder_3590_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3706_io_ci = FullAdder_3591_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_199_io_a = FullAdder_3591_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_199_io_b = FullAdder_3592_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_200_io_a = FullAdder_3592_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_200_io_b = HalfAdder_171_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3707_io_a = FullAdder_3429_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3707_io_b = FullAdder_3593_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3707_io_ci = FullAdder_3594_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3708_io_a = FullAdder_3430_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3708_io_b = FullAdder_3594_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3708_io_ci = HalfAdder_172_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3709_io_a = HalfAdder_137_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3709_io_b = HalfAdder_138_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3709_io_ci = FullAdder_3598_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_201_io_a = HalfAdder_173_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_201_io_b = FullAdder_3599_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3710_io_a = HalfAdder_141_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3710_io_b = HalfAdder_142_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3710_io_ci = HalfAdder_174_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_202_io_a = HalfAdder_144_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_202_io_b = FullAdder_3600_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_203_io_a = HalfAdder_146_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_203_io_b = HalfAdder_176_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3711_io_a = HalfAdder_146_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3711_io_b = HalfAdder_147_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3711_io_ci = HalfAdder_177_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_204_io_a = HalfAdder_177_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_204_io_b = HalfAdder_178_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_205_io_a = HalfAdder_178_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_205_io_b = FullAdder_3601_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3712_io_a = FullAdder_3437_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3712_io_b = FullAdder_3438_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3712_io_ci = FullAdder_3603_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_206_io_a = HalfAdder_179_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_206_io_b = FullAdder_3605_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_207_io_a = FullAdder_3606_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_207_io_b = FullAdder_3607_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_208_io_a = HalfAdder_180_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_208_io_b = FullAdder_3608_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3713_io_a = FullAdder_3446_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3713_io_b = FullAdder_3608_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3713_io_ci = FullAdder_3609_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_209_io_a = FullAdder_3609_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_209_io_b = FullAdder_3610_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3714_io_a = HalfAdder_152_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3714_io_b = FullAdder_3612_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3714_io_ci = HalfAdder_181_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_210_io_a = FullAdder_3450_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_210_io_b = HalfAdder_181_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3715_io_a = FullAdder_3451_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3715_io_b = FullAdder_3613_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3715_io_ci = FullAdder_3614_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3716_io_a = FullAdder_3452_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3716_io_b = FullAdder_3453_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3716_io_ci = FullAdder_3614_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3717_io_a = HalfAdder_153_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3717_io_b = FullAdder_3615_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3717_io_ci = FullAdder_3616_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3718_io_a = FullAdder_3456_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3718_io_b = FullAdder_3616_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3718_io_ci = FullAdder_3617_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3719_io_a = FullAdder_3457_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3719_io_b = FullAdder_3458_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3719_io_ci = FullAdder_3617_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3720_io_a = HalfAdder_154_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3720_io_b = FullAdder_3618_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3720_io_ci = HalfAdder_182_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_211_io_a = FullAdder_3461_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_211_io_b = HalfAdder_182_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_212_io_a = HalfAdder_183_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_212_io_b = FullAdder_3619_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_213_io_a = FullAdder_3619_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_213_io_b = FullAdder_3620_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3721_io_a = FullAdder_3463_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3721_io_b = FullAdder_3464_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3721_io_ci = FullAdder_3620_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3722_io_a = FullAdder_3465_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3722_io_b = FullAdder_3466_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3722_io_ci = FullAdder_3621_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3723_io_a = FullAdder_3622_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3723_io_b = HalfAdder_184_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3723_io_ci = HalfAdder_185_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_214_io_a = FullAdder_3468_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_214_io_b = HalfAdder_185_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_215_io_a = HalfAdder_186_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_215_io_b = FullAdder_3623_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3724_io_a = FullAdder_3470_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3724_io_b = FullAdder_3623_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3724_io_ci = FullAdder_3624_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3725_io_a = FullAdder_3624_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3725_io_b = HalfAdder_187_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3725_io_ci = FullAdder_3625_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3726_io_a = FullAdder_3473_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3726_io_b = FullAdder_3474_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3726_io_ci = FullAdder_3625_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3727_io_a = FullAdder_3476_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3727_io_b = FullAdder_3626_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3727_io_ci = HalfAdder_188_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_216_io_a = FullAdder_3478_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_216_io_b = HalfAdder_188_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_217_io_a = HalfAdder_189_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_217_io_b = FullAdder_3627_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3728_io_a = FullAdder_3479_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3728_io_b = FullAdder_3480_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3728_io_ci = FullAdder_3627_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3729_io_a = FullAdder_3481_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3729_io_b = FullAdder_3482_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3729_io_ci = FullAdder_3628_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3730_io_a = HalfAdder_158_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3730_io_b = FullAdder_3629_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3730_io_ci = FullAdder_3630_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3731_io_a = FullAdder_3631_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3731_io_b = HalfAdder_190_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3731_io_ci = FullAdder_3632_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3732_io_a = FullAdder_3632_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3732_io_b = FullAdder_3633_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3732_io_ci = FullAdder_3634_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3733_io_a = HalfAdder_159_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3733_io_b = FullAdder_3634_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3733_io_ci = FullAdder_3635_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3734_io_a = FullAdder_3491_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3734_io_b = FullAdder_3492_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3734_io_ci = FullAdder_3636_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3735_io_a = HalfAdder_160_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3735_io_b = FullAdder_3637_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3735_io_ci = FullAdder_3638_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3736_io_a = FullAdder_3639_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3736_io_b = FullAdder_3640_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3736_io_ci = FullAdder_3641_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3737_io_a = FullAdder_3641_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3737_io_b = HalfAdder_191_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3737_io_ci = FullAdder_3642_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3738_io_a = FullAdder_3642_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3738_io_b = FullAdder_3643_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3738_io_ci = FullAdder_3644_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3739_io_a = FullAdder_3644_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3739_io_b = FullAdder_3645_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3739_io_ci = FullAdder_3646_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3740_io_a = HalfAdder_162_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3740_io_b = FullAdder_3646_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3740_io_ci = FullAdder_3647_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3741_io_a = FullAdder_3648_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3741_io_b = FullAdder_3649_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3741_io_ci = FullAdder_3650_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3742_io_a = HalfAdder_166_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3742_io_b = FullAdder_3650_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3742_io_ci = FullAdder_3651_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3743_io_a = HalfAdder_192_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3743_io_b = HalfAdder_193_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3743_io_ci = HalfAdder_194_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_218_io_a = FullAdder_3510_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_218_io_b = HalfAdder_192_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_219_io_a = HalfAdder_193_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_219_io_b = HalfAdder_194_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_220_io_a = FullAdder_3652_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_220_io_b = FullAdder_3653_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3744_io_a = FullAdder_3513_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3744_io_b = FullAdder_3652_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3744_io_ci = FullAdder_3653_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_221_io_a = FullAdder_3654_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_221_io_b = FullAdder_3655_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3745_io_a = FullAdder_3654_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3745_io_b = FullAdder_3655_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3745_io_ci = FullAdder_3656_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3746_io_a = FullAdder_3656_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3746_io_b = FullAdder_3657_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3746_io_ci = FullAdder_3658_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3747_io_a = FullAdder_3658_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3747_io_b = FullAdder_3659_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3747_io_ci = FullAdder_3660_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3748_io_a = FullAdder_3660_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3748_io_b = HalfAdder_195_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3748_io_ci = FullAdder_3661_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3749_io_a = FullAdder_3661_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3749_io_b = FullAdder_3662_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3749_io_ci = FullAdder_3663_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3750_io_a = FullAdder_3529_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3750_io_b = FullAdder_3663_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3750_io_ci = FullAdder_3664_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3751_io_a = FullAdder_3665_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3751_io_b = FullAdder_3666_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3751_io_ci = FullAdder_3667_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3752_io_a = FullAdder_3667_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3752_io_b = FullAdder_3668_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3752_io_ci = FullAdder_3669_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3753_io_a = FullAdder_3535_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3753_io_b = FullAdder_3536_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3753_io_ci = FullAdder_3669_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3754_io_a = FullAdder_3670_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3754_io_b = FullAdder_3671_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3754_io_ci = FullAdder_3672_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3755_io_a = FullAdder_3540_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3755_io_b = FullAdder_3541_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3755_io_ci = FullAdder_3672_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3756_io_a = FullAdder_3673_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3756_io_b = FullAdder_3674_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3756_io_ci = FullAdder_3675_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3757_io_a = FullAdder_3675_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3757_io_b = FullAdder_3676_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3757_io_ci = FullAdder_3677_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3758_io_a = FullAdder_3546_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3758_io_b = FullAdder_3547_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3758_io_ci = FullAdder_3677_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3759_io_a = FullAdder_3678_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3759_io_b = HalfAdder_196_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3759_io_ci = FullAdder_3679_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3760_io_a = FullAdder_3550_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3760_io_b = FullAdder_3551_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3760_io_ci = FullAdder_3679_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3761_io_a = FullAdder_3680_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3761_io_b = FullAdder_3681_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3761_io_ci = FullAdder_3682_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3762_io_a = FullAdder_3682_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3762_io_b = HalfAdder_197_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3762_io_ci = FullAdder_3683_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3763_io_a = FullAdder_3557_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3763_io_b = FullAdder_3683_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3763_io_ci = FullAdder_3684_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3764_io_a = FullAdder_3558_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3764_io_b = FullAdder_3559_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3764_io_ci = FullAdder_3684_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3765_io_a = FullAdder_3560_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3765_io_b = FullAdder_3561_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3765_io_ci = FullAdder_3685_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3766_io_a = FullAdder_3563_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3766_io_b = FullAdder_3686_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3766_io_ci = FullAdder_3687_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3767_io_a = FullAdder_3564_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3767_io_b = FullAdder_3565_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3767_io_ci = FullAdder_3687_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3768_io_a = HalfAdder_168_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3768_io_b = FullAdder_3688_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3768_io_ci = FullAdder_3689_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_222_io_a = FullAdder_3568_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_222_io_b = FullAdder_3689_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3769_io_a = FullAdder_3569_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3769_io_b = FullAdder_3570_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3769_io_ci = FullAdder_3690_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3770_io_a = FullAdder_3572_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3770_io_b = FullAdder_3573_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3770_io_ci = FullAdder_3692_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3771_io_a = FullAdder_3575_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3771_io_b = FullAdder_3693_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3771_io_ci = FullAdder_3694_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3772_io_a = HalfAdder_169_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3772_io_b = FullAdder_3694_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3772_io_ci = FullAdder_3695_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_223_io_a = FullAdder_3695_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_223_io_b = FullAdder_3696_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3773_io_a = FullAdder_3578_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3773_io_b = HalfAdder_170_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3773_io_ci = FullAdder_3696_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_224_io_a = FullAdder_3697_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_224_io_b = FullAdder_3698_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3774_io_a = FullAdder_3581_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3774_io_b = FullAdder_3698_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3774_io_ci = FullAdder_3699_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_225_io_a = FullAdder_3700_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_225_io_b = FullAdder_3701_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3775_io_a = FullAdder_3584_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3775_io_b = FullAdder_3585_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3775_io_ci = FullAdder_3702_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3776_io_a = FullAdder_3586_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3776_io_b = FullAdder_3702_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3776_io_ci = HalfAdder_198_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_226_io_a = HalfAdder_198_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_226_io_b = FullAdder_3703_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3777_io_a = FullAdder_3588_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3777_io_b = FullAdder_3703_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3777_io_ci = FullAdder_3704_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3778_io_a = HalfAdder_171_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3778_io_b = FullAdder_3593_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3778_io_ci = FullAdder_3707_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3779_io_a = FullAdder_3597_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3779_io_b = FullAdder_3598_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3779_io_ci = FullAdder_3709_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3780_io_a = HalfAdder_173_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3780_io_b = FullAdder_3709_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3780_io_ci = HalfAdder_201_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3781_io_a = HalfAdder_140_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3781_io_b = HalfAdder_141_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3781_io_ci = FullAdder_3710_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_227_io_a = HalfAdder_175_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_227_io_b = HalfAdder_202_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3782_io_a = FullAdder_3600_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3782_io_b = HalfAdder_176_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3782_io_ci = HalfAdder_203_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_228_io_a = HalfAdder_203_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_228_io_b = FullAdder_3711_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_229_io_a = HalfAdder_204_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_229_io_b = HalfAdder_205_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3783_io_a = FullAdder_3436_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3783_io_b = FullAdder_3437_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3783_io_ci = FullAdder_3712_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3784_io_a = FullAdder_3604_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3784_io_b = HalfAdder_179_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3784_io_ci = HalfAdder_206_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3785_io_a = FullAdder_3605_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3785_io_b = FullAdder_3606_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3785_io_ci = HalfAdder_207_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3786_io_a = FullAdder_3607_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3786_io_b = HalfAdder_180_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3786_io_ci = HalfAdder_208_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_230_io_a = HalfAdder_208_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_230_io_b = FullAdder_3713_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3787_io_a = FullAdder_3611_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3787_io_b = FullAdder_3612_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3787_io_ci = FullAdder_3714_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_231_io_a = FullAdder_3613_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_231_io_b = HalfAdder_210_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3788_io_a = FullAdder_3615_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3788_io_b = FullAdder_3716_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3788_io_ci = FullAdder_3717_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3789_io_a = FullAdder_3618_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3789_io_b = FullAdder_3719_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3789_io_ci = FullAdder_3720_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3790_io_a = HalfAdder_183_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3790_io_b = FullAdder_3720_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3790_io_ci = HalfAdder_211_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_232_io_a = HalfAdder_211_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_232_io_b = HalfAdder_212_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3791_io_a = FullAdder_3621_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3791_io_b = FullAdder_3721_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3791_io_ci = FullAdder_3722_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3792_io_a = FullAdder_3622_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3792_io_b = HalfAdder_184_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3792_io_ci = FullAdder_3722_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3793_io_a = HalfAdder_186_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3793_io_b = FullAdder_3723_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3793_io_ci = HalfAdder_214_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_233_io_a = HalfAdder_214_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_233_io_b = HalfAdder_215_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3794_io_a = HalfAdder_187_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3794_io_b = FullAdder_3724_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3794_io_ci = FullAdder_3725_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_234_io_a = FullAdder_3725_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_234_io_b = FullAdder_3726_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3795_io_a = FullAdder_3626_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3795_io_b = FullAdder_3726_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3795_io_ci = FullAdder_3727_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3796_io_a = HalfAdder_189_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3796_io_b = FullAdder_3727_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3796_io_ci = HalfAdder_216_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_235_io_a = HalfAdder_216_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_235_io_b = HalfAdder_217_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3797_io_a = FullAdder_3628_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3797_io_b = FullAdder_3728_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3797_io_ci = FullAdder_3729_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3798_io_a = FullAdder_3629_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3798_io_b = FullAdder_3630_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3798_io_ci = FullAdder_3729_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3799_io_a = FullAdder_3631_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3799_io_b = HalfAdder_190_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3799_io_ci = FullAdder_3730_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3800_io_a = FullAdder_3633_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3800_io_b = FullAdder_3731_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3800_io_ci = FullAdder_3732_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3801_io_a = FullAdder_3635_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3801_io_b = FullAdder_3732_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3801_io_ci = FullAdder_3733_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3802_io_a = FullAdder_3636_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3802_io_b = FullAdder_3733_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3802_io_ci = FullAdder_3734_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3803_io_a = FullAdder_3637_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3803_io_b = FullAdder_3638_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3803_io_ci = FullAdder_3734_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3804_io_a = FullAdder_3639_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3804_io_b = FullAdder_3640_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3804_io_ci = FullAdder_3735_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3805_io_a = HalfAdder_191_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3805_io_b = FullAdder_3736_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3805_io_ci = FullAdder_3737_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3806_io_a = FullAdder_3643_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3806_io_b = FullAdder_3737_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3806_io_ci = FullAdder_3738_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3807_io_a = FullAdder_3645_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3807_io_b = FullAdder_3738_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3807_io_ci = FullAdder_3739_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3808_io_a = FullAdder_3647_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3808_io_b = FullAdder_3739_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3808_io_ci = FullAdder_3740_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3809_io_a = FullAdder_3648_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3809_io_b = FullAdder_3649_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3809_io_ci = FullAdder_3740_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3810_io_a = FullAdder_3651_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3810_io_b = FullAdder_3741_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3810_io_ci = FullAdder_3742_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3811_io_a = FullAdder_3742_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3811_io_b = FullAdder_3743_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3811_io_ci = HalfAdder_218_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_236_io_a = HalfAdder_219_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_236_io_b = HalfAdder_220_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_237_io_a = HalfAdder_218_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_237_io_b = HalfAdder_219_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_238_io_a = HalfAdder_220_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_238_io_b = FullAdder_3744_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3812_io_a = FullAdder_3744_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3812_io_b = HalfAdder_221_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3812_io_ci = FullAdder_3745_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3813_io_a = FullAdder_3657_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3813_io_b = FullAdder_3745_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3813_io_ci = FullAdder_3746_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3814_io_a = FullAdder_3659_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3814_io_b = FullAdder_3746_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3814_io_ci = FullAdder_3747_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3815_io_a = HalfAdder_195_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3815_io_b = FullAdder_3747_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3815_io_ci = FullAdder_3748_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_239_io_a = FullAdder_3662_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_239_io_b = FullAdder_3748_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3816_io_a = FullAdder_3664_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3816_io_b = FullAdder_3749_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3816_io_ci = FullAdder_3750_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3817_io_a = FullAdder_3665_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3817_io_b = FullAdder_3666_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3817_io_ci = FullAdder_3750_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3818_io_a = FullAdder_3668_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3818_io_b = FullAdder_3751_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3818_io_ci = FullAdder_3752_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3819_io_a = FullAdder_3670_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3819_io_b = FullAdder_3671_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3819_io_ci = FullAdder_3753_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3820_io_a = FullAdder_3673_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3820_io_b = FullAdder_3674_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3820_io_ci = FullAdder_3755_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3821_io_a = FullAdder_3676_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3821_io_b = FullAdder_3756_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3821_io_ci = FullAdder_3757_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3822_io_a = FullAdder_3678_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3822_io_b = HalfAdder_196_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3822_io_ci = FullAdder_3758_io_s; // @[wallace.scala 71:19]
  assign HalfAdder_240_io_a = FullAdder_3759_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_240_io_b = FullAdder_3760_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3823_io_a = FullAdder_3680_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3823_io_b = FullAdder_3681_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3823_io_ci = FullAdder_3760_io_s; // @[wallace.scala 71:19]
  assign FullAdder_3824_io_a = HalfAdder_197_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3824_io_b = FullAdder_3761_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3824_io_ci = FullAdder_3762_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_241_io_a = FullAdder_3763_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_241_io_b = FullAdder_3764_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3825_io_a = FullAdder_3685_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3825_io_b = FullAdder_3764_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3825_io_ci = FullAdder_3765_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3826_io_a = FullAdder_3686_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3826_io_b = FullAdder_3765_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3826_io_ci = FullAdder_3766_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3827_io_a = FullAdder_3688_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3827_io_b = FullAdder_3767_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3827_io_ci = FullAdder_3768_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_242_io_a = FullAdder_3690_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_242_io_b = HalfAdder_222_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3828_io_a = FullAdder_3691_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3828_io_b = FullAdder_3692_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3828_io_ci = FullAdder_3770_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3829_io_a = FullAdder_3693_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3829_io_b = FullAdder_3770_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3829_io_ci = FullAdder_3771_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_243_io_a = FullAdder_3772_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_243_io_b = HalfAdder_223_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3830_io_a = FullAdder_3697_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3830_io_b = FullAdder_3773_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3830_io_ci = HalfAdder_224_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_244_io_a = HalfAdder_224_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_244_io_b = FullAdder_3774_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3831_io_a = FullAdder_3699_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3831_io_b = FullAdder_3700_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3831_io_ci = HalfAdder_225_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_245_io_a = FullAdder_3701_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_245_io_b = FullAdder_3775_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_246_io_a = HalfAdder_226_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_246_io_b = FullAdder_3777_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_247_io_a = HalfAdder_200_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_247_io_b = FullAdder_3778_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3832_io_a = FullAdder_3596_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3832_io_b = FullAdder_3597_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3832_io_ci = FullAdder_3779_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3833_io_a = HalfAdder_139_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3833_io_b = HalfAdder_140_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3833_io_ci = FullAdder_3781_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_248_io_a = HalfAdder_202_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_248_io_b = FullAdder_3782_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3834_io_a = FullAdder_3711_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3834_io_b = HalfAdder_204_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3834_io_ci = HalfAdder_229_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3835_io_a = HalfAdder_150_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3835_io_b = FullAdder_3436_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3835_io_ci = FullAdder_3783_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3836_io_a = FullAdder_3603_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3836_io_b = FullAdder_3604_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3836_io_ci = FullAdder_3784_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3837_io_a = FullAdder_3610_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3837_io_b = FullAdder_3611_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3837_io_ci = FullAdder_3787_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3838_io_a = FullAdder_3714_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3838_io_b = HalfAdder_210_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3838_io_ci = HalfAdder_231_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_249_io_a = FullAdder_3715_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_249_io_b = HalfAdder_231_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3839_io_a = FullAdder_3715_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3839_io_b = FullAdder_3716_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3839_io_ci = FullAdder_3788_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3840_io_a = FullAdder_3718_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3840_io_b = FullAdder_3719_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3840_io_ci = FullAdder_3789_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3841_io_a = HalfAdder_212_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3841_io_b = FullAdder_3790_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3841_io_ci = HalfAdder_232_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_250_io_a = HalfAdder_213_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_250_io_b = HalfAdder_232_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3842_io_a = HalfAdder_213_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3842_io_b = FullAdder_3721_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3842_io_ci = FullAdder_3791_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3843_io_a = FullAdder_3723_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3843_io_b = FullAdder_3792_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3843_io_ci = FullAdder_3793_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3844_io_a = HalfAdder_215_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3844_io_b = FullAdder_3793_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3844_io_ci = HalfAdder_233_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_251_io_a = FullAdder_3724_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_251_io_b = HalfAdder_233_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_252_io_a = HalfAdder_234_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_252_io_b = FullAdder_3795_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3845_io_a = HalfAdder_217_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3845_io_b = FullAdder_3796_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3845_io_ci = HalfAdder_235_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_253_io_a = FullAdder_3728_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_253_io_b = HalfAdder_235_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3846_io_a = FullAdder_3730_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3846_io_b = FullAdder_3798_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3846_io_ci = FullAdder_3799_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3847_io_a = FullAdder_3731_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3847_io_b = FullAdder_3799_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3847_io_ci = FullAdder_3800_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_254_io_a = FullAdder_3800_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_254_io_b = FullAdder_3801_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3848_io_a = FullAdder_3735_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3848_io_b = FullAdder_3803_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3848_io_ci = FullAdder_3804_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3849_io_a = FullAdder_3736_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3849_io_b = FullAdder_3804_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3849_io_ci = FullAdder_3805_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_255_io_a = FullAdder_3805_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_255_io_b = FullAdder_3806_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_256_io_a = FullAdder_3806_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_256_io_b = FullAdder_3807_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3850_io_a = FullAdder_3741_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3850_io_b = FullAdder_3809_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3850_io_ci = FullAdder_3810_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3851_io_a = FullAdder_3743_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3851_io_b = FullAdder_3810_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3851_io_ci = FullAdder_3811_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3852_io_a = FullAdder_3811_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3852_io_b = HalfAdder_236_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3852_io_ci = HalfAdder_237_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_257_io_a = HalfAdder_221_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_257_io_b = HalfAdder_237_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_258_io_a = HalfAdder_238_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_258_io_b = FullAdder_3812_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_259_io_a = FullAdder_3812_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_259_io_b = FullAdder_3813_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_260_io_a = FullAdder_3814_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_260_io_b = FullAdder_3815_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_261_io_a = FullAdder_3749_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_261_io_b = HalfAdder_239_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3853_io_a = FullAdder_3751_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3853_io_b = FullAdder_3817_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3853_io_ci = FullAdder_3818_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3854_io_a = FullAdder_3752_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3854_io_b = FullAdder_3753_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3854_io_ci = FullAdder_3819_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3855_io_a = FullAdder_3754_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3855_io_b = FullAdder_3755_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3855_io_ci = FullAdder_3820_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3856_io_a = FullAdder_3756_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3856_io_b = FullAdder_3820_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3856_io_ci = FullAdder_3821_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3857_io_a = FullAdder_3757_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3857_io_b = FullAdder_3758_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3857_io_ci = FullAdder_3822_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3858_io_a = FullAdder_3759_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3858_io_b = FullAdder_3822_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3858_io_ci = HalfAdder_240_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3859_io_a = FullAdder_3761_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3859_io_b = FullAdder_3823_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3859_io_ci = FullAdder_3824_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3860_io_a = FullAdder_3762_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3860_io_b = FullAdder_3763_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3860_io_ci = HalfAdder_241_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3861_io_a = FullAdder_3766_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3861_io_b = FullAdder_3767_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3861_io_ci = FullAdder_3827_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3862_io_a = FullAdder_3768_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3862_io_b = HalfAdder_222_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3862_io_ci = HalfAdder_242_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_262_io_a = FullAdder_3769_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_262_io_b = HalfAdder_242_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3863_io_a = FullAdder_3691_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3863_io_b = FullAdder_3769_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3863_io_ci = FullAdder_3828_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3864_io_a = FullAdder_3771_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3864_io_b = FullAdder_3772_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3864_io_ci = HalfAdder_243_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3865_io_a = HalfAdder_223_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3865_io_b = FullAdder_3773_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3865_io_ci = FullAdder_3830_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_263_io_a = HalfAdder_225_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_263_io_b = HalfAdder_245_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3866_io_a = FullAdder_3776_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3866_io_b = HalfAdder_226_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3866_io_ci = HalfAdder_246_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3867_io_a = HalfAdder_199_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3867_io_b = HalfAdder_200_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3867_io_ci = HalfAdder_247_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3868_io_a = FullAdder_3432_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3868_io_b = FullAdder_3596_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3868_io_ci = FullAdder_3832_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_264_io_a = HalfAdder_227_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_264_io_b = HalfAdder_248_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_265_io_a = HalfAdder_228_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_265_io_b = FullAdder_3834_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_266_io_a = HalfAdder_209_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_266_io_b = FullAdder_3837_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3869_io_a = FullAdder_3717_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3869_io_b = FullAdder_3718_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3869_io_ci = FullAdder_3840_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3870_io_a = FullAdder_3789_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3870_io_b = FullAdder_3790_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3870_io_ci = FullAdder_3841_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3871_io_a = FullAdder_3791_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3871_io_b = FullAdder_3792_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3871_io_ci = FullAdder_3843_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_267_io_a = FullAdder_3794_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_267_io_b = HalfAdder_251_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3872_io_a = FullAdder_3794_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3872_io_b = HalfAdder_234_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3872_io_ci = HalfAdder_252_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3873_io_a = FullAdder_3795_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3873_io_b = FullAdder_3796_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3873_io_ci = FullAdder_3845_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_268_io_a = FullAdder_3845_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_268_io_b = HalfAdder_253_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_269_io_a = FullAdder_3797_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_269_io_b = HalfAdder_253_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3874_io_a = FullAdder_3797_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3874_io_b = FullAdder_3798_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3874_io_ci = FullAdder_3846_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3875_io_a = FullAdder_3802_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3875_io_b = FullAdder_3803_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3875_io_ci = FullAdder_3848_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3876_io_a = FullAdder_3808_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3876_io_b = FullAdder_3809_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3876_io_ci = FullAdder_3850_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_270_io_a = HalfAdder_236_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_270_io_b = FullAdder_3851_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3877_io_a = HalfAdder_238_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3877_io_b = FullAdder_3852_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3877_io_ci = HalfAdder_257_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_271_io_a = HalfAdder_257_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_271_io_b = HalfAdder_258_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3878_io_a = FullAdder_3813_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3878_io_b = FullAdder_3814_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3878_io_ci = HalfAdder_260_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3879_io_a = FullAdder_3815_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3879_io_b = HalfAdder_239_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3879_io_ci = HalfAdder_261_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_272_io_a = FullAdder_3816_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_272_io_b = HalfAdder_261_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3880_io_a = FullAdder_3816_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3880_io_b = FullAdder_3817_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3880_io_ci = FullAdder_3853_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3881_io_a = FullAdder_3754_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3881_io_b = FullAdder_3819_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3881_io_ci = FullAdder_3855_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3882_io_a = HalfAdder_240_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3882_io_b = FullAdder_3823_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3882_io_ci = FullAdder_3859_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_273_io_a = HalfAdder_243_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_273_io_b = FullAdder_3865_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3883_io_a = FullAdder_3775_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3883_io_b = FullAdder_3776_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3883_io_ci = FullAdder_3866_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3884_io_a = FullAdder_3706_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3884_io_b = HalfAdder_199_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3884_io_ci = FullAdder_3867_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3885_io_a = FullAdder_3432_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3885_io_b = FullAdder_3595_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3885_io_ci = FullAdder_3868_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3886_io_a = FullAdder_3782_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3886_io_b = HalfAdder_228_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3886_io_ci = HalfAdder_265_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3887_io_a = FullAdder_3713_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3887_io_b = HalfAdder_209_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3887_io_ci = HalfAdder_266_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3888_io_a = FullAdder_3844_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3888_io_b = HalfAdder_251_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3888_io_ci = HalfAdder_267_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_274_io_a = HalfAdder_252_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_274_io_b = FullAdder_3873_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_275_io_a = HalfAdder_268_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_275_io_b = HalfAdder_269_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3889_io_a = FullAdder_3801_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3889_io_b = FullAdder_3802_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3889_io_ci = FullAdder_3875_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3890_io_a = FullAdder_3807_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3890_io_b = FullAdder_3808_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3890_io_ci = FullAdder_3876_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3891_io_a = FullAdder_3850_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3891_io_b = FullAdder_3851_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3891_io_ci = HalfAdder_270_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_276_io_a = FullAdder_3852_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_276_io_b = HalfAdder_270_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3892_io_a = HalfAdder_258_io_co; // @[wallace.scala 69:18]
  assign FullAdder_3892_io_b = FullAdder_3877_io_s; // @[wallace.scala 70:18]
  assign FullAdder_3892_io_ci = HalfAdder_271_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_277_io_a = HalfAdder_259_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_277_io_b = HalfAdder_271_io_s; // @[wallace.scala 60:18]
  assign HalfAdder_278_io_a = HalfAdder_259_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_278_io_b = FullAdder_3878_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_279_io_a = HalfAdder_272_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_279_io_b = FullAdder_3880_io_co; // @[wallace.scala 60:18]
  assign HalfAdder_280_io_a = HalfAdder_245_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_280_io_b = FullAdder_3883_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3893_io_a = FullAdder_3705_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3893_io_b = FullAdder_3706_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3893_io_ci = FullAdder_3884_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3894_io_a = HalfAdder_172_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3894_io_b = FullAdder_3595_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3894_io_ci = FullAdder_3885_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_281_io_a = HalfAdder_248_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_281_io_b = FullAdder_3886_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3895_io_a = FullAdder_3843_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3895_io_b = FullAdder_3844_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3895_io_ci = FullAdder_3888_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3896_io_a = FullAdder_3873_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3896_io_b = HalfAdder_268_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3896_io_ci = HalfAdder_275_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_282_io_a = FullAdder_3877_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_282_io_b = HalfAdder_276_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3897_io_a = FullAdder_3879_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3897_io_b = HalfAdder_272_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3897_io_ci = HalfAdder_279_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3898_io_a = FullAdder_3704_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3898_io_b = FullAdder_3705_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3898_io_ci = FullAdder_3893_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_283_io_a = HalfAdder_264_io_s; // @[wallace.scala 59:18]
  assign HalfAdder_283_io_b = HalfAdder_281_io_co; // @[wallace.scala 60:18]
  assign FullAdder_3899_io_a = FullAdder_3891_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3899_io_b = HalfAdder_276_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3899_io_ci = HalfAdder_282_io_co; // @[wallace.scala 71:19]
  assign HalfAdder_284_io_a = FullAdder_3892_io_co; // @[wallace.scala 59:18]
  assign HalfAdder_284_io_b = HalfAdder_282_io_s; // @[wallace.scala 60:18]
  assign FullAdder_3900_io_a = HalfAdder_260_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3900_io_b = FullAdder_3879_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3900_io_ci = FullAdder_3897_io_co; // @[wallace.scala 71:19]
  assign FullAdder_3901_io_a = FullAdder_3876_io_s; // @[wallace.scala 69:18]
  assign FullAdder_3901_io_b = FullAdder_3891_io_co; // @[wallace.scala 70:18]
  assign FullAdder_3901_io_ci = FullAdder_3899_io_co; // @[wallace.scala 71:19]
endmodule
module MUL(
  input  [63:0]  io_multiplicand,
  input  [63:0]  io_multiplier,
  output [126:0] io_outs
);
  wire [63:0] pp_io_multiplicand; // @[mul.scala 26:18]
  wire [63:0] pp_io_multiplier; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_0; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_1; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_2; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_3; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_4; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_5; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_6; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_7; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_8; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_9; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_10; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_11; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_12; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_13; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_14; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_15; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_16; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_17; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_18; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_19; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_20; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_21; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_22; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_23; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_24; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_25; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_26; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_27; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_28; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_29; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_30; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_31; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_32; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_33; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_34; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_35; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_36; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_37; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_38; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_39; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_40; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_41; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_42; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_43; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_44; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_45; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_46; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_47; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_48; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_49; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_50; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_51; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_52; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_53; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_54; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_55; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_56; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_57; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_58; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_59; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_60; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_61; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_62; // @[mul.scala 26:18]
  wire [63:0] pp_io_outs_63; // @[mul.scala 26:18]
  wire [63:0] wt_io_pp_0; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_1; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_2; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_3; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_4; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_5; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_6; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_7; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_8; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_9; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_10; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_11; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_12; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_13; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_14; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_15; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_16; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_17; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_18; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_19; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_20; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_21; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_22; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_23; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_24; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_25; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_26; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_27; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_28; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_29; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_30; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_31; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_32; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_33; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_34; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_35; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_36; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_37; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_38; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_39; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_40; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_41; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_42; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_43; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_44; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_45; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_46; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_47; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_48; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_49; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_50; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_51; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_52; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_53; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_54; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_55; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_56; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_57; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_58; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_59; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_60; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_61; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_62; // @[mul.scala 30:18]
  wire [63:0] wt_io_pp_63; // @[mul.scala 30:18]
  wire [127:0] wt_io_augend; // @[mul.scala 30:18]
  wire [127:0] wt_io_addend; // @[mul.scala 30:18]
  wire [127:0] _T_1 = wt_io_augend + wt_io_addend; // @[mul.scala 37:27]
  PartialProd pp ( // @[mul.scala 26:18]
    .io_multiplicand(pp_io_multiplicand),
    .io_multiplier(pp_io_multiplier),
    .io_outs_0(pp_io_outs_0),
    .io_outs_1(pp_io_outs_1),
    .io_outs_2(pp_io_outs_2),
    .io_outs_3(pp_io_outs_3),
    .io_outs_4(pp_io_outs_4),
    .io_outs_5(pp_io_outs_5),
    .io_outs_6(pp_io_outs_6),
    .io_outs_7(pp_io_outs_7),
    .io_outs_8(pp_io_outs_8),
    .io_outs_9(pp_io_outs_9),
    .io_outs_10(pp_io_outs_10),
    .io_outs_11(pp_io_outs_11),
    .io_outs_12(pp_io_outs_12),
    .io_outs_13(pp_io_outs_13),
    .io_outs_14(pp_io_outs_14),
    .io_outs_15(pp_io_outs_15),
    .io_outs_16(pp_io_outs_16),
    .io_outs_17(pp_io_outs_17),
    .io_outs_18(pp_io_outs_18),
    .io_outs_19(pp_io_outs_19),
    .io_outs_20(pp_io_outs_20),
    .io_outs_21(pp_io_outs_21),
    .io_outs_22(pp_io_outs_22),
    .io_outs_23(pp_io_outs_23),
    .io_outs_24(pp_io_outs_24),
    .io_outs_25(pp_io_outs_25),
    .io_outs_26(pp_io_outs_26),
    .io_outs_27(pp_io_outs_27),
    .io_outs_28(pp_io_outs_28),
    .io_outs_29(pp_io_outs_29),
    .io_outs_30(pp_io_outs_30),
    .io_outs_31(pp_io_outs_31),
    .io_outs_32(pp_io_outs_32),
    .io_outs_33(pp_io_outs_33),
    .io_outs_34(pp_io_outs_34),
    .io_outs_35(pp_io_outs_35),
    .io_outs_36(pp_io_outs_36),
    .io_outs_37(pp_io_outs_37),
    .io_outs_38(pp_io_outs_38),
    .io_outs_39(pp_io_outs_39),
    .io_outs_40(pp_io_outs_40),
    .io_outs_41(pp_io_outs_41),
    .io_outs_42(pp_io_outs_42),
    .io_outs_43(pp_io_outs_43),
    .io_outs_44(pp_io_outs_44),
    .io_outs_45(pp_io_outs_45),
    .io_outs_46(pp_io_outs_46),
    .io_outs_47(pp_io_outs_47),
    .io_outs_48(pp_io_outs_48),
    .io_outs_49(pp_io_outs_49),
    .io_outs_50(pp_io_outs_50),
    .io_outs_51(pp_io_outs_51),
    .io_outs_52(pp_io_outs_52),
    .io_outs_53(pp_io_outs_53),
    .io_outs_54(pp_io_outs_54),
    .io_outs_55(pp_io_outs_55),
    .io_outs_56(pp_io_outs_56),
    .io_outs_57(pp_io_outs_57),
    .io_outs_58(pp_io_outs_58),
    .io_outs_59(pp_io_outs_59),
    .io_outs_60(pp_io_outs_60),
    .io_outs_61(pp_io_outs_61),
    .io_outs_62(pp_io_outs_62),
    .io_outs_63(pp_io_outs_63)
  );
  Wallace wt ( // @[mul.scala 30:18]
    .io_pp_0(wt_io_pp_0),
    .io_pp_1(wt_io_pp_1),
    .io_pp_2(wt_io_pp_2),
    .io_pp_3(wt_io_pp_3),
    .io_pp_4(wt_io_pp_4),
    .io_pp_5(wt_io_pp_5),
    .io_pp_6(wt_io_pp_6),
    .io_pp_7(wt_io_pp_7),
    .io_pp_8(wt_io_pp_8),
    .io_pp_9(wt_io_pp_9),
    .io_pp_10(wt_io_pp_10),
    .io_pp_11(wt_io_pp_11),
    .io_pp_12(wt_io_pp_12),
    .io_pp_13(wt_io_pp_13),
    .io_pp_14(wt_io_pp_14),
    .io_pp_15(wt_io_pp_15),
    .io_pp_16(wt_io_pp_16),
    .io_pp_17(wt_io_pp_17),
    .io_pp_18(wt_io_pp_18),
    .io_pp_19(wt_io_pp_19),
    .io_pp_20(wt_io_pp_20),
    .io_pp_21(wt_io_pp_21),
    .io_pp_22(wt_io_pp_22),
    .io_pp_23(wt_io_pp_23),
    .io_pp_24(wt_io_pp_24),
    .io_pp_25(wt_io_pp_25),
    .io_pp_26(wt_io_pp_26),
    .io_pp_27(wt_io_pp_27),
    .io_pp_28(wt_io_pp_28),
    .io_pp_29(wt_io_pp_29),
    .io_pp_30(wt_io_pp_30),
    .io_pp_31(wt_io_pp_31),
    .io_pp_32(wt_io_pp_32),
    .io_pp_33(wt_io_pp_33),
    .io_pp_34(wt_io_pp_34),
    .io_pp_35(wt_io_pp_35),
    .io_pp_36(wt_io_pp_36),
    .io_pp_37(wt_io_pp_37),
    .io_pp_38(wt_io_pp_38),
    .io_pp_39(wt_io_pp_39),
    .io_pp_40(wt_io_pp_40),
    .io_pp_41(wt_io_pp_41),
    .io_pp_42(wt_io_pp_42),
    .io_pp_43(wt_io_pp_43),
    .io_pp_44(wt_io_pp_44),
    .io_pp_45(wt_io_pp_45),
    .io_pp_46(wt_io_pp_46),
    .io_pp_47(wt_io_pp_47),
    .io_pp_48(wt_io_pp_48),
    .io_pp_49(wt_io_pp_49),
    .io_pp_50(wt_io_pp_50),
    .io_pp_51(wt_io_pp_51),
    .io_pp_52(wt_io_pp_52),
    .io_pp_53(wt_io_pp_53),
    .io_pp_54(wt_io_pp_54),
    .io_pp_55(wt_io_pp_55),
    .io_pp_56(wt_io_pp_56),
    .io_pp_57(wt_io_pp_57),
    .io_pp_58(wt_io_pp_58),
    .io_pp_59(wt_io_pp_59),
    .io_pp_60(wt_io_pp_60),
    .io_pp_61(wt_io_pp_61),
    .io_pp_62(wt_io_pp_62),
    .io_pp_63(wt_io_pp_63),
    .io_augend(wt_io_augend),
    .io_addend(wt_io_addend)
  );
  assign io_outs = _T_1[126:0]; // @[mul.scala 37:11]
  assign pp_io_multiplicand = io_multiplicand; // @[mul.scala 27:22]
  assign pp_io_multiplier = io_multiplier; // @[mul.scala 28:20]
  assign wt_io_pp_0 = pp_io_outs_0; // @[mul.scala 31:12]
  assign wt_io_pp_1 = pp_io_outs_1; // @[mul.scala 31:12]
  assign wt_io_pp_2 = pp_io_outs_2; // @[mul.scala 31:12]
  assign wt_io_pp_3 = pp_io_outs_3; // @[mul.scala 31:12]
  assign wt_io_pp_4 = pp_io_outs_4; // @[mul.scala 31:12]
  assign wt_io_pp_5 = pp_io_outs_5; // @[mul.scala 31:12]
  assign wt_io_pp_6 = pp_io_outs_6; // @[mul.scala 31:12]
  assign wt_io_pp_7 = pp_io_outs_7; // @[mul.scala 31:12]
  assign wt_io_pp_8 = pp_io_outs_8; // @[mul.scala 31:12]
  assign wt_io_pp_9 = pp_io_outs_9; // @[mul.scala 31:12]
  assign wt_io_pp_10 = pp_io_outs_10; // @[mul.scala 31:12]
  assign wt_io_pp_11 = pp_io_outs_11; // @[mul.scala 31:12]
  assign wt_io_pp_12 = pp_io_outs_12; // @[mul.scala 31:12]
  assign wt_io_pp_13 = pp_io_outs_13; // @[mul.scala 31:12]
  assign wt_io_pp_14 = pp_io_outs_14; // @[mul.scala 31:12]
  assign wt_io_pp_15 = pp_io_outs_15; // @[mul.scala 31:12]
  assign wt_io_pp_16 = pp_io_outs_16; // @[mul.scala 31:12]
  assign wt_io_pp_17 = pp_io_outs_17; // @[mul.scala 31:12]
  assign wt_io_pp_18 = pp_io_outs_18; // @[mul.scala 31:12]
  assign wt_io_pp_19 = pp_io_outs_19; // @[mul.scala 31:12]
  assign wt_io_pp_20 = pp_io_outs_20; // @[mul.scala 31:12]
  assign wt_io_pp_21 = pp_io_outs_21; // @[mul.scala 31:12]
  assign wt_io_pp_22 = pp_io_outs_22; // @[mul.scala 31:12]
  assign wt_io_pp_23 = pp_io_outs_23; // @[mul.scala 31:12]
  assign wt_io_pp_24 = pp_io_outs_24; // @[mul.scala 31:12]
  assign wt_io_pp_25 = pp_io_outs_25; // @[mul.scala 31:12]
  assign wt_io_pp_26 = pp_io_outs_26; // @[mul.scala 31:12]
  assign wt_io_pp_27 = pp_io_outs_27; // @[mul.scala 31:12]
  assign wt_io_pp_28 = pp_io_outs_28; // @[mul.scala 31:12]
  assign wt_io_pp_29 = pp_io_outs_29; // @[mul.scala 31:12]
  assign wt_io_pp_30 = pp_io_outs_30; // @[mul.scala 31:12]
  assign wt_io_pp_31 = pp_io_outs_31; // @[mul.scala 31:12]
  assign wt_io_pp_32 = pp_io_outs_32; // @[mul.scala 31:12]
  assign wt_io_pp_33 = pp_io_outs_33; // @[mul.scala 31:12]
  assign wt_io_pp_34 = pp_io_outs_34; // @[mul.scala 31:12]
  assign wt_io_pp_35 = pp_io_outs_35; // @[mul.scala 31:12]
  assign wt_io_pp_36 = pp_io_outs_36; // @[mul.scala 31:12]
  assign wt_io_pp_37 = pp_io_outs_37; // @[mul.scala 31:12]
  assign wt_io_pp_38 = pp_io_outs_38; // @[mul.scala 31:12]
  assign wt_io_pp_39 = pp_io_outs_39; // @[mul.scala 31:12]
  assign wt_io_pp_40 = pp_io_outs_40; // @[mul.scala 31:12]
  assign wt_io_pp_41 = pp_io_outs_41; // @[mul.scala 31:12]
  assign wt_io_pp_42 = pp_io_outs_42; // @[mul.scala 31:12]
  assign wt_io_pp_43 = pp_io_outs_43; // @[mul.scala 31:12]
  assign wt_io_pp_44 = pp_io_outs_44; // @[mul.scala 31:12]
  assign wt_io_pp_45 = pp_io_outs_45; // @[mul.scala 31:12]
  assign wt_io_pp_46 = pp_io_outs_46; // @[mul.scala 31:12]
  assign wt_io_pp_47 = pp_io_outs_47; // @[mul.scala 31:12]
  assign wt_io_pp_48 = pp_io_outs_48; // @[mul.scala 31:12]
  assign wt_io_pp_49 = pp_io_outs_49; // @[mul.scala 31:12]
  assign wt_io_pp_50 = pp_io_outs_50; // @[mul.scala 31:12]
  assign wt_io_pp_51 = pp_io_outs_51; // @[mul.scala 31:12]
  assign wt_io_pp_52 = pp_io_outs_52; // @[mul.scala 31:12]
  assign wt_io_pp_53 = pp_io_outs_53; // @[mul.scala 31:12]
  assign wt_io_pp_54 = pp_io_outs_54; // @[mul.scala 31:12]
  assign wt_io_pp_55 = pp_io_outs_55; // @[mul.scala 31:12]
  assign wt_io_pp_56 = pp_io_outs_56; // @[mul.scala 31:12]
  assign wt_io_pp_57 = pp_io_outs_57; // @[mul.scala 31:12]
  assign wt_io_pp_58 = pp_io_outs_58; // @[mul.scala 31:12]
  assign wt_io_pp_59 = pp_io_outs_59; // @[mul.scala 31:12]
  assign wt_io_pp_60 = pp_io_outs_60; // @[mul.scala 31:12]
  assign wt_io_pp_61 = pp_io_outs_61; // @[mul.scala 31:12]
  assign wt_io_pp_62 = pp_io_outs_62; // @[mul.scala 31:12]
  assign wt_io_pp_63 = pp_io_outs_63; // @[mul.scala 31:12]
endmodule
