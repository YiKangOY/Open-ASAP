module kn32 (in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, out30, out31, out32, );
input in0;
input in1;
input in2;
input in3;
input in4;
input in5;
input in6;
input in7;
input in8;
input in9;
input in10;
input in11;
input in12;
input in13;
input in14;
input in15;
input in16;
input in17;
input in18;
input in19;
input in20;
input in21;
input in22;
input in23;
input in24;
input in25;
input in26;
input in27;
input in28;
input in29;
input in30;
input in31;
input in32;
input in33;
input in34;
input in35;
input in36;
input in37;
input in38;
input in39;
input in40;
input in41;
input in42;
input in43;
input in44;
input in45;
input in46;
input in47;
input in48;
input in49;
input in50;
input in51;
input in52;
input in53;
input in54;
input in55;
input in56;
input in57;
input in58;
input in59;
input in60;
input in61;
input in62;
input in63;
output out0;
output out1;
output out2;
output out3;
output out4;
output out5;
output out6;
output out7;
output out8;
output out9;
output out10;
output out11;
output out12;
output out13;
output out14;
output out15;
output out16;
output out17;
output out18;
output out19;
output out20;
output out21;
output out22;
output out23;
output out24;
output out25;
output out26;
output out27;
output out28;
output out29;
output out30;
output out31;
output out32;
wire var0;
wire var1;
wire var2;
wire var3;
wire var4;
wire var5;
wire var6;
wire var7;
wire var8;
wire var9;
wire var10;
wire var11;
wire var12;
wire var13;
wire var14;
wire var15;
wire var16;
wire var17;
wire var18;
wire var19;
wire var20;
wire var21;
wire var22;
wire var23;
wire var24;
wire var25;
wire var26;
wire var27;
wire var28;
wire var29;
wire var30;
wire var31;
wire var32;
wire var33;
wire var34;
wire var35;
wire var36;
wire var37;
wire var38;
wire var39;
wire var40;
wire var41;
wire var42;
wire var43;
wire var44;
wire var45;
wire var46;
wire var47;
wire var48;
wire var49;
wire var50;
wire var51;
wire var52;
wire var53;
wire var54;
wire var55;
wire var56;
wire var57;
wire var58;
wire var59;
wire var60;
wire var61;
wire var62;
wire var63;
wire var64;
wire var65;
wire var66;
wire var67;
wire var68;
wire var69;
wire var70;
wire var71;
wire var72;
wire var73;
wire var74;
wire var75;
wire var76;
wire var77;
wire var78;
wire var79;
wire var80;
wire var81;
wire var82;
wire var83;
wire var84;
wire var85;
wire var86;
wire var87;
wire var88;
wire var89;
wire var90;
wire var91;
wire var92;
wire var93;
wire var94;
wire var95;
wire var96;
wire var97;
wire var98;
wire var99;
wire var100;
wire var101;
wire var102;
wire var103;
wire var104;
wire var105;
wire var106;
wire var107;
wire var108;
wire var109;
wire var110;
wire var111;
wire var112;
wire var113;
wire var114;
wire var115;
wire var116;
wire var117;
wire var118;
wire var119;
wire var120;
wire var121;
wire var122;
wire var123;
wire var124;
wire var125;
wire var126;
wire var127;
wire var128;
wire var129;
wire var130;
wire var131;
wire var132;
wire var133;
wire var134;
wire var135;
wire var136;
wire var137;
wire var138;
wire var139;
wire var140;
wire var141;
wire var142;
wire var143;
wire var144;
wire var145;
wire var146;
wire var147;
wire var148;
wire var149;
wire var150;
wire var151;
wire var152;
wire var153;
wire var154;
wire var155;
wire var156;
wire var157;
wire var158;
wire var159;
wire var160;
wire var161;
wire var162;
wire var163;
wire var164;
wire var165;
wire var166;
wire var167;
wire var168;
wire var169;
wire var170;
wire var171;
wire var172;
wire var173;
wire var174;
wire var175;
wire var176;
wire var177;
wire var178;
wire var179;
wire var180;
wire var181;
wire var182;
wire var183;
wire var184;
wire var185;
wire var186;
wire var187;
wire var188;
wire var189;
wire var190;
wire var191;
wire var192;
wire var193;
wire var194;
wire var195;
wire var196;
wire var197;
wire var198;
wire var199;
wire var200;
wire var201;
wire var202;
wire var203;
wire var204;
wire var205;
wire var206;
wire var207;
wire var208;
wire var209;
wire var210;
wire var211;
wire var212;
wire var213;
wire var214;
wire var215;
wire var216;
wire var217;
wire var218;
wire var219;
wire var220;
wire var221;
wire var222;
wire var223;
wire var224;
wire var225;
wire var226;
wire var227;
wire var228;
wire var229;
wire var230;
wire var231;
wire var232;
wire var233;
wire var234;
wire var235;
wire var236;
wire var237;
wire var238;
wire var239;
wire var240;
wire var241;
wire var242;
wire var243;
wire var244;
wire var245;
wire var246;
wire var247;
wire var248;
wire var249;
wire var250;
wire var251;
wire var252;
wire var253;
wire var254;
wire var255;
wire var256;
wire var257;
wire var258;
wire var259;
wire var260;
wire var261;
wire var262;
wire var263;
wire var264;
wire var265;
wire var266;
wire var267;
wire var268;
wire var269;
wire var270;
wire var271;
wire var272;
wire var273;
wire var274;
wire var275;
wire var276;
wire var277;
wire var278;
wire var279;
wire var280;
wire var281;
wire var282;
wire var283;
wire var284;
wire var285;
wire var286;
wire var287;
wire var288;
wire var289;
wire var290;
wire var291;
wire var292;
wire var293;
wire var294;
wire var295;
wire var296;
wire var297;
wire var298;
wire var299;
wire var300;
wire var301;
wire var302;
wire var303;
wire var304;
wire var305;
wire var306;
wire var307;
wire var308;
wire var309;
wire var310;
wire var311;
wire var312;
wire var313;
wire var314;
wire var315;
wire var316;
wire var317;
wire var318;
wire var319;
wire var320;
wire var321;
wire var322;
wire var323;
wire var324;
wire var325;
wire var326;
wire var327;
wire var328;
wire var329;
wire var330;
wire var331;
wire var332;
wire var333;
wire var334;
wire var335;
wire var336;
wire var337;
wire var338;
wire var339;
wire var340;
wire var341;
wire var342;
wire var343;
wire var344;
wire var345;
wire var346;
wire var347;
wire var348;
wire var349;
wire var350;
wire var351;
wire var352;
wire var353;
wire var354;
wire var355;
wire var356;
wire var357;
wire var358;
wire var359;
wire var360;
wire var361;
wire var362;
wire var363;
wire var364;
wire var365;
wire var366;
wire var367;
wire var368;
wire var369;
wire var370;
wire var371;
wire var372;
wire var373;
wire var374;
wire var375;
wire var376;
wire var377;
wire var378;
wire var379;
wire var380;
wire var381;
wire var382;
wire var383;
wire var384;
wire var385;
wire var386;
wire var387;
wire var388;
wire var389;
wire var390;
wire var391;
wire var392;
wire var393;
wire var394;
wire var395;
wire var396;
wire var397;
wire var398;
wire var399;
wire var400;
wire var401;
wire var402;
wire var403;
wire var404;
wire var405;
wire var406;
wire var407;
wire var408;
wire var409;
wire var410;
wire var411;
wire var412;
wire var413;
wire var414;
wire var415;
wire var416;
wire var417;
wire var418;
wire var419;
wire var420;
wire var421;
wire var422;
wire var423;
wire var424;
wire var425;
wire var426;
assign var0 = in63 & in31;
assign var1 = in62 & in30;
assign var2 = in61 & in29;
assign var3 = in60 & in28;
assign var4 = in59 & in27;
assign var5 = in58 & in26;
assign var6 = in57 & in25;
assign var7 = in56 & in24;
assign var8 = in55 & in23;
assign var9 = in54 & in22;
assign var10 = in53 & in21;
assign var11 = in52 & in20;
assign var12 = in51 & in19;
assign var13 = in50 & in18;
assign var14 = in49 & in17;
assign var15 = in48 & in16;
assign var16 = in47 & in15;
assign var17 = in46 & in14;
assign var18 = in45 & in13;
assign var19 = in44 & in12;
assign var20 = in43 & in11;
assign var21 = in42 & in10;
assign var22 = in41 & in9;
assign var23 = in40 & in8;
assign var24 = in39 & in7;
assign var25 = in38 & in6;
assign var26 = in37 & in5;
assign var27 = in36 & in4;
assign var28 = in35 & in3;
assign var29 = in34 & in2;
assign var30 = in33 & in1;
assign var31 = in32 & in0;
assign var32 = in63 ^ in31;
assign var33 = in62 ^ in30;
assign var34 = in61 ^ in29;
assign var35 = in60 ^ in28;
assign var36 = in59 ^ in27;
assign var37 = in58 ^ in26;
assign var38 = in57 ^ in25;
assign var39 = in56 ^ in24;
assign var40 = in55 ^ in23;
assign var41 = in54 ^ in22;
assign var42 = in53 ^ in21;
assign var43 = in52 ^ in20;
assign var44 = in51 ^ in19;
assign var45 = in50 ^ in18;
assign var46 = in49 ^ in17;
assign var47 = in48 ^ in16;
assign var48 = in47 ^ in15;
assign var49 = in46 ^ in14;
assign var50 = in45 ^ in13;
assign var51 = in44 ^ in12;
assign var52 = in43 ^ in11;
assign var53 = in42 ^ in10;
assign var54 = in41 ^ in9;
assign var55 = in40 ^ in8;
assign var56 = in39 ^ in7;
assign var57 = in38 ^ in6;
assign var58 = in37 ^ in5;
assign var59 = in36 ^ in4;
assign var60 = in35 ^ in3;
assign var61 = in34 ^ in2;
assign var62 = in33 ^ in1;
assign var63 = in32 ^ in0;
assign var64 = var63 & var30;
assign var65 = var31 | var64;
assign var66 = var63 & var62;
assign var67 = var62 & var29;
assign var68 = var30 | var67;
assign var69 = var62 & var61;
assign var70 = var61 & var28;
assign var71 = var29 | var70;
assign var72 = var61 & var60;
assign var73 = var60 & var27;
assign var74 = var28 | var73;
assign var75 = var60 & var59;
assign var76 = var59 & var26;
assign var77 = var27 | var76;
assign var78 = var59 & var58;
assign var79 = var58 & var25;
assign var80 = var26 | var79;
assign var81 = var58 & var57;
assign var82 = var57 & var24;
assign var83 = var25 | var82;
assign var84 = var57 & var56;
assign var85 = var56 & var23;
assign var86 = var24 | var85;
assign var87 = var56 & var55;
assign var88 = var55 & var22;
assign var89 = var23 | var88;
assign var90 = var55 & var54;
assign var91 = var54 & var21;
assign var92 = var22 | var91;
assign var93 = var54 & var53;
assign var94 = var53 & var20;
assign var95 = var21 | var94;
assign var96 = var53 & var52;
assign var97 = var52 & var19;
assign var98 = var20 | var97;
assign var99 = var52 & var51;
assign var100 = var51 & var18;
assign var101 = var19 | var100;
assign var102 = var51 & var50;
assign var103 = var50 & var17;
assign var104 = var18 | var103;
assign var105 = var50 & var49;
assign var106 = var49 & var16;
assign var107 = var17 | var106;
assign var108 = var49 & var48;
assign var109 = var48 & var15;
assign var110 = var16 | var109;
assign var111 = var48 & var47;
assign var112 = var47 & var14;
assign var113 = var15 | var112;
assign var114 = var47 & var46;
assign var115 = var46 & var13;
assign var116 = var14 | var115;
assign var117 = var46 & var45;
assign var118 = var45 & var12;
assign var119 = var13 | var118;
assign var120 = var45 & var44;
assign var121 = var44 & var11;
assign var122 = var12 | var121;
assign var123 = var44 & var43;
assign var124 = var43 & var10;
assign var125 = var11 | var124;
assign var126 = var43 & var42;
assign var127 = var42 & var9;
assign var128 = var10 | var127;
assign var129 = var42 & var41;
assign var130 = var41 & var8;
assign var131 = var9 | var130;
assign var132 = var41 & var40;
assign var133 = var40 & var7;
assign var134 = var8 | var133;
assign var135 = var40 & var39;
assign var136 = var39 & var6;
assign var137 = var7 | var136;
assign var138 = var39 & var38;
assign var139 = var38 & var5;
assign var140 = var6 | var139;
assign var141 = var38 & var37;
assign var142 = var37 & var4;
assign var143 = var5 | var142;
assign var144 = var37 & var36;
assign var145 = var36 & var3;
assign var146 = var4 | var145;
assign var147 = var36 & var35;
assign var148 = var35 & var2;
assign var149 = var3 | var148;
assign var150 = var35 & var34;
assign var151 = var34 & var1;
assign var152 = var2 | var151;
assign var153 = var34 & var33;
assign var154 = var33 & var0;
assign var155 = var1 | var154;
assign var156 = var66 & var71;
assign var157 = var65 | var156;
assign var158 = var66 & var72;
assign var159 = var69 & var74;
assign var160 = var68 | var159;
assign var161 = var69 & var75;
assign var162 = var72 & var77;
assign var163 = var71 | var162;
assign var164 = var72 & var78;
assign var165 = var75 & var80;
assign var166 = var74 | var165;
assign var167 = var75 & var81;
assign var168 = var78 & var83;
assign var169 = var77 | var168;
assign var170 = var78 & var84;
assign var171 = var81 & var86;
assign var172 = var80 | var171;
assign var173 = var81 & var87;
assign var174 = var84 & var89;
assign var175 = var83 | var174;
assign var176 = var84 & var90;
assign var177 = var87 & var92;
assign var178 = var86 | var177;
assign var179 = var87 & var93;
assign var180 = var90 & var95;
assign var181 = var89 | var180;
assign var182 = var90 & var96;
assign var183 = var93 & var98;
assign var184 = var92 | var183;
assign var185 = var93 & var99;
assign var186 = var96 & var101;
assign var187 = var95 | var186;
assign var188 = var96 & var102;
assign var189 = var99 & var104;
assign var190 = var98 | var189;
assign var191 = var99 & var105;
assign var192 = var102 & var107;
assign var193 = var101 | var192;
assign var194 = var102 & var108;
assign var195 = var105 & var110;
assign var196 = var104 | var195;
assign var197 = var105 & var111;
assign var198 = var108 & var113;
assign var199 = var107 | var198;
assign var200 = var108 & var114;
assign var201 = var111 & var116;
assign var202 = var110 | var201;
assign var203 = var111 & var117;
assign var204 = var114 & var119;
assign var205 = var113 | var204;
assign var206 = var114 & var120;
assign var207 = var117 & var122;
assign var208 = var116 | var207;
assign var209 = var117 & var123;
assign var210 = var120 & var125;
assign var211 = var119 | var210;
assign var212 = var120 & var126;
assign var213 = var123 & var128;
assign var214 = var122 | var213;
assign var215 = var123 & var129;
assign var216 = var126 & var131;
assign var217 = var125 | var216;
assign var218 = var126 & var132;
assign var219 = var129 & var134;
assign var220 = var128 | var219;
assign var221 = var129 & var135;
assign var222 = var132 & var137;
assign var223 = var131 | var222;
assign var224 = var132 & var138;
assign var225 = var135 & var140;
assign var226 = var134 | var225;
assign var227 = var135 & var141;
assign var228 = var138 & var143;
assign var229 = var137 | var228;
assign var230 = var138 & var144;
assign var231 = var141 & var146;
assign var232 = var140 | var231;
assign var233 = var141 & var147;
assign var234 = var144 & var149;
assign var235 = var143 | var234;
assign var236 = var144 & var150;
assign var237 = var147 & var152;
assign var238 = var146 | var237;
assign var239 = var147 & var153;
assign var240 = var150 & var155;
assign var241 = var149 | var240;
assign var242 = var153 & var0;
assign var243 = var152 | var242;
assign var244 = var158 & var169;
assign var245 = var157 | var244;
assign var246 = var158 & var170;
assign var247 = var161 & var172;
assign var248 = var160 | var247;
assign var249 = var161 & var173;
assign var250 = var164 & var175;
assign var251 = var163 | var250;
assign var252 = var164 & var176;
assign var253 = var167 & var178;
assign var254 = var166 | var253;
assign var255 = var167 & var179;
assign var256 = var170 & var181;
assign var257 = var169 | var256;
assign var258 = var170 & var182;
assign var259 = var173 & var184;
assign var260 = var172 | var259;
assign var261 = var173 & var185;
assign var262 = var176 & var187;
assign var263 = var175 | var262;
assign var264 = var176 & var188;
assign var265 = var179 & var190;
assign var266 = var178 | var265;
assign var267 = var179 & var191;
assign var268 = var182 & var193;
assign var269 = var181 | var268;
assign var270 = var182 & var194;
assign var271 = var185 & var196;
assign var272 = var184 | var271;
assign var273 = var185 & var197;
assign var274 = var188 & var199;
assign var275 = var187 | var274;
assign var276 = var188 & var200;
assign var277 = var191 & var202;
assign var278 = var190 | var277;
assign var279 = var191 & var203;
assign var280 = var194 & var205;
assign var281 = var193 | var280;
assign var282 = var194 & var206;
assign var283 = var197 & var208;
assign var284 = var196 | var283;
assign var285 = var197 & var209;
assign var286 = var200 & var211;
assign var287 = var199 | var286;
assign var288 = var200 & var212;
assign var289 = var203 & var214;
assign var290 = var202 | var289;
assign var291 = var203 & var215;
assign var292 = var206 & var217;
assign var293 = var205 | var292;
assign var294 = var206 & var218;
assign var295 = var209 & var220;
assign var296 = var208 | var295;
assign var297 = var209 & var221;
assign var298 = var212 & var223;
assign var299 = var211 | var298;
assign var300 = var212 & var224;
assign var301 = var215 & var226;
assign var302 = var214 | var301;
assign var303 = var215 & var227;
assign var304 = var218 & var229;
assign var305 = var217 | var304;
assign var306 = var218 & var230;
assign var307 = var221 & var232;
assign var308 = var220 | var307;
assign var309 = var221 & var233;
assign var310 = var224 & var235;
assign var311 = var223 | var310;
assign var312 = var224 & var236;
assign var313 = var227 & var238;
assign var314 = var226 | var313;
assign var315 = var227 & var239;
assign var316 = var230 & var241;
assign var317 = var229 | var316;
assign var318 = var233 & var243;
assign var319 = var232 | var318;
assign var320 = var236 & var155;
assign var321 = var235 | var320;
assign var322 = var239 & var0;
assign var323 = var238 | var322;
assign var324 = var246 & var269;
assign var325 = var245 | var324;
assign var326 = var246 & var270;
assign var327 = var249 & var272;
assign var328 = var248 | var327;
assign var329 = var249 & var273;
assign var330 = var252 & var275;
assign var331 = var251 | var330;
assign var332 = var252 & var276;
assign var333 = var255 & var278;
assign var334 = var254 | var333;
assign var335 = var255 & var279;
assign var336 = var258 & var281;
assign var337 = var257 | var336;
assign var338 = var258 & var282;
assign var339 = var261 & var284;
assign var340 = var260 | var339;
assign var341 = var261 & var285;
assign var342 = var264 & var287;
assign var343 = var263 | var342;
assign var344 = var264 & var288;
assign var345 = var267 & var290;
assign var346 = var266 | var345;
assign var347 = var267 & var291;
assign var348 = var294 & var317;
assign var349 = var293 | var348;
assign var350 = var297 & var319;
assign var351 = var296 | var350;
assign var352 = var300 & var321;
assign var353 = var299 | var352;
assign var354 = var303 & var323;
assign var355 = var302 | var354;
assign var356 = var306 & var241;
assign var357 = var305 | var356;
assign var358 = var309 & var243;
assign var359 = var308 | var358;
assign var360 = var312 & var155;
assign var361 = var311 | var360;
assign var362 = var315 & var0;
assign var363 = var314 | var362;
assign var364 = var326 & var349;
assign var365 = var325 | var364;
assign var366 = var329 & var349;
assign var367 = var328 | var366;
assign var368 = var332 & var349;
assign var369 = var331 | var368;
assign var370 = var335 & var349;
assign var371 = var334 | var370;
assign var372 = var338 & var349;
assign var373 = var337 | var372;
assign var374 = var341 & var349;
assign var375 = var340 | var374;
assign var376 = var344 & var349;
assign var377 = var343 | var376;
assign var378 = var347 & var349;
assign var379 = var346 | var378;
assign var380 = var270 & var349;
assign var381 = var269 | var380;
assign var382 = var273 & var349;
assign var383 = var272 | var382;
assign var384 = var276 & var349;
assign var385 = var275 | var384;
assign var386 = var279 & var349;
assign var387 = var278 | var386;
assign var388 = var282 & var349;
assign var389 = var281 | var388;
assign var390 = var285 & var349;
assign var391 = var284 | var390;
assign var392 = var288 & var349;
assign var393 = var287 | var392;
assign var394 = var291 & var349;
assign var395 = var290 | var394;
assign var396 = var33 ^ var0;
assign var397 = var34 ^ var155;
assign var398 = var35 ^ var243;
assign var399 = var36 ^ var241;
assign var400 = var37 ^ var323;
assign var401 = var38 ^ var321;
assign var402 = var39 ^ var319;
assign var403 = var40 ^ var317;
assign var404 = var41 ^ var363;
assign var405 = var42 ^ var361;
assign var406 = var43 ^ var359;
assign var407 = var44 ^ var357;
assign var408 = var45 ^ var355;
assign var409 = var46 ^ var353;
assign var410 = var47 ^ var351;
assign var411 = var48 ^ var349;
assign var412 = var49 ^ var395;
assign var413 = var50 ^ var393;
assign var414 = var51 ^ var391;
assign var415 = var52 ^ var389;
assign var416 = var53 ^ var387;
assign var417 = var54 ^ var385;
assign var418 = var55 ^ var383;
assign var419 = var56 ^ var381;
assign var420 = var57 ^ var379;
assign var421 = var58 ^ var377;
assign var422 = var59 ^ var375;
assign var423 = var60 ^ var373;
assign var424 = var61 ^ var371;
assign var425 = var62 ^ var369;
assign var426 = var63 ^ var367;
assign out0 = var365;
assign out1 = var426;
assign out2 = var425;
assign out3 = var424;
assign out4 = var423;
assign out5 = var422;
assign out6 = var421;
assign out7 = var420;
assign out8 = var419;
assign out9 = var418;
assign out10 = var417;
assign out11 = var416;
assign out12 = var415;
assign out13 = var414;
assign out14 = var413;
assign out15 = var412;
assign out16 = var411;
assign out17 = var410;
assign out18 = var409;
assign out19 = var408;
assign out20 = var407;
assign out21 = var406;
assign out22 = var405;
assign out23 = var404;
assign out24 = var403;
assign out25 = var402;
assign out26 = var401;
assign out27 = var400;
assign out28 = var399;
assign out29 = var398;
assign out30 = var397;
assign out31 = var396;
assign out32 = var32;
endmodule 
